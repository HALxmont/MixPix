magic
tech sky130B
magscale 1 2
timestamp 1668043855
<< viali >>
rect 5273 57409 5307 57443
rect 15209 57409 15243 57443
rect 25145 57409 25179 57443
rect 35081 57409 35115 57443
rect 45017 57409 45051 57443
rect 55321 57409 55355 57443
rect 64889 57409 64923 57443
rect 67005 57409 67039 57443
rect 67649 57409 67683 57443
rect 68109 56797 68143 56831
rect 67649 55097 67683 55131
rect 67649 53941 67683 53975
rect 68109 52445 68143 52479
rect 68109 51357 68143 51391
rect 67649 49725 67683 49759
rect 67649 48501 67683 48535
rect 68109 47005 68143 47039
rect 68109 45917 68143 45951
rect 67649 44217 67683 44251
rect 67649 43061 67683 43095
rect 68109 41565 68143 41599
rect 68109 40477 68143 40511
rect 67649 38777 67683 38811
rect 67649 37621 67683 37655
rect 68109 36125 68143 36159
rect 68109 35037 68143 35071
rect 67649 33337 67683 33371
rect 67649 32181 67683 32215
rect 20913 31909 20947 31943
rect 21373 31841 21407 31875
rect 20545 31773 20579 31807
rect 21603 31773 21637 31807
rect 21738 31773 21772 31807
rect 21854 31770 21888 31804
rect 22017 31773 22051 31807
rect 23121 31773 23155 31807
rect 23305 31773 23339 31807
rect 15117 31705 15151 31739
rect 15301 31705 15335 31739
rect 20729 31705 20763 31739
rect 22569 31705 22603 31739
rect 15485 31637 15519 31671
rect 19349 31637 19383 31671
rect 23489 31637 23523 31671
rect 13001 31365 13035 31399
rect 3994 31297 4028 31331
rect 12817 31297 12851 31331
rect 15393 31297 15427 31331
rect 15485 31297 15519 31331
rect 15577 31297 15611 31331
rect 15761 31297 15795 31331
rect 17417 31297 17451 31331
rect 17601 31297 17635 31331
rect 18521 31297 18555 31331
rect 18613 31297 18647 31331
rect 18705 31297 18739 31331
rect 18889 31297 18923 31331
rect 19349 31297 19383 31331
rect 19533 31297 19567 31331
rect 19625 31297 19659 31331
rect 19717 31297 19751 31331
rect 23489 31297 23523 31331
rect 23673 31297 23707 31331
rect 23784 31297 23818 31331
rect 23877 31297 23911 31331
rect 4261 31229 4295 31263
rect 17785 31229 17819 31263
rect 16773 31161 16807 31195
rect 24133 31161 24167 31195
rect 2881 31093 2915 31127
rect 13185 31093 13219 31127
rect 15117 31093 15151 31127
rect 18245 31093 18279 31127
rect 19993 31093 20027 31127
rect 24593 31093 24627 31127
rect 15485 30889 15519 30923
rect 19625 30889 19659 30923
rect 6745 30685 6779 30719
rect 11437 30685 11471 30719
rect 14105 30685 14139 30719
rect 16405 30685 16439 30719
rect 16672 30685 16706 30719
rect 19257 30685 19291 30719
rect 22486 30685 22520 30719
rect 22753 30685 22787 30719
rect 68109 30685 68143 30719
rect 7012 30617 7046 30651
rect 9505 30617 9539 30651
rect 9689 30617 9723 30651
rect 11704 30617 11738 30651
rect 14372 30617 14406 30651
rect 19441 30617 19475 30651
rect 8125 30549 8159 30583
rect 9873 30549 9907 30583
rect 12817 30549 12851 30583
rect 17785 30549 17819 30583
rect 21373 30549 21407 30583
rect 24501 30345 24535 30379
rect 1593 30277 1627 30311
rect 2605 30277 2639 30311
rect 13185 30277 13219 30311
rect 15577 30277 15611 30311
rect 20646 30277 20680 30311
rect 21833 30277 21867 30311
rect 1777 30209 1811 30243
rect 2789 30209 2823 30243
rect 4445 30209 4479 30243
rect 4712 30209 4746 30243
rect 9321 30209 9355 30243
rect 9781 30209 9815 30243
rect 13461 30209 13495 30243
rect 13550 30212 13584 30246
rect 13650 30209 13684 30243
rect 13829 30209 13863 30243
rect 15393 30209 15427 30243
rect 15669 30209 15703 30243
rect 15761 30209 15795 30243
rect 22017 30209 22051 30243
rect 23774 30209 23808 30243
rect 24041 30209 24075 30243
rect 25614 30209 25648 30243
rect 25881 30209 25915 30243
rect 14933 30141 14967 30175
rect 20913 30141 20947 30175
rect 5825 30073 5859 30107
rect 8033 30073 8067 30107
rect 14381 30073 14415 30107
rect 22661 30073 22695 30107
rect 1961 30005 1995 30039
rect 2421 30005 2455 30039
rect 15945 30005 15979 30039
rect 19533 30005 19567 30039
rect 22201 30005 22235 30039
rect 2605 29801 2639 29835
rect 10977 29801 11011 29835
rect 22569 29801 22603 29835
rect 1409 29733 1443 29767
rect 12081 29733 12115 29767
rect 14197 29665 14231 29699
rect 1961 29597 1995 29631
rect 2145 29597 2179 29631
rect 2237 29597 2271 29631
rect 2329 29597 2363 29631
rect 7297 29597 7331 29631
rect 7481 29597 7515 29631
rect 9597 29597 9631 29631
rect 12265 29597 12299 29631
rect 13185 29597 13219 29631
rect 13274 29597 13308 29631
rect 13369 29597 13403 29631
rect 13553 29597 13587 29631
rect 17233 29597 17267 29631
rect 17325 29597 17359 29631
rect 17601 29597 17635 29631
rect 18061 29597 18095 29631
rect 18209 29597 18243 29631
rect 18337 29597 18371 29631
rect 18526 29597 18560 29631
rect 19257 29597 19291 29631
rect 19405 29597 19439 29631
rect 19722 29597 19756 29631
rect 21925 29597 21959 29631
rect 22088 29597 22122 29631
rect 22188 29594 22222 29628
rect 22293 29597 22327 29631
rect 26985 29597 27019 29631
rect 68109 29597 68143 29631
rect 3801 29529 3835 29563
rect 3985 29529 4019 29563
rect 6193 29529 6227 29563
rect 8125 29529 8159 29563
rect 8309 29529 8343 29563
rect 9864 29529 9898 29563
rect 12449 29529 12483 29563
rect 17417 29529 17451 29563
rect 18429 29529 18463 29563
rect 19533 29529 19567 29563
rect 19625 29529 19659 29563
rect 20361 29529 20395 29563
rect 26718 29529 26752 29563
rect 4169 29461 4203 29495
rect 7113 29461 7147 29495
rect 7941 29461 7975 29495
rect 12909 29461 12943 29495
rect 16589 29461 16623 29495
rect 17049 29461 17083 29495
rect 18705 29461 18739 29495
rect 19901 29461 19935 29495
rect 25605 29461 25639 29495
rect 3065 29257 3099 29291
rect 7113 29257 7147 29291
rect 10241 29257 10275 29291
rect 11529 29257 11563 29291
rect 15393 29257 15427 29291
rect 15945 29257 15979 29291
rect 16865 29257 16899 29291
rect 14289 29189 14323 29223
rect 17233 29189 17267 29223
rect 27353 29189 27387 29223
rect 2421 29121 2455 29155
rect 2605 29121 2639 29155
rect 2697 29121 2731 29155
rect 2789 29121 2823 29155
rect 4077 29121 4111 29155
rect 4344 29121 4378 29155
rect 6469 29121 6503 29155
rect 6653 29121 6687 29155
rect 6745 29121 6779 29155
rect 6837 29121 6871 29155
rect 7757 29121 7791 29155
rect 8024 29121 8058 29155
rect 9597 29121 9631 29155
rect 9781 29121 9815 29155
rect 9873 29121 9907 29155
rect 9965 29121 9999 29155
rect 12653 29121 12687 29155
rect 15209 29121 15243 29155
rect 16037 29121 16071 29155
rect 17049 29121 17083 29155
rect 17141 29121 17175 29155
rect 17417 29121 17451 29155
rect 18981 29121 19015 29155
rect 19129 29121 19163 29155
rect 19257 29121 19291 29155
rect 19349 29121 19383 29155
rect 19446 29121 19480 29155
rect 24878 29121 24912 29155
rect 25145 29121 25179 29155
rect 29101 29121 29135 29155
rect 29561 29121 29595 29155
rect 12909 29053 12943 29087
rect 3617 28985 3651 29019
rect 5457 28985 5491 29019
rect 9137 28985 9171 29019
rect 19625 28985 19659 29019
rect 23765 28985 23799 29019
rect 17969 28917 18003 28951
rect 18429 28917 18463 28951
rect 4445 28713 4479 28747
rect 8125 28713 8159 28747
rect 6929 28577 6963 28611
rect 21465 28577 21499 28611
rect 23397 28577 23431 28611
rect 25789 28577 25823 28611
rect 1685 28509 1719 28543
rect 3801 28509 3835 28543
rect 3985 28509 4019 28543
rect 4077 28509 4111 28543
rect 4169 28509 4203 28543
rect 7481 28509 7515 28543
rect 7665 28509 7699 28543
rect 7757 28509 7791 28543
rect 7849 28509 7883 28543
rect 9965 28509 9999 28543
rect 13001 28509 13035 28543
rect 13369 28509 13403 28543
rect 14473 28509 14507 28543
rect 16773 28509 16807 28543
rect 16921 28509 16955 28543
rect 17141 28509 17175 28543
rect 17238 28509 17272 28543
rect 17877 28509 17911 28543
rect 29009 28509 29043 28543
rect 1869 28441 1903 28475
rect 10232 28441 10266 28475
rect 13185 28441 13219 28475
rect 13277 28441 13311 28475
rect 17049 28441 17083 28475
rect 21198 28441 21232 28475
rect 23130 28441 23164 28475
rect 26034 28441 26068 28475
rect 28742 28441 28776 28475
rect 2053 28373 2087 28407
rect 3249 28373 3283 28407
rect 6285 28373 6319 28407
rect 9413 28373 9447 28407
rect 11345 28373 11379 28407
rect 13553 28373 13587 28407
rect 15761 28373 15795 28407
rect 17417 28373 17451 28407
rect 20085 28373 20119 28407
rect 22017 28373 22051 28407
rect 27169 28373 27203 28407
rect 27629 28373 27663 28407
rect 10149 28169 10183 28203
rect 13093 28169 13127 28203
rect 20729 28169 20763 28203
rect 22017 28169 22051 28203
rect 25789 28169 25823 28203
rect 12817 28101 12851 28135
rect 19257 28101 19291 28135
rect 1869 28033 1903 28067
rect 2053 28033 2087 28067
rect 2145 28033 2179 28067
rect 2237 28033 2271 28067
rect 2973 28033 3007 28067
rect 7665 28033 7699 28067
rect 9505 28033 9539 28067
rect 9689 28033 9723 28067
rect 9781 28033 9815 28067
rect 9873 28033 9907 28067
rect 12541 28033 12575 28067
rect 12725 28033 12759 28067
rect 12909 28033 12943 28067
rect 15229 28033 15263 28067
rect 15485 28033 15519 28067
rect 18357 28033 18391 28067
rect 19441 28033 19475 28067
rect 19625 28033 19659 28067
rect 20085 28033 20119 28067
rect 20248 28036 20282 28070
rect 20348 28036 20382 28070
rect 20499 28033 20533 28067
rect 22293 28033 22327 28067
rect 22385 28033 22419 28067
rect 22477 28033 22511 28067
rect 22661 28033 22695 28067
rect 25145 28033 25179 28067
rect 25324 28033 25358 28067
rect 25424 28039 25458 28073
rect 25513 28033 25547 28067
rect 30398 28033 30432 28067
rect 30665 28033 30699 28067
rect 18613 27965 18647 27999
rect 21281 27965 21315 27999
rect 67649 27897 67683 27931
rect 2513 27829 2547 27863
rect 7205 27829 7239 27863
rect 13553 27829 13587 27863
rect 14105 27829 14139 27863
rect 15945 27829 15979 27863
rect 16681 27829 16715 27863
rect 17233 27829 17267 27863
rect 23213 27829 23247 27863
rect 26249 27829 26283 27863
rect 29285 27829 29319 27863
rect 10057 27625 10091 27659
rect 21465 27625 21499 27659
rect 25697 27625 25731 27659
rect 14105 27557 14139 27591
rect 23857 27557 23891 27591
rect 24593 27557 24627 27591
rect 28273 27557 28307 27591
rect 11069 27489 11103 27523
rect 16313 27489 16347 27523
rect 19349 27489 19383 27523
rect 20177 27489 20211 27523
rect 20453 27489 20487 27523
rect 22477 27489 22511 27523
rect 2237 27421 2271 27455
rect 3801 27421 3835 27455
rect 3985 27421 4019 27455
rect 4077 27421 4111 27455
rect 4169 27421 4203 27455
rect 5457 27421 5491 27455
rect 5713 27421 5747 27455
rect 7297 27421 7331 27455
rect 7481 27421 7515 27455
rect 7576 27415 7610 27449
rect 7665 27421 7699 27455
rect 9873 27421 9907 27455
rect 11336 27421 11370 27455
rect 13369 27421 13403 27455
rect 14381 27421 14415 27455
rect 14473 27421 14507 27455
rect 14565 27421 14599 27455
rect 14749 27421 14783 27455
rect 16037 27421 16071 27455
rect 16773 27421 16807 27455
rect 16921 27421 16955 27455
rect 17238 27421 17272 27455
rect 19257 27421 19291 27455
rect 19441 27421 19475 27455
rect 22109 27421 22143 27455
rect 22293 27421 22327 27455
rect 23213 27421 23247 27455
rect 23376 27421 23410 27455
rect 23476 27421 23510 27455
rect 23581 27421 23615 27455
rect 25053 27421 25087 27455
rect 25237 27421 25271 27455
rect 25329 27421 25363 27455
rect 25421 27421 25455 27455
rect 27629 27421 27663 27455
rect 27792 27421 27826 27455
rect 27892 27421 27926 27455
rect 27997 27421 28031 27455
rect 2881 27353 2915 27387
rect 3065 27353 3099 27387
rect 3249 27353 3283 27387
rect 9689 27353 9723 27387
rect 13553 27353 13587 27387
rect 17049 27353 17083 27387
rect 17141 27353 17175 27387
rect 17969 27353 18003 27387
rect 26157 27353 26191 27387
rect 26341 27353 26375 27387
rect 2053 27285 2087 27319
rect 4445 27285 4479 27319
rect 6837 27285 6871 27319
rect 7941 27285 7975 27319
rect 12449 27285 12483 27319
rect 13185 27285 13219 27319
rect 17417 27285 17451 27319
rect 18613 27285 18647 27319
rect 26525 27285 26559 27319
rect 27077 27285 27111 27319
rect 2145 27081 2179 27115
rect 5457 27081 5491 27115
rect 9413 27081 9447 27115
rect 12817 27081 12851 27115
rect 14657 27081 14691 27115
rect 15485 27081 15519 27115
rect 18981 27081 19015 27115
rect 21189 27081 21223 27115
rect 23489 27081 23523 27115
rect 25053 27081 25087 27115
rect 26341 27081 26375 27115
rect 27629 27081 27663 27115
rect 28457 27081 28491 27115
rect 4344 27013 4378 27047
rect 7840 27013 7874 27047
rect 12633 27013 12667 27047
rect 13461 27013 13495 27047
rect 17601 27013 17635 27047
rect 18337 27013 18371 27047
rect 18521 27013 18555 27047
rect 20177 27013 20211 27047
rect 23305 27013 23339 27047
rect 24685 27013 24719 27047
rect 2329 26945 2363 26979
rect 3341 26945 3375 26979
rect 6929 26945 6963 26979
rect 9597 26945 9631 26979
rect 9781 26945 9815 26979
rect 12449 26945 12483 26979
rect 13277 26945 13311 26979
rect 13553 26945 13587 26979
rect 13645 26945 13679 26979
rect 14841 26945 14875 26979
rect 15025 26945 15059 26979
rect 15761 26945 15795 26979
rect 15853 26945 15887 26979
rect 15945 26945 15979 26979
rect 16129 26945 16163 26979
rect 16681 26945 16715 26979
rect 16865 26945 16899 26979
rect 17509 26945 17543 26979
rect 17693 26945 17727 26979
rect 18153 26945 18187 26979
rect 19211 26945 19245 26979
rect 19349 26945 19383 26979
rect 19441 26945 19475 26979
rect 19625 26945 19659 26979
rect 20361 26945 20395 26979
rect 21005 26945 21039 26979
rect 23121 26945 23155 26979
rect 24869 26945 24903 26979
rect 26985 26945 27019 26979
rect 27148 26945 27182 26979
rect 27261 26945 27295 26979
rect 27353 26945 27387 26979
rect 28089 26945 28123 26979
rect 28273 26945 28307 26979
rect 3617 26877 3651 26911
rect 4077 26877 4111 26911
rect 7573 26877 7607 26911
rect 8953 26809 8987 26843
rect 13829 26809 13863 26843
rect 20545 26809 20579 26843
rect 7113 26741 7147 26775
rect 17049 26741 17083 26775
rect 67649 26741 67683 26775
rect 5825 26537 5859 26571
rect 26893 26537 26927 26571
rect 14657 26469 14691 26503
rect 17417 26469 17451 26503
rect 21373 26469 21407 26503
rect 2605 26401 2639 26435
rect 7021 26401 7055 26435
rect 19993 26401 20027 26435
rect 30389 26401 30423 26435
rect 2881 26333 2915 26367
rect 3893 26333 3927 26367
rect 4445 26333 4479 26367
rect 7297 26333 7331 26367
rect 7941 26333 7975 26367
rect 8125 26333 8159 26367
rect 11805 26333 11839 26367
rect 14105 26333 14139 26367
rect 14473 26333 14507 26367
rect 15485 26333 15519 26367
rect 15577 26333 15611 26367
rect 15669 26333 15703 26367
rect 15853 26333 15887 26367
rect 16773 26333 16807 26367
rect 16921 26333 16955 26367
rect 17049 26333 17083 26367
rect 17238 26333 17272 26367
rect 17877 26333 17911 26367
rect 18153 26333 18187 26367
rect 19441 26333 19475 26367
rect 20269 26333 20303 26367
rect 22753 26333 22787 26367
rect 26065 26333 26099 26367
rect 26709 26333 26743 26367
rect 4690 26265 4724 26299
rect 8953 26265 8987 26299
rect 11560 26265 11594 26299
rect 14289 26265 14323 26299
rect 14381 26265 14415 26299
rect 17141 26265 17175 26299
rect 22486 26265 22520 26299
rect 23489 26265 23523 26299
rect 23673 26265 23707 26299
rect 25798 26265 25832 26299
rect 26525 26265 26559 26299
rect 30656 26265 30690 26299
rect 7757 26197 7791 26231
rect 10425 26197 10459 26231
rect 15209 26197 15243 26231
rect 19257 26197 19291 26231
rect 23857 26197 23891 26231
rect 24685 26197 24719 26231
rect 31769 26197 31803 26231
rect 13185 25993 13219 26027
rect 18153 25993 18187 26027
rect 20821 25993 20855 26027
rect 22477 25993 22511 26027
rect 24869 25993 24903 26027
rect 26341 25993 26375 26027
rect 30757 25993 30791 26027
rect 2053 25925 2087 25959
rect 6745 25925 6779 25959
rect 12072 25925 12106 25959
rect 19533 25925 19567 25959
rect 27721 25925 27755 25959
rect 29294 25925 29328 25959
rect 31401 25925 31435 25959
rect 1869 25857 1903 25891
rect 3994 25857 4028 25891
rect 4261 25857 4295 25891
rect 8493 25857 8527 25891
rect 8953 25857 8987 25891
rect 9209 25857 9243 25891
rect 11805 25857 11839 25891
rect 14657 25857 14691 25891
rect 15577 25857 15611 25891
rect 16957 25857 16991 25891
rect 18705 25857 18739 25891
rect 18889 25857 18923 25891
rect 21833 25857 21867 25891
rect 22017 25857 22051 25891
rect 22109 25857 22143 25891
rect 22201 25857 22235 25891
rect 22937 25857 22971 25891
rect 24225 25857 24259 25891
rect 24388 25857 24422 25891
rect 24504 25857 24538 25891
rect 24613 25857 24647 25891
rect 27077 25857 27111 25891
rect 27261 25857 27295 25891
rect 27353 25857 27387 25891
rect 27445 25857 27479 25891
rect 29561 25857 29595 25891
rect 30113 25857 30147 25891
rect 30297 25857 30331 25891
rect 30392 25857 30426 25891
rect 30527 25857 30561 25891
rect 31217 25857 31251 25891
rect 15301 25789 15335 25823
rect 16681 25789 16715 25823
rect 2237 25653 2271 25687
rect 2881 25653 2915 25687
rect 10333 25653 10367 25687
rect 13645 25653 13679 25687
rect 14841 25653 14875 25687
rect 19073 25653 19107 25687
rect 23673 25653 23707 25687
rect 28181 25653 28215 25687
rect 31585 25653 31619 25687
rect 2973 25449 3007 25483
rect 6745 25449 6779 25483
rect 8401 25449 8435 25483
rect 12909 25449 12943 25483
rect 20637 25449 20671 25483
rect 27353 25449 27387 25483
rect 29929 25449 29963 25483
rect 18337 25381 18371 25415
rect 30389 25381 30423 25415
rect 1869 25313 1903 25347
rect 14105 25313 14139 25347
rect 1685 25245 1719 25279
rect 2329 25245 2363 25279
rect 2513 25245 2547 25279
rect 2605 25245 2639 25279
rect 2697 25245 2731 25279
rect 5365 25245 5399 25279
rect 7297 25245 7331 25279
rect 7757 25245 7791 25279
rect 7920 25245 7954 25279
rect 8020 25242 8054 25276
rect 8171 25245 8205 25279
rect 8953 25245 8987 25279
rect 9137 25245 9171 25279
rect 13165 25245 13199 25279
rect 13274 25245 13308 25279
rect 13374 25245 13408 25279
rect 13553 25245 13587 25279
rect 14381 25245 14415 25279
rect 17049 25245 17083 25279
rect 17142 25245 17176 25279
rect 17325 25245 17359 25279
rect 17533 25245 17567 25279
rect 18521 25245 18555 25279
rect 18613 25245 18647 25279
rect 19533 25245 19567 25279
rect 19717 25245 19751 25279
rect 19809 25245 19843 25279
rect 19901 25245 19935 25279
rect 22017 25245 22051 25279
rect 23857 25245 23891 25279
rect 25421 25245 25455 25279
rect 27169 25245 27203 25279
rect 30941 25245 30975 25279
rect 31125 25239 31159 25273
rect 31220 25245 31254 25279
rect 31309 25245 31343 25279
rect 33425 25245 33459 25279
rect 68109 25245 68143 25279
rect 1501 25177 1535 25211
rect 5632 25177 5666 25211
rect 17417 25177 17451 25211
rect 20177 25177 20211 25211
rect 21750 25177 21784 25211
rect 23590 25177 23624 25211
rect 25605 25177 25639 25211
rect 26985 25177 27019 25211
rect 31585 25177 31619 25211
rect 33158 25177 33192 25211
rect 3893 25109 3927 25143
rect 9321 25109 9355 25143
rect 9873 25109 9907 25143
rect 15945 25109 15979 25143
rect 17693 25109 17727 25143
rect 22477 25109 22511 25143
rect 25789 25109 25823 25143
rect 26341 25109 26375 25143
rect 32045 25109 32079 25143
rect 12633 24905 12667 24939
rect 23489 24905 23523 24939
rect 24961 24905 24995 24939
rect 31125 24905 31159 24939
rect 1409 24837 1443 24871
rect 1777 24837 1811 24871
rect 18061 24837 18095 24871
rect 30757 24837 30791 24871
rect 1593 24769 1627 24803
rect 2237 24769 2271 24803
rect 2421 24769 2455 24803
rect 2513 24769 2547 24803
rect 2651 24769 2685 24803
rect 3801 24769 3835 24803
rect 4068 24769 4102 24803
rect 7113 24769 7147 24803
rect 8493 24769 8527 24803
rect 8677 24769 8711 24803
rect 8769 24769 8803 24803
rect 8861 24769 8895 24803
rect 9853 24769 9887 24803
rect 12081 24769 12115 24803
rect 12265 24769 12299 24803
rect 12357 24769 12391 24803
rect 12449 24769 12483 24803
rect 13645 24769 13679 24803
rect 15862 24769 15896 24803
rect 16129 24769 16163 24803
rect 19726 24769 19760 24803
rect 19993 24769 20027 24803
rect 23765 24769 23799 24803
rect 23854 24769 23888 24803
rect 23954 24769 23988 24803
rect 24133 24769 24167 24803
rect 25053 24769 25087 24803
rect 25605 24769 25639 24803
rect 25789 24769 25823 24803
rect 25884 24769 25918 24803
rect 25973 24769 26007 24803
rect 28098 24769 28132 24803
rect 29101 24769 29135 24803
rect 29193 24769 29227 24803
rect 29285 24769 29319 24803
rect 29469 24769 29503 24803
rect 30113 24769 30147 24803
rect 30297 24769 30331 24803
rect 30941 24769 30975 24803
rect 2881 24701 2915 24735
rect 6837 24701 6871 24735
rect 9137 24701 9171 24735
rect 9597 24701 9631 24735
rect 13921 24701 13955 24735
rect 26249 24701 26283 24735
rect 28365 24701 28399 24735
rect 29929 24701 29963 24735
rect 5181 24565 5215 24599
rect 10977 24565 11011 24599
rect 14749 24565 14783 24599
rect 18613 24565 18647 24599
rect 20545 24565 20579 24599
rect 21833 24565 21867 24599
rect 26985 24565 27019 24599
rect 28825 24565 28859 24599
rect 3801 24361 3835 24395
rect 7021 24361 7055 24395
rect 8309 24361 8343 24395
rect 12725 24361 12759 24395
rect 13553 24361 13587 24395
rect 19257 24361 19291 24395
rect 23765 24361 23799 24395
rect 26801 24361 26835 24395
rect 30573 24361 30607 24395
rect 10793 24293 10827 24327
rect 21281 24293 21315 24327
rect 2973 24225 3007 24259
rect 3249 24225 3283 24259
rect 18429 24225 18463 24259
rect 22201 24225 22235 24259
rect 7277 24157 7311 24191
rect 7389 24157 7423 24191
rect 7486 24157 7520 24191
rect 7665 24157 7699 24191
rect 8125 24157 8159 24191
rect 9413 24157 9447 24191
rect 12541 24157 12575 24191
rect 14289 24157 14323 24191
rect 15485 24157 15519 24191
rect 15761 24157 15795 24191
rect 16681 24157 16715 24191
rect 16829 24157 16863 24191
rect 17049 24157 17083 24191
rect 17146 24157 17180 24191
rect 18245 24157 18279 24191
rect 19533 24157 19567 24191
rect 19625 24157 19659 24191
rect 19717 24157 19751 24191
rect 19901 24157 19935 24191
rect 22661 24157 22695 24191
rect 23581 24157 23615 24191
rect 27721 24157 27755 24191
rect 27905 24157 27939 24191
rect 27997 24157 28031 24191
rect 28089 24157 28123 24191
rect 31125 24157 31159 24191
rect 31288 24157 31322 24191
rect 31401 24157 31435 24191
rect 31539 24157 31573 24191
rect 33977 24157 34011 24191
rect 68109 24157 68143 24191
rect 1593 24089 1627 24123
rect 1777 24089 1811 24123
rect 4353 24089 4387 24123
rect 6285 24089 6319 24123
rect 9658 24089 9692 24123
rect 12357 24089 12391 24123
rect 16957 24089 16991 24123
rect 18061 24089 18095 24123
rect 20545 24089 20579 24123
rect 21097 24089 21131 24123
rect 22017 24089 22051 24123
rect 23397 24089 23431 24123
rect 25513 24089 25547 24123
rect 31769 24089 31803 24123
rect 33710 24089 33744 24123
rect 1961 24021 1995 24055
rect 5733 24021 5767 24055
rect 6377 24021 6411 24055
rect 14381 24021 14415 24055
rect 17325 24021 17359 24055
rect 22845 24021 22879 24055
rect 24777 24021 24811 24055
rect 28365 24021 28399 24055
rect 32597 24021 32631 24055
rect 3709 23817 3743 23851
rect 5457 23817 5491 23851
rect 8861 23817 8895 23851
rect 9321 23817 9355 23851
rect 15485 23817 15519 23851
rect 27353 23817 27387 23851
rect 27905 23817 27939 23851
rect 31309 23817 31343 23851
rect 4261 23749 4295 23783
rect 17509 23749 17543 23783
rect 19441 23749 19475 23783
rect 27169 23749 27203 23783
rect 28816 23749 28850 23783
rect 3065 23681 3099 23715
rect 3249 23681 3283 23715
rect 3341 23681 3375 23715
rect 3479 23681 3513 23715
rect 5641 23681 5675 23715
rect 6929 23681 6963 23715
rect 8217 23681 8251 23715
rect 8401 23681 8435 23715
rect 8493 23681 8527 23715
rect 8585 23681 8619 23715
rect 12449 23681 12483 23715
rect 12633 23681 12667 23715
rect 13553 23681 13587 23715
rect 13645 23681 13679 23715
rect 13737 23681 13771 23715
rect 13921 23681 13955 23715
rect 14841 23681 14875 23715
rect 15025 23681 15059 23715
rect 15117 23681 15151 23715
rect 15209 23681 15243 23715
rect 17141 23681 17175 23715
rect 17289 23681 17323 23715
rect 17417 23681 17451 23715
rect 17606 23681 17640 23715
rect 19257 23681 19291 23715
rect 22109 23681 22143 23715
rect 23581 23681 23615 23715
rect 24593 23681 24627 23715
rect 26985 23681 27019 23715
rect 30941 23681 30975 23715
rect 31125 23681 31159 23715
rect 2329 23613 2363 23647
rect 2605 23613 2639 23647
rect 4997 23613 5031 23647
rect 5825 23613 5859 23647
rect 7205 23613 7239 23647
rect 12817 23613 12851 23647
rect 16037 23613 16071 23647
rect 18797 23613 18831 23647
rect 19625 23613 19659 23647
rect 23305 23613 23339 23647
rect 24869 23613 24903 23647
rect 25329 23613 25363 23647
rect 25605 23613 25639 23647
rect 28549 23613 28583 23647
rect 6377 23545 6411 23579
rect 17785 23545 17819 23579
rect 21189 23545 21223 23579
rect 13277 23477 13311 23511
rect 22201 23477 22235 23511
rect 29929 23477 29963 23511
rect 30481 23477 30515 23511
rect 1685 23273 1719 23307
rect 6653 23273 6687 23307
rect 7205 23273 7239 23307
rect 8401 23273 8435 23307
rect 13001 23273 13035 23307
rect 14657 23273 14691 23307
rect 15669 23273 15703 23307
rect 21925 23273 21959 23307
rect 25605 23273 25639 23307
rect 5641 23205 5675 23239
rect 13553 23205 13587 23239
rect 9781 23137 9815 23171
rect 17325 23137 17359 23171
rect 26985 23137 27019 23171
rect 27629 23137 27663 23171
rect 29837 23137 29871 23171
rect 1869 23069 1903 23103
rect 2329 23069 2363 23103
rect 2492 23069 2526 23103
rect 2605 23069 2639 23103
rect 2697 23069 2731 23103
rect 3801 23069 3835 23103
rect 6561 23069 6595 23103
rect 6745 23069 6779 23103
rect 7389 23069 7423 23103
rect 7573 23069 7607 23103
rect 8033 23069 8067 23103
rect 8953 23069 8987 23103
rect 11621 23069 11655 23103
rect 14473 23069 14507 23103
rect 15117 23069 15151 23103
rect 15485 23069 15519 23103
rect 17601 23069 17635 23103
rect 19441 23069 19475 23103
rect 19625 23069 19659 23103
rect 19717 23069 19751 23103
rect 19809 23069 19843 23103
rect 20545 23069 20579 23103
rect 22661 23069 22695 23103
rect 22845 23069 22879 23103
rect 22937 23069 22971 23103
rect 23029 23069 23063 23103
rect 26729 23069 26763 23103
rect 29561 23069 29595 23103
rect 30849 23069 30883 23103
rect 31585 23069 31619 23103
rect 2973 23001 3007 23035
rect 4046 23001 4080 23035
rect 5825 23001 5859 23035
rect 8217 23001 8251 23035
rect 9137 23001 9171 23035
rect 10026 23001 10060 23035
rect 11888 23001 11922 23035
rect 14289 23001 14323 23035
rect 15301 23001 15335 23035
rect 15393 23001 15427 23035
rect 18613 23001 18647 23035
rect 20790 23001 20824 23035
rect 27896 23001 27930 23035
rect 31830 23001 31864 23035
rect 5181 22933 5215 22967
rect 9321 22933 9355 22967
rect 11161 22933 11195 22967
rect 16221 22933 16255 22967
rect 20085 22933 20119 22967
rect 23305 22933 23339 22967
rect 23765 22933 23799 22967
rect 29009 22933 29043 22967
rect 31033 22933 31067 22967
rect 32965 22933 32999 22967
rect 9505 22729 9539 22763
rect 14197 22729 14231 22763
rect 26157 22729 26191 22763
rect 28089 22729 28123 22763
rect 30849 22729 30883 22763
rect 2421 22661 2455 22695
rect 3126 22661 3160 22695
rect 13829 22661 13863 22695
rect 13921 22661 13955 22695
rect 15025 22661 15059 22695
rect 17816 22661 17850 22695
rect 18613 22661 18647 22695
rect 24326 22661 24360 22695
rect 25329 22661 25363 22695
rect 29193 22661 29227 22695
rect 1777 22593 1811 22627
rect 1961 22593 1995 22627
rect 2053 22593 2087 22627
rect 2191 22593 2225 22627
rect 2881 22593 2915 22627
rect 4997 22593 5031 22627
rect 5089 22593 5123 22627
rect 5181 22593 5215 22627
rect 5365 22593 5399 22627
rect 7113 22593 7147 22627
rect 7205 22593 7239 22627
rect 7297 22593 7331 22627
rect 7481 22593 7515 22627
rect 8125 22593 8159 22627
rect 8309 22593 8343 22627
rect 8861 22593 8895 22627
rect 9045 22593 9079 22627
rect 9137 22593 9171 22627
rect 9229 22593 9263 22627
rect 9965 22593 9999 22627
rect 13645 22593 13679 22627
rect 14013 22593 14047 22627
rect 14657 22593 14691 22627
rect 14750 22593 14784 22627
rect 14933 22593 14967 22627
rect 15163 22593 15197 22627
rect 15853 22593 15887 22627
rect 18889 22593 18923 22627
rect 18981 22593 19015 22627
rect 19073 22593 19107 22627
rect 19257 22593 19291 22627
rect 20729 22593 20763 22627
rect 25513 22593 25547 22627
rect 26249 22593 26283 22627
rect 27445 22593 27479 22627
rect 27629 22593 27663 22627
rect 27721 22593 27755 22627
rect 27813 22593 27847 22627
rect 29377 22593 29411 22627
rect 30205 22593 30239 22627
rect 30389 22593 30423 22627
rect 30481 22593 30515 22627
rect 30619 22593 30653 22627
rect 31493 22593 31527 22627
rect 32137 22593 32171 22627
rect 7941 22525 7975 22559
rect 18061 22525 18095 22559
rect 21005 22525 21039 22559
rect 21833 22525 21867 22559
rect 22109 22525 22143 22559
rect 24593 22525 24627 22559
rect 29009 22525 29043 22559
rect 4261 22457 4295 22491
rect 31309 22457 31343 22491
rect 67649 22457 67683 22491
rect 4721 22389 4755 22423
rect 6837 22389 6871 22423
rect 15301 22389 15335 22423
rect 15945 22389 15979 22423
rect 16681 22389 16715 22423
rect 23213 22389 23247 22423
rect 2053 22185 2087 22219
rect 5089 22185 5123 22219
rect 18705 22185 18739 22219
rect 22753 22185 22787 22219
rect 23305 22185 23339 22219
rect 27629 22185 27663 22219
rect 30389 22185 30423 22219
rect 3065 22049 3099 22083
rect 7297 22049 7331 22083
rect 21649 22049 21683 22083
rect 26249 22049 26283 22083
rect 30941 22049 30975 22083
rect 1685 21981 1719 22015
rect 1869 21981 1903 22015
rect 5457 21981 5491 22015
rect 7021 21981 7055 22015
rect 14933 21981 14967 22015
rect 15209 21981 15243 22015
rect 15301 21981 15335 22015
rect 16313 21981 16347 22015
rect 16461 21981 16495 22015
rect 16681 21981 16715 22015
rect 16778 21981 16812 22015
rect 17417 21981 17451 22015
rect 18337 21981 18371 22015
rect 18521 21981 18555 22015
rect 20637 21981 20671 22015
rect 21925 21981 21959 22015
rect 22385 21981 22419 22015
rect 23213 21981 23247 22015
rect 23397 21981 23431 22015
rect 26525 21981 26559 22015
rect 30021 21981 30055 22015
rect 34161 21981 34195 22015
rect 5273 21913 5307 21947
rect 9137 21913 9171 21947
rect 9321 21913 9355 21947
rect 9873 21913 9907 21947
rect 10057 21913 10091 21947
rect 15117 21913 15151 21947
rect 16589 21913 16623 21947
rect 22569 21913 22603 21947
rect 25605 21913 25639 21947
rect 25789 21913 25823 21947
rect 30205 21913 30239 21947
rect 31208 21913 31242 21947
rect 33894 21913 33928 21947
rect 36369 21913 36403 21947
rect 2513 21845 2547 21879
rect 3985 21845 4019 21879
rect 6009 21845 6043 21879
rect 7757 21845 7791 21879
rect 8953 21845 8987 21879
rect 10241 21845 10275 21879
rect 14381 21845 14415 21879
rect 15485 21845 15519 21879
rect 16957 21845 16991 21879
rect 19349 21845 19383 21879
rect 25053 21845 25087 21879
rect 32321 21845 32355 21879
rect 32781 21845 32815 21879
rect 35909 21845 35943 21879
rect 37657 21845 37691 21879
rect 2973 21641 3007 21675
rect 6377 21641 6411 21675
rect 7113 21641 7147 21675
rect 13829 21641 13863 21675
rect 16773 21641 16807 21675
rect 17969 21641 18003 21675
rect 21281 21641 21315 21675
rect 28641 21641 28675 21675
rect 31125 21641 31159 21675
rect 4712 21573 4746 21607
rect 11621 21573 11655 21607
rect 11805 21573 11839 21607
rect 23581 21573 23615 21607
rect 24317 21573 24351 21607
rect 25513 21573 25547 21607
rect 33149 21573 33183 21607
rect 3157 21505 3191 21539
rect 3709 21505 3743 21539
rect 4445 21505 4479 21539
rect 6377 21505 6411 21539
rect 6561 21505 6595 21539
rect 7921 21505 7955 21539
rect 9853 21505 9887 21539
rect 12449 21505 12483 21539
rect 12716 21505 12750 21539
rect 15577 21505 15611 21539
rect 16957 21505 16991 21539
rect 17877 21505 17911 21539
rect 19818 21505 19852 21539
rect 20085 21505 20119 21539
rect 21097 21505 21131 21539
rect 22661 21505 22695 21539
rect 23305 21505 23339 21539
rect 23489 21505 23523 21539
rect 23673 21505 23707 21539
rect 25145 21505 25179 21539
rect 25293 21505 25327 21539
rect 25421 21505 25455 21539
rect 25610 21505 25644 21539
rect 26433 21505 26467 21539
rect 27261 21505 27295 21539
rect 27353 21505 27387 21539
rect 27445 21505 27479 21539
rect 27629 21505 27663 21539
rect 28549 21505 28583 21539
rect 28733 21505 28767 21539
rect 29193 21505 29227 21539
rect 30481 21505 30515 21539
rect 30665 21505 30699 21539
rect 30757 21505 30791 21539
rect 30849 21505 30883 21539
rect 32965 21505 32999 21539
rect 34529 21505 34563 21539
rect 34713 21505 34747 21539
rect 36470 21505 36504 21539
rect 36737 21505 36771 21539
rect 7665 21437 7699 21471
rect 9597 21437 9631 21471
rect 20913 21437 20947 21471
rect 22385 21437 22419 21471
rect 29469 21437 29503 21471
rect 5825 21369 5859 21403
rect 10977 21369 11011 21403
rect 23857 21369 23891 21403
rect 35357 21369 35391 21403
rect 2053 21301 2087 21335
rect 3801 21301 3835 21335
rect 9045 21301 9079 21335
rect 11989 21301 12023 21335
rect 18705 21301 18739 21335
rect 25789 21301 25823 21335
rect 26985 21301 27019 21335
rect 33333 21301 33367 21335
rect 34897 21301 34931 21335
rect 67649 21301 67683 21335
rect 8033 21097 8067 21131
rect 9597 21097 9631 21131
rect 12357 21097 12391 21131
rect 16589 21097 16623 21131
rect 19901 21097 19935 21131
rect 21649 21097 21683 21131
rect 22661 21097 22695 21131
rect 29009 21097 29043 21131
rect 30389 21097 30423 21131
rect 33609 21097 33643 21131
rect 35633 21097 35667 21131
rect 9045 21029 9079 21063
rect 17049 21029 17083 21063
rect 23765 21029 23799 21063
rect 34161 21029 34195 21063
rect 6193 20961 6227 20995
rect 6653 20961 6687 20995
rect 18705 20961 18739 20995
rect 26801 20961 26835 20995
rect 28641 20961 28675 20995
rect 32413 20961 32447 20995
rect 38025 20961 38059 20995
rect 2329 20893 2363 20927
rect 2605 20893 2639 20927
rect 9827 20893 9861 20927
rect 9965 20893 9999 20927
rect 10057 20893 10091 20927
rect 10241 20893 10275 20927
rect 11713 20893 11747 20927
rect 11897 20893 11931 20927
rect 11992 20893 12026 20927
rect 12081 20893 12115 20927
rect 15485 20893 15519 20927
rect 19257 20893 19291 20927
rect 19441 20893 19475 20927
rect 19533 20893 19567 20927
rect 19625 20893 19659 20927
rect 21097 20893 21131 20927
rect 22569 20893 22603 20927
rect 22753 20893 22787 20927
rect 23213 20893 23247 20927
rect 23489 20893 23523 20927
rect 23581 20893 23615 20927
rect 24409 20893 24443 20927
rect 25140 20893 25174 20927
rect 25329 20893 25363 20927
rect 25512 20893 25546 20927
rect 25605 20893 25639 20927
rect 27068 20893 27102 20927
rect 28825 20893 28859 20927
rect 30021 20893 30055 20927
rect 32965 20893 32999 20927
rect 33149 20893 33183 20927
rect 33241 20893 33275 20927
rect 33333 20893 33367 20927
rect 34989 20893 35023 20927
rect 35173 20893 35207 20927
rect 35265 20893 35299 20927
rect 35357 20893 35391 20927
rect 3985 20825 4019 20859
rect 4445 20825 4479 20859
rect 6920 20825 6954 20859
rect 11161 20825 11195 20859
rect 15240 20825 15274 20859
rect 17601 20825 17635 20859
rect 18337 20825 18371 20859
rect 18521 20825 18555 20859
rect 21741 20825 21775 20859
rect 23397 20825 23431 20859
rect 25237 20825 25271 20859
rect 30205 20825 30239 20859
rect 37758 20825 37792 20859
rect 3249 20757 3283 20791
rect 14105 20757 14139 20791
rect 20453 20757 20487 20791
rect 20913 20757 20947 20791
rect 24961 20757 24995 20791
rect 28181 20757 28215 20791
rect 30849 20757 30883 20791
rect 31953 20757 31987 20791
rect 36093 20757 36127 20791
rect 36645 20757 36679 20791
rect 7297 20553 7331 20587
rect 7757 20553 7791 20587
rect 10977 20553 11011 20587
rect 15485 20553 15519 20587
rect 27721 20553 27755 20587
rect 28549 20553 28583 20587
rect 35725 20553 35759 20587
rect 4813 20485 4847 20519
rect 6377 20485 6411 20519
rect 11529 20485 11563 20519
rect 11713 20485 11747 20519
rect 12694 20485 12728 20519
rect 17785 20485 17819 20519
rect 18153 20485 18187 20519
rect 23489 20485 23523 20519
rect 23581 20485 23615 20519
rect 25605 20485 25639 20519
rect 30941 20485 30975 20519
rect 34161 20485 34195 20519
rect 34345 20485 34379 20519
rect 1961 20417 1995 20451
rect 2145 20417 2179 20451
rect 3056 20417 3090 20451
rect 4629 20417 4663 20451
rect 7113 20417 7147 20451
rect 8033 20417 8067 20451
rect 8125 20417 8159 20451
rect 8217 20417 8251 20451
rect 8401 20417 8435 20451
rect 10333 20417 10367 20451
rect 10496 20420 10530 20454
rect 10609 20417 10643 20451
rect 10747 20417 10781 20451
rect 11897 20417 11931 20451
rect 15761 20417 15795 20451
rect 15853 20417 15887 20451
rect 15945 20417 15979 20451
rect 16141 20417 16175 20451
rect 16957 20417 16991 20451
rect 17049 20417 17083 20451
rect 17141 20417 17175 20451
rect 17325 20417 17359 20451
rect 17969 20417 18003 20451
rect 20729 20417 20763 20451
rect 23305 20417 23339 20451
rect 23673 20417 23707 20451
rect 25467 20417 25501 20451
rect 25697 20417 25731 20451
rect 25825 20417 25859 20451
rect 25973 20417 26007 20451
rect 27905 20417 27939 20451
rect 28089 20417 28123 20451
rect 29285 20417 29319 20451
rect 31493 20417 31527 20451
rect 33250 20417 33284 20451
rect 33977 20417 34011 20451
rect 35081 20417 35115 20451
rect 35265 20417 35299 20451
rect 35357 20417 35391 20451
rect 35449 20417 35483 20451
rect 36185 20417 36219 20451
rect 38209 20417 38243 20451
rect 38465 20417 38499 20451
rect 2796 20349 2830 20383
rect 6929 20349 6963 20383
rect 12449 20349 12483 20383
rect 20453 20349 20487 20383
rect 33517 20349 33551 20383
rect 4169 20281 4203 20315
rect 5825 20281 5859 20315
rect 8861 20281 8895 20315
rect 13829 20281 13863 20315
rect 22753 20281 22787 20315
rect 23857 20281 23891 20315
rect 37473 20281 37507 20315
rect 1777 20213 1811 20247
rect 4997 20213 5031 20247
rect 9413 20213 9447 20247
rect 16681 20213 16715 20247
rect 19073 20213 19107 20247
rect 19901 20213 19935 20247
rect 21833 20213 21867 20247
rect 25329 20213 25363 20247
rect 32137 20213 32171 20247
rect 39589 20213 39623 20247
rect 2513 20009 2547 20043
rect 13093 20009 13127 20043
rect 15577 20009 15611 20043
rect 19257 20009 19291 20043
rect 31769 20009 31803 20043
rect 10609 19941 10643 19975
rect 27813 19941 27847 19975
rect 29745 19941 29779 19975
rect 35633 19941 35667 19975
rect 2973 19873 3007 19907
rect 5457 19873 5491 19907
rect 16865 19873 16899 19907
rect 22753 19873 22787 19907
rect 1869 19805 1903 19839
rect 2053 19805 2087 19839
rect 2145 19805 2179 19839
rect 2237 19805 2271 19839
rect 4353 19805 4387 19839
rect 4537 19805 4571 19839
rect 4629 19805 4663 19839
rect 4721 19805 4755 19839
rect 9229 19805 9263 19839
rect 11345 19805 11379 19839
rect 11805 19805 11839 19839
rect 15393 19805 15427 19839
rect 16221 19805 16255 19839
rect 17121 19805 17155 19839
rect 19441 19805 19475 19839
rect 19533 19805 19567 19839
rect 19809 19805 19843 19839
rect 20269 19805 20303 19839
rect 20453 19805 20487 19839
rect 20545 19805 20579 19839
rect 20637 19805 20671 19839
rect 23213 19805 23247 19839
rect 23397 19805 23431 19839
rect 23489 19805 23523 19839
rect 23581 19805 23615 19839
rect 24409 19805 24443 19839
rect 25232 19805 25266 19839
rect 25421 19805 25455 19839
rect 25604 19805 25638 19839
rect 25697 19805 25731 19839
rect 26433 19805 26467 19839
rect 26617 19805 26651 19839
rect 26709 19805 26743 19839
rect 26801 19805 26835 19839
rect 28365 19805 28399 19839
rect 28549 19805 28583 19839
rect 28641 19805 28675 19839
rect 28733 19805 28767 19839
rect 29561 19805 29595 19839
rect 30297 19805 30331 19839
rect 31125 19805 31159 19839
rect 31309 19805 31343 19839
rect 31401 19805 31435 19839
rect 31539 19805 31573 19839
rect 32229 19805 32263 19839
rect 34897 19805 34931 19839
rect 37013 19805 37047 19839
rect 68109 19805 68143 19839
rect 4997 19737 5031 19771
rect 5702 19737 5736 19771
rect 7389 19737 7423 19771
rect 7573 19737 7607 19771
rect 8033 19737 8067 19771
rect 8217 19737 8251 19771
rect 9474 19737 9508 19771
rect 15209 19737 15243 19771
rect 19625 19737 19659 19771
rect 20913 19737 20947 19771
rect 22486 19737 22520 19771
rect 23857 19737 23891 19771
rect 25329 19737 25363 19771
rect 30481 19737 30515 19771
rect 30665 19737 30699 19771
rect 34713 19737 34747 19771
rect 36746 19737 36780 19771
rect 37473 19737 37507 19771
rect 37657 19737 37691 19771
rect 6837 19669 6871 19703
rect 8401 19669 8435 19703
rect 18245 19669 18279 19703
rect 21373 19669 21407 19703
rect 24593 19669 24627 19703
rect 25053 19669 25087 19703
rect 27077 19669 27111 19703
rect 29009 19669 29043 19703
rect 34161 19669 34195 19703
rect 35081 19669 35115 19703
rect 37841 19669 37875 19703
rect 1685 19465 1719 19499
rect 9137 19465 9171 19499
rect 16773 19465 16807 19499
rect 22983 19465 23017 19499
rect 26249 19465 26283 19499
rect 30481 19465 30515 19499
rect 35817 19465 35851 19499
rect 38209 19465 38243 19499
rect 2789 19397 2823 19431
rect 3678 19397 3712 19431
rect 14933 19397 14967 19431
rect 19257 19397 19291 19431
rect 20361 19397 20395 19431
rect 31309 19397 31343 19431
rect 2145 19329 2179 19363
rect 2329 19329 2363 19363
rect 2421 19329 2455 19363
rect 2513 19329 2547 19363
rect 3433 19329 3467 19363
rect 7297 19329 7331 19363
rect 8493 19329 8527 19363
rect 8656 19329 8690 19363
rect 8769 19329 8803 19363
rect 8907 19329 8941 19363
rect 12357 19329 12391 19363
rect 14749 19329 14783 19363
rect 15669 19329 15703 19363
rect 15761 19329 15795 19363
rect 15853 19332 15887 19366
rect 16037 19329 16071 19363
rect 18981 19329 19015 19363
rect 19165 19329 19199 19363
rect 19349 19329 19383 19363
rect 20545 19329 20579 19363
rect 24685 19329 24719 19363
rect 26985 19329 27019 19363
rect 27241 19329 27275 19363
rect 29101 19329 29135 19363
rect 29357 19329 29391 19363
rect 34446 19329 34480 19363
rect 35173 19329 35207 19363
rect 35357 19329 35391 19363
rect 35449 19329 35483 19363
rect 35541 19329 35575 19363
rect 37565 19329 37599 19363
rect 37749 19329 37783 19363
rect 37841 19329 37875 19363
rect 37933 19329 37967 19363
rect 39385 19329 39419 19363
rect 6561 19261 6595 19295
rect 7021 19261 7055 19295
rect 9689 19261 9723 19295
rect 12633 19261 12667 19295
rect 14565 19261 14599 19295
rect 17325 19261 17359 19295
rect 20729 19261 20763 19295
rect 21189 19261 21223 19295
rect 22753 19261 22787 19295
rect 24961 19261 24995 19295
rect 34713 19261 34747 19295
rect 39129 19261 39163 19295
rect 10241 19193 10275 19227
rect 31493 19193 31527 19227
rect 4813 19125 4847 19159
rect 13093 19125 13127 19159
rect 15393 19125 15427 19159
rect 19533 19125 19567 19159
rect 22293 19125 22327 19159
rect 28365 19125 28399 19159
rect 33333 19125 33367 19159
rect 36277 19125 36311 19159
rect 40509 19125 40543 19159
rect 2513 18921 2547 18955
rect 3065 18921 3099 18955
rect 21005 18921 21039 18955
rect 27353 18921 27387 18955
rect 29561 18921 29595 18955
rect 39221 18921 39255 18955
rect 35081 18853 35115 18887
rect 6653 18785 6687 18819
rect 7481 18785 7515 18819
rect 8953 18785 8987 18819
rect 19533 18785 19567 18819
rect 22845 18785 22879 18819
rect 25973 18785 26007 18819
rect 28917 18785 28951 18819
rect 32321 18785 32355 18819
rect 38117 18785 38151 18819
rect 2145 18717 2179 18751
rect 6377 18717 6411 18751
rect 7389 18717 7423 18751
rect 7573 18717 7607 18751
rect 8033 18717 8067 18751
rect 8217 18717 8251 18751
rect 9229 18717 9263 18751
rect 10241 18717 10275 18751
rect 10977 18717 11011 18751
rect 15485 18717 15519 18751
rect 16405 18717 16439 18751
rect 16681 18717 16715 18751
rect 16773 18717 16807 18751
rect 17509 18717 17543 18751
rect 18153 18717 18187 18751
rect 18337 18717 18371 18751
rect 18429 18717 18463 18751
rect 18521 18717 18555 18751
rect 19257 18717 19291 18751
rect 20637 18717 20671 18751
rect 20821 18717 20855 18751
rect 21741 18717 21775 18751
rect 21833 18717 21867 18751
rect 21925 18717 21959 18751
rect 22109 18717 22143 18751
rect 22569 18717 22603 18751
rect 25706 18717 25740 18751
rect 27537 18717 27571 18751
rect 28825 18717 28859 18751
rect 29009 18717 29043 18751
rect 29745 18717 29779 18751
rect 33149 18717 33183 18751
rect 33425 18717 33459 18751
rect 38577 18717 38611 18751
rect 38756 18717 38790 18751
rect 38853 18717 38887 18751
rect 38945 18717 38979 18751
rect 39865 18717 39899 18751
rect 68109 18717 68143 18751
rect 2329 18649 2363 18683
rect 5365 18649 5399 18683
rect 8401 18649 8435 18683
rect 11244 18649 11278 18683
rect 12817 18649 12851 18683
rect 13001 18649 13035 18683
rect 15240 18649 15274 18683
rect 16589 18649 16623 18683
rect 21465 18649 21499 18683
rect 27721 18649 27755 18683
rect 29929 18649 29963 18683
rect 30481 18649 30515 18683
rect 32054 18649 32088 18683
rect 36369 18649 36403 18683
rect 10425 18581 10459 18615
rect 12357 18581 12391 18615
rect 13185 18581 13219 18615
rect 14105 18581 14139 18615
rect 16957 18581 16991 18615
rect 17601 18581 17635 18615
rect 18705 18581 18739 18615
rect 24593 18581 24627 18615
rect 28365 18581 28399 18615
rect 30941 18581 30975 18615
rect 35909 18581 35943 18615
rect 8217 18377 8251 18411
rect 11529 18377 11563 18411
rect 14105 18377 14139 18411
rect 22201 18377 22235 18411
rect 27721 18377 27755 18411
rect 38117 18377 38151 18411
rect 2513 18309 2547 18343
rect 8861 18309 8895 18343
rect 9045 18309 9079 18343
rect 15853 18309 15887 18343
rect 20269 18309 20303 18343
rect 22017 18309 22051 18343
rect 24142 18309 24176 18343
rect 30849 18309 30883 18343
rect 34253 18309 34287 18343
rect 37749 18309 37783 18343
rect 1869 18241 1903 18275
rect 2048 18241 2082 18275
rect 2145 18241 2179 18275
rect 2283 18241 2317 18275
rect 2973 18241 3007 18275
rect 3229 18241 3263 18275
rect 7490 18241 7524 18275
rect 7757 18241 7791 18275
rect 8401 18241 8435 18275
rect 9689 18241 9723 18275
rect 11805 18241 11839 18275
rect 11897 18241 11931 18275
rect 11989 18241 12023 18275
rect 12173 18241 12207 18275
rect 12981 18241 13015 18275
rect 16037 18241 16071 18275
rect 17187 18241 17221 18275
rect 17325 18241 17359 18275
rect 17417 18241 17451 18275
rect 17600 18241 17634 18275
rect 17693 18241 17727 18275
rect 18705 18241 18739 18275
rect 20131 18241 20165 18275
rect 20361 18241 20395 18275
rect 20544 18241 20578 18275
rect 20637 18241 20671 18275
rect 21281 18241 21315 18275
rect 21833 18241 21867 18275
rect 26341 18241 26375 18275
rect 29009 18241 29043 18275
rect 29653 18241 29687 18275
rect 29837 18241 29871 18275
rect 31033 18241 31067 18275
rect 32137 18241 32171 18275
rect 34437 18241 34471 18275
rect 35357 18241 35391 18275
rect 35613 18241 35647 18275
rect 37933 18241 37967 18275
rect 39293 18241 39327 18275
rect 9965 18173 9999 18207
rect 12725 18173 12759 18207
rect 18429 18173 18463 18207
rect 24409 18173 24443 18207
rect 26065 18173 26099 18207
rect 28273 18173 28307 18207
rect 28825 18173 28859 18207
rect 29745 18173 29779 18207
rect 32781 18173 32815 18207
rect 33057 18173 33091 18207
rect 39037 18173 39071 18207
rect 23029 18105 23063 18139
rect 29193 18105 29227 18139
rect 32321 18105 32355 18139
rect 4353 18037 4387 18071
rect 6377 18037 6411 18071
rect 9229 18037 9263 18071
rect 17049 18037 17083 18071
rect 19993 18037 20027 18071
rect 21097 18037 21131 18071
rect 30389 18037 30423 18071
rect 31217 18037 31251 18071
rect 34069 18037 34103 18071
rect 36737 18037 36771 18071
rect 40417 18037 40451 18071
rect 2697 17833 2731 17867
rect 10057 17833 10091 17867
rect 24777 17833 24811 17867
rect 33885 17833 33919 17867
rect 35357 17833 35391 17867
rect 37289 17833 37323 17867
rect 38485 17833 38519 17867
rect 4169 17697 4203 17731
rect 7021 17697 7055 17731
rect 14565 17697 14599 17731
rect 27905 17697 27939 17731
rect 29653 17697 29687 17731
rect 30941 17697 30975 17731
rect 32781 17697 32815 17731
rect 4353 17629 4387 17663
rect 7297 17629 7331 17663
rect 9413 17629 9447 17663
rect 9597 17626 9631 17660
rect 9689 17629 9723 17663
rect 9827 17629 9861 17663
rect 13001 17629 13035 17663
rect 16865 17629 16899 17663
rect 16954 17629 16988 17663
rect 17049 17629 17083 17663
rect 17233 17629 17267 17663
rect 18153 17629 18187 17663
rect 18337 17629 18371 17663
rect 18521 17629 18555 17663
rect 19533 17629 19567 17663
rect 20315 17629 20349 17663
rect 20453 17629 20487 17663
rect 20728 17629 20762 17663
rect 20821 17629 20855 17663
rect 24593 17629 24627 17663
rect 29009 17629 29043 17663
rect 29929 17629 29963 17663
rect 31125 17629 31159 17663
rect 31309 17629 31343 17663
rect 32505 17629 32539 17663
rect 33241 17629 33275 17663
rect 33425 17629 33459 17663
rect 33517 17629 33551 17663
rect 33655 17629 33689 17663
rect 35633 17629 35667 17663
rect 35725 17629 35759 17663
rect 35817 17629 35851 17663
rect 36001 17629 36035 17663
rect 36829 17629 36863 17663
rect 37841 17629 37875 17663
rect 38025 17629 38059 17663
rect 38120 17629 38154 17663
rect 38209 17629 38243 17663
rect 39129 17629 39163 17663
rect 4537 17561 4571 17595
rect 8309 17561 8343 17595
rect 12817 17561 12851 17595
rect 14832 17561 14866 17595
rect 16589 17561 16623 17595
rect 18429 17561 18463 17595
rect 19349 17561 19383 17595
rect 19717 17561 19751 17595
rect 20545 17561 20579 17595
rect 21373 17561 21407 17595
rect 21925 17561 21959 17595
rect 24409 17561 24443 17595
rect 25329 17561 25363 17595
rect 25881 17561 25915 17595
rect 26065 17561 26099 17595
rect 27638 17561 27672 17595
rect 36645 17561 36679 17595
rect 38945 17561 38979 17595
rect 39313 17561 39347 17595
rect 6193 17493 6227 17527
rect 11345 17493 11379 17527
rect 13185 17493 13219 17527
rect 15945 17493 15979 17527
rect 18705 17493 18739 17527
rect 20177 17493 20211 17527
rect 23213 17493 23247 17527
rect 26525 17493 26559 17527
rect 28825 17493 28859 17527
rect 34805 17493 34839 17527
rect 36461 17493 36495 17527
rect 4629 17289 4663 17323
rect 5825 17289 5859 17323
rect 15669 17289 15703 17323
rect 17049 17289 17083 17323
rect 27353 17289 27387 17323
rect 31493 17289 31527 17323
rect 33057 17289 33091 17323
rect 6561 17221 6595 17255
rect 16865 17221 16899 17255
rect 20729 17221 20763 17255
rect 28457 17221 28491 17255
rect 28641 17221 28675 17255
rect 29653 17221 29687 17255
rect 32137 17221 32171 17255
rect 32321 17221 32355 17255
rect 38485 17221 38519 17255
rect 39466 17221 39500 17255
rect 1869 17153 1903 17187
rect 2053 17153 2087 17187
rect 5181 17153 5215 17187
rect 5344 17153 5378 17187
rect 5457 17153 5491 17187
rect 5549 17153 5583 17187
rect 6745 17153 6779 17187
rect 7205 17153 7239 17187
rect 7389 17153 7423 17187
rect 7481 17153 7515 17187
rect 7573 17153 7607 17187
rect 8316 17153 8350 17187
rect 8565 17153 8599 17187
rect 10517 17153 10551 17187
rect 10701 17153 10735 17187
rect 11529 17153 11563 17187
rect 11785 17153 11819 17187
rect 13369 17153 13403 17187
rect 13553 17153 13587 17187
rect 13645 17153 13679 17187
rect 13737 17153 13771 17187
rect 14473 17153 14507 17187
rect 15117 17153 15151 17187
rect 15853 17153 15887 17187
rect 16681 17153 16715 17187
rect 18889 17153 18923 17187
rect 19073 17153 19107 17187
rect 19165 17153 19199 17187
rect 19257 17153 19291 17187
rect 20591 17153 20625 17187
rect 20821 17153 20855 17187
rect 20949 17153 20983 17187
rect 21097 17153 21131 17187
rect 23314 17153 23348 17187
rect 24501 17153 24535 17187
rect 25145 17153 25179 17187
rect 25329 17153 25363 17187
rect 26433 17153 26467 17187
rect 27629 17153 27663 17187
rect 27718 17156 27752 17190
rect 27813 17153 27847 17187
rect 27997 17153 28031 17187
rect 28825 17153 28859 17187
rect 29561 17153 29595 17187
rect 29745 17153 29779 17187
rect 29929 17153 29963 17187
rect 30849 17153 30883 17187
rect 31033 17153 31067 17187
rect 31125 17153 31159 17187
rect 31263 17153 31297 17187
rect 34170 17153 34204 17187
rect 34437 17153 34471 17187
rect 35541 17153 35575 17187
rect 37841 17153 37875 17187
rect 38025 17153 38059 17187
rect 38120 17156 38154 17190
rect 38229 17153 38263 17187
rect 39221 17153 39255 17187
rect 7849 17085 7883 17119
rect 17509 17085 17543 17119
rect 23581 17085 23615 17119
rect 35265 17085 35299 17119
rect 6377 17017 6411 17051
rect 12909 17017 12943 17051
rect 19441 17017 19475 17051
rect 22201 17017 22235 17051
rect 24685 17017 24719 17051
rect 67649 17017 67683 17051
rect 2237 16949 2271 16983
rect 9689 16949 9723 16983
rect 10885 16949 10919 16983
rect 14013 16949 14047 16983
rect 20453 16949 20487 16983
rect 25513 16949 25547 16983
rect 29377 16949 29411 16983
rect 32505 16949 32539 16983
rect 37289 16949 37323 16983
rect 40601 16949 40635 16983
rect 3249 16745 3283 16779
rect 5181 16745 5215 16779
rect 7849 16745 7883 16779
rect 11345 16745 11379 16779
rect 15485 16745 15519 16779
rect 22109 16745 22143 16779
rect 34805 16745 34839 16779
rect 38117 16745 38151 16779
rect 5917 16677 5951 16711
rect 8309 16677 8343 16711
rect 20545 16677 20579 16711
rect 23765 16677 23799 16711
rect 35265 16677 35299 16711
rect 14105 16609 14139 16643
rect 16037 16609 16071 16643
rect 25789 16609 25823 16643
rect 28549 16609 28583 16643
rect 29837 16609 29871 16643
rect 33057 16609 33091 16643
rect 36645 16609 36679 16643
rect 2053 16541 2087 16575
rect 2232 16541 2266 16575
rect 2332 16535 2366 16569
rect 2467 16541 2501 16575
rect 3801 16541 3835 16575
rect 5733 16541 5767 16575
rect 6469 16541 6503 16575
rect 6837 16541 6871 16575
rect 10241 16541 10275 16575
rect 10425 16541 10459 16575
rect 10517 16541 10551 16575
rect 10655 16541 10689 16575
rect 12403 16541 12437 16575
rect 12633 16541 12667 16575
rect 14361 16541 14395 16575
rect 16773 16541 16807 16575
rect 16865 16541 16899 16575
rect 16957 16541 16991 16575
rect 17141 16541 17175 16575
rect 18337 16541 18371 16575
rect 18429 16541 18463 16575
rect 18521 16541 18555 16575
rect 18705 16541 18739 16575
rect 19625 16541 19659 16575
rect 21465 16541 21499 16575
rect 21628 16541 21662 16575
rect 21741 16541 21775 16575
rect 21833 16541 21867 16575
rect 29561 16541 29595 16575
rect 31033 16541 31067 16575
rect 31401 16541 31435 16575
rect 32781 16541 32815 16575
rect 33701 16541 33735 16575
rect 2697 16473 2731 16507
rect 4046 16473 4080 16507
rect 6653 16473 6687 16507
rect 6745 16473 6779 16507
rect 7481 16473 7515 16507
rect 7665 16473 7699 16507
rect 10885 16473 10919 16507
rect 19257 16473 19291 16507
rect 19441 16473 19475 16507
rect 25544 16473 25578 16507
rect 26801 16473 26835 16507
rect 31125 16473 31159 16507
rect 31217 16473 31251 16507
rect 33517 16473 33551 16507
rect 36378 16473 36412 16507
rect 37749 16473 37783 16507
rect 37933 16473 37967 16507
rect 7021 16405 7055 16439
rect 16497 16405 16531 16439
rect 18061 16405 18095 16439
rect 24409 16405 24443 16439
rect 26341 16405 26375 16439
rect 30849 16405 30883 16439
rect 33885 16405 33919 16439
rect 8677 16201 8711 16235
rect 14381 16201 14415 16235
rect 17049 16201 17083 16235
rect 17969 16201 18003 16235
rect 21833 16201 21867 16235
rect 23213 16201 23247 16235
rect 25789 16201 25823 16235
rect 29929 16201 29963 16235
rect 32965 16201 32999 16235
rect 34529 16201 34563 16235
rect 35909 16201 35943 16235
rect 5181 16133 5215 16167
rect 7389 16133 7423 16167
rect 12817 16133 12851 16167
rect 15301 16133 15335 16167
rect 16681 16133 16715 16167
rect 19901 16133 19935 16167
rect 19993 16133 20027 16167
rect 23857 16133 23891 16167
rect 24041 16133 24075 16167
rect 24869 16133 24903 16167
rect 28641 16133 28675 16167
rect 31125 16133 31159 16167
rect 38393 16133 38427 16167
rect 40334 16133 40368 16167
rect 2053 16065 2087 16099
rect 2237 16065 2271 16099
rect 2329 16065 2363 16099
rect 2467 16065 2501 16099
rect 3157 16065 3191 16099
rect 4905 16065 4939 16099
rect 5089 16065 5123 16099
rect 5273 16065 5307 16099
rect 6377 16065 6411 16099
rect 6561 16065 6595 16099
rect 7573 16065 7607 16099
rect 12633 16065 12667 16099
rect 15025 16065 15059 16099
rect 15209 16065 15243 16099
rect 15393 16065 15427 16099
rect 16865 16065 16899 16099
rect 19625 16065 19659 16099
rect 19718 16065 19752 16099
rect 20090 16065 20124 16099
rect 21281 16065 21315 16099
rect 24685 16065 24719 16099
rect 26065 16065 26099 16099
rect 26157 16065 26191 16099
rect 26249 16065 26283 16099
rect 26433 16065 26467 16099
rect 27905 16065 27939 16099
rect 31033 16065 31067 16099
rect 31217 16065 31251 16099
rect 31401 16065 31435 16099
rect 32321 16065 32355 16099
rect 32505 16065 32539 16099
rect 32597 16065 32631 16099
rect 32689 16065 32723 16099
rect 33885 16065 33919 16099
rect 34069 16065 34103 16099
rect 34161 16065 34195 16099
rect 34253 16065 34287 16099
rect 35725 16065 35759 16099
rect 37749 16065 37783 16099
rect 37912 16065 37946 16099
rect 38012 16065 38046 16099
rect 38117 16065 38151 16099
rect 21189 15997 21223 16031
rect 28181 15997 28215 16031
rect 40601 15997 40635 16031
rect 5457 15929 5491 15963
rect 8033 15929 8067 15963
rect 15577 15929 15611 15963
rect 2697 15861 2731 15895
rect 6469 15861 6503 15895
rect 7205 15861 7239 15895
rect 12173 15861 12207 15895
rect 13001 15861 13035 15895
rect 13553 15861 13587 15895
rect 20269 15861 20303 15895
rect 20913 15861 20947 15895
rect 21097 15861 21131 15895
rect 24501 15861 24535 15895
rect 30849 15861 30883 15895
rect 36645 15861 36679 15895
rect 39221 15861 39255 15895
rect 67649 15861 67683 15895
rect 2237 15657 2271 15691
rect 7113 15657 7147 15691
rect 10885 15657 10919 15691
rect 15761 15657 15795 15691
rect 18705 15657 18739 15691
rect 20775 15657 20809 15691
rect 21833 15657 21867 15691
rect 22293 15657 22327 15691
rect 25881 15657 25915 15691
rect 27353 15657 27387 15691
rect 29561 15657 29595 15691
rect 35449 15657 35483 15691
rect 38853 15657 38887 15691
rect 25697 15589 25731 15623
rect 26893 15589 26927 15623
rect 33701 15589 33735 15623
rect 6193 15521 6227 15555
rect 6469 15521 6503 15555
rect 7573 15521 7607 15555
rect 9045 15521 9079 15555
rect 25973 15521 26007 15555
rect 36921 15521 36955 15555
rect 41245 15521 41279 15555
rect 1869 15453 1903 15487
rect 3801 15453 3835 15487
rect 4057 15453 4091 15487
rect 6929 15453 6963 15487
rect 7849 15453 7883 15487
rect 8953 15453 8987 15487
rect 9137 15453 9171 15487
rect 12173 15453 12207 15487
rect 12909 15453 12943 15487
rect 13001 15453 13035 15487
rect 13093 15453 13127 15487
rect 13277 15453 13311 15487
rect 14565 15453 14599 15487
rect 15945 15453 15979 15487
rect 16405 15453 16439 15487
rect 17325 15453 17359 15487
rect 17592 15453 17626 15487
rect 19441 15453 19475 15487
rect 19534 15453 19568 15487
rect 19717 15453 19751 15487
rect 19947 15453 19981 15487
rect 20545 15453 20579 15487
rect 22017 15453 22051 15487
rect 22109 15453 22143 15487
rect 22293 15453 22327 15487
rect 25053 15453 25087 15487
rect 26065 15453 26099 15487
rect 27077 15453 27111 15487
rect 27169 15453 27203 15487
rect 28273 15453 28307 15487
rect 28365 15453 28399 15487
rect 28641 15453 28675 15487
rect 30205 15453 30239 15487
rect 32597 15453 32631 15487
rect 32760 15453 32794 15487
rect 32876 15453 32910 15487
rect 32965 15453 32999 15487
rect 35633 15453 35667 15487
rect 35725 15453 35759 15487
rect 36001 15453 36035 15487
rect 36553 15453 36587 15487
rect 37381 15453 37415 15487
rect 37560 15453 37594 15487
rect 37660 15453 37694 15487
rect 37749 15453 37783 15487
rect 40978 15453 41012 15487
rect 2053 15385 2087 15419
rect 14749 15385 14783 15419
rect 19809 15385 19843 15419
rect 24869 15385 24903 15419
rect 27353 15385 27387 15419
rect 28457 15385 28491 15419
rect 30450 15385 30484 15419
rect 35817 15385 35851 15419
rect 36737 15385 36771 15419
rect 38025 15385 38059 15419
rect 38485 15385 38519 15419
rect 38669 15385 38703 15419
rect 5181 15317 5215 15351
rect 12633 15317 12667 15351
rect 20085 15317 20119 15351
rect 25237 15317 25271 15351
rect 28089 15317 28123 15351
rect 31585 15317 31619 15351
rect 32137 15317 32171 15351
rect 33241 15317 33275 15351
rect 39865 15317 39899 15351
rect 8033 15113 8067 15147
rect 10333 15113 10367 15147
rect 15669 15113 15703 15147
rect 18061 15113 18095 15147
rect 28917 15113 28951 15147
rect 29561 15113 29595 15147
rect 30849 15113 30883 15147
rect 32505 15113 32539 15147
rect 33057 15113 33091 15147
rect 35909 15113 35943 15147
rect 2145 15045 2179 15079
rect 5365 15045 5399 15079
rect 6745 15045 6779 15079
rect 11713 15045 11747 15079
rect 12786 15045 12820 15079
rect 25053 15045 25087 15079
rect 26157 15045 26191 15079
rect 28098 15045 28132 15079
rect 31309 15045 31343 15079
rect 32137 15045 32171 15079
rect 32321 15045 32355 15079
rect 34170 15045 34204 15079
rect 35173 15045 35207 15079
rect 36277 15045 36311 15079
rect 1961 14977 1995 15011
rect 5089 14977 5123 15011
rect 5273 14977 5307 15011
rect 5457 14977 5491 15011
rect 8953 14977 8987 15011
rect 9220 14977 9254 15011
rect 11897 14977 11931 15011
rect 14381 14977 14415 15011
rect 16681 14977 16715 15011
rect 16937 14977 16971 15011
rect 20453 14977 20487 15011
rect 20729 14977 20763 15011
rect 22017 14977 22051 15011
rect 22293 14977 22327 15011
rect 24061 14977 24095 15011
rect 25513 14977 25547 15011
rect 25676 14983 25710 15017
rect 25776 14983 25810 15017
rect 25881 14977 25915 15011
rect 28365 14977 28399 15011
rect 29837 14977 29871 15011
rect 29929 14977 29963 15011
rect 30021 14977 30055 15011
rect 30205 14977 30239 15011
rect 30665 14977 30699 15011
rect 31493 14977 31527 15011
rect 35081 14977 35115 15011
rect 35265 14977 35299 15011
rect 35449 14977 35483 15011
rect 36093 14977 36127 15011
rect 36185 14977 36219 15011
rect 36461 14977 36495 15011
rect 37381 14977 37415 15011
rect 12541 14909 12575 14943
rect 22201 14909 22235 14943
rect 24317 14909 24351 14943
rect 34437 14909 34471 14943
rect 5641 14841 5675 14875
rect 13921 14841 13955 14875
rect 22937 14841 22971 14875
rect 26985 14841 27019 14875
rect 37841 14841 37875 14875
rect 1777 14773 1811 14807
rect 12081 14773 12115 14807
rect 22293 14773 22327 14807
rect 22477 14773 22511 14807
rect 34897 14773 34931 14807
rect 7297 14569 7331 14603
rect 9873 14569 9907 14603
rect 11989 14569 12023 14603
rect 17233 14569 17267 14603
rect 22293 14569 22327 14603
rect 25053 14569 25087 14603
rect 2881 14501 2915 14535
rect 9321 14501 9355 14535
rect 22109 14501 22143 14535
rect 26801 14501 26835 14535
rect 29929 14501 29963 14535
rect 30481 14501 30515 14535
rect 30941 14501 30975 14535
rect 4077 14433 4111 14467
rect 10609 14433 10643 14467
rect 22385 14433 22419 14467
rect 1777 14365 1811 14399
rect 1961 14365 1995 14399
rect 2053 14365 2087 14399
rect 2145 14365 2179 14399
rect 3801 14365 3835 14399
rect 5089 14365 5123 14399
rect 5273 14365 5307 14399
rect 5365 14365 5399 14399
rect 5457 14365 5491 14399
rect 6653 14365 6687 14399
rect 6837 14365 6871 14399
rect 6929 14365 6963 14399
rect 7021 14365 7055 14399
rect 7757 14365 7791 14399
rect 7941 14365 7975 14399
rect 8033 14365 8067 14399
rect 8125 14365 8159 14399
rect 14841 14365 14875 14399
rect 15025 14365 15059 14399
rect 15117 14365 15151 14399
rect 15209 14365 15243 14399
rect 15853 14365 15887 14399
rect 15946 14365 15980 14399
rect 16318 14365 16352 14399
rect 17141 14365 17175 14399
rect 17325 14365 17359 14399
rect 20729 14365 20763 14399
rect 22477 14365 22511 14399
rect 25329 14365 25363 14399
rect 25421 14365 25455 14399
rect 25513 14365 25547 14399
rect 25697 14365 25731 14399
rect 28089 14365 28123 14399
rect 28181 14365 28215 14399
rect 28457 14365 28491 14399
rect 31677 14365 31711 14399
rect 31953 14365 31987 14399
rect 37657 14365 37691 14399
rect 37836 14359 37870 14393
rect 37936 14365 37970 14399
rect 38045 14365 38079 14399
rect 38945 14365 38979 14399
rect 68109 14365 68143 14399
rect 8953 14297 8987 14331
rect 9137 14297 9171 14331
rect 10876 14297 10910 14331
rect 14197 14297 14231 14331
rect 16129 14297 16163 14331
rect 16221 14297 16255 14331
rect 26249 14297 26283 14331
rect 28273 14297 28307 14331
rect 29561 14297 29595 14331
rect 29745 14297 29779 14331
rect 31125 14297 31159 14331
rect 34161 14297 34195 14331
rect 36829 14297 36863 14331
rect 38761 14297 38795 14331
rect 2421 14229 2455 14263
rect 5733 14229 5767 14263
rect 8401 14229 8435 14263
rect 12817 14229 12851 14263
rect 13369 14229 13403 14263
rect 15393 14229 15427 14263
rect 16497 14229 16531 14263
rect 17509 14229 17543 14263
rect 20269 14229 20303 14263
rect 20913 14229 20947 14263
rect 24593 14229 24627 14263
rect 27905 14229 27939 14263
rect 29009 14229 29043 14263
rect 32965 14229 32999 14263
rect 35541 14229 35575 14263
rect 38301 14229 38335 14263
rect 39129 14229 39163 14263
rect 4077 14025 4111 14059
rect 6745 14025 6779 14059
rect 10793 14025 10827 14059
rect 11529 14025 11563 14059
rect 13921 14025 13955 14059
rect 24041 14025 24075 14059
rect 33701 14025 33735 14059
rect 35265 14025 35299 14059
rect 37749 14025 37783 14059
rect 38945 14025 38979 14059
rect 7205 13957 7239 13991
rect 9658 13957 9692 13991
rect 14841 13957 14875 13991
rect 15945 13957 15979 13991
rect 25973 13957 26007 13991
rect 28089 13957 28123 13991
rect 31217 13957 31251 13991
rect 33793 13957 33827 13991
rect 34621 13957 34655 13991
rect 37565 13957 37599 13991
rect 40058 13957 40092 13991
rect 2697 13889 2731 13923
rect 2953 13889 2987 13923
rect 4537 13889 4571 13923
rect 4813 13889 4847 13923
rect 6469 13889 6503 13923
rect 6561 13889 6595 13923
rect 7389 13889 7423 13923
rect 8677 13889 8711 13923
rect 9413 13889 9447 13923
rect 11805 13889 11839 13923
rect 11897 13889 11931 13923
rect 11989 13889 12023 13923
rect 12173 13889 12207 13923
rect 13093 13889 13127 13923
rect 14105 13889 14139 13923
rect 14657 13889 14691 13923
rect 15577 13889 15611 13923
rect 15761 13889 15795 13923
rect 16681 13889 16715 13923
rect 16865 13889 16899 13923
rect 18061 13889 18095 13923
rect 18317 13889 18351 13923
rect 19901 13889 19935 13923
rect 20168 13889 20202 13923
rect 22293 13889 22327 13923
rect 22937 13889 22971 13923
rect 23581 13889 23615 13923
rect 23857 13889 23891 13923
rect 25053 13889 25087 13923
rect 25145 13889 25179 13923
rect 25237 13889 25271 13923
rect 25421 13889 25455 13923
rect 27077 13889 27111 13923
rect 27997 13889 28031 13923
rect 28181 13889 28215 13923
rect 28365 13889 28399 13923
rect 31401 13889 31435 13923
rect 32643 13889 32677 13923
rect 32778 13889 32812 13923
rect 32894 13889 32928 13923
rect 33057 13889 33091 13923
rect 34805 13889 34839 13923
rect 36378 13889 36412 13923
rect 36645 13889 36679 13923
rect 37381 13889 37415 13923
rect 40325 13889 40359 13923
rect 1961 13821 1995 13855
rect 2237 13821 2271 13855
rect 7573 13821 7607 13855
rect 8953 13821 8987 13855
rect 22477 13821 22511 13855
rect 23673 13821 23707 13855
rect 28825 13821 28859 13855
rect 29101 13821 29135 13855
rect 30665 13821 30699 13855
rect 34437 13821 34471 13855
rect 13277 13753 13311 13787
rect 17049 13753 17083 13787
rect 27813 13753 27847 13787
rect 31585 13753 31619 13787
rect 16681 13685 16715 13719
rect 19441 13685 19475 13719
rect 21281 13685 21315 13719
rect 23857 13685 23891 13719
rect 24777 13685 24811 13719
rect 32413 13685 32447 13719
rect 2973 13481 3007 13515
rect 4629 13481 4663 13515
rect 9321 13481 9355 13515
rect 12541 13481 12575 13515
rect 13553 13481 13587 13515
rect 17325 13481 17359 13515
rect 19441 13481 19475 13515
rect 21281 13481 21315 13515
rect 36001 13481 36035 13515
rect 37381 13481 37415 13515
rect 6469 13413 6503 13447
rect 13461 13413 13495 13447
rect 14473 13413 14507 13447
rect 16589 13413 16623 13447
rect 16773 13413 16807 13447
rect 30573 13413 30607 13447
rect 34805 13413 34839 13447
rect 5089 13345 5123 13379
rect 7113 13345 7147 13379
rect 10241 13345 10275 13379
rect 15301 13345 15335 13379
rect 18613 13345 18647 13379
rect 23489 13345 23523 13379
rect 25605 13345 25639 13379
rect 34161 13345 34195 13379
rect 4261 13277 4295 13311
rect 5356 13277 5390 13311
rect 7941 13277 7975 13311
rect 9965 13277 9999 13311
rect 11529 13277 11563 13311
rect 11805 13277 11839 13311
rect 11897 13277 11931 13311
rect 15393 13277 15427 13311
rect 15577 13277 15611 13311
rect 18337 13277 18371 13311
rect 19533 13277 19567 13311
rect 19625 13277 19659 13311
rect 21097 13277 21131 13311
rect 23233 13277 23267 13311
rect 25329 13277 25363 13311
rect 26249 13277 26283 13311
rect 28641 13277 28675 13311
rect 28733 13277 28767 13311
rect 29009 13277 29043 13311
rect 29745 13277 29779 13311
rect 29837 13277 29871 13311
rect 30113 13277 30147 13311
rect 31953 13277 31987 13311
rect 35357 13277 35391 13311
rect 35541 13277 35575 13311
rect 35633 13277 35667 13311
rect 35725 13277 35759 13311
rect 37841 13277 37875 13311
rect 38025 13277 38059 13311
rect 38117 13277 38151 13311
rect 38209 13277 38243 13311
rect 39313 13277 39347 13311
rect 40233 13277 40267 13311
rect 68109 13277 68143 13311
rect 2237 13209 2271 13243
rect 2421 13209 2455 13243
rect 4445 13209 4479 13243
rect 7297 13209 7331 13243
rect 8125 13209 8159 13243
rect 9413 13209 9447 13243
rect 11713 13209 11747 13243
rect 13093 13209 13127 13243
rect 14105 13209 14139 13243
rect 16313 13209 16347 13243
rect 26494 13209 26528 13243
rect 28825 13209 28859 13243
rect 29929 13209 29963 13243
rect 31708 13209 31742 13243
rect 33894 13209 33928 13243
rect 2053 13141 2087 13175
rect 8309 13141 8343 13175
rect 12081 13141 12115 13175
rect 14565 13141 14599 13175
rect 19257 13141 19291 13175
rect 20637 13141 20671 13175
rect 22109 13141 22143 13175
rect 27629 13141 27663 13175
rect 28457 13141 28491 13175
rect 29561 13141 29595 13175
rect 32781 13141 32815 13175
rect 38485 13141 38519 13175
rect 41521 13141 41555 13175
rect 4537 12937 4571 12971
rect 5273 12937 5307 12971
rect 6469 12937 6503 12971
rect 18061 12937 18095 12971
rect 20085 12937 20119 12971
rect 22385 12937 22419 12971
rect 24133 12937 24167 12971
rect 24961 12937 24995 12971
rect 26065 12937 26099 12971
rect 26985 12937 27019 12971
rect 28089 12937 28123 12971
rect 39865 12937 39899 12971
rect 10517 12869 10551 12903
rect 11713 12869 11747 12903
rect 22017 12869 22051 12903
rect 24777 12869 24811 12903
rect 27261 12869 27295 12903
rect 27353 12869 27387 12903
rect 32413 12869 32447 12903
rect 35725 12869 35759 12903
rect 40978 12869 41012 12903
rect 2697 12801 2731 12835
rect 3157 12801 3191 12835
rect 3413 12801 3447 12835
rect 6653 12801 6687 12835
rect 7941 12801 7975 12835
rect 8657 12801 8691 12835
rect 10241 12801 10275 12835
rect 10425 12801 10459 12835
rect 10609 12801 10643 12835
rect 11529 12801 11563 12835
rect 11805 12801 11839 12835
rect 11897 12801 11931 12835
rect 12725 12801 12759 12835
rect 12909 12801 12943 12835
rect 13737 12801 13771 12835
rect 15301 12801 15335 12835
rect 17601 12801 17635 12835
rect 18337 12801 18371 12835
rect 18429 12801 18463 12835
rect 18521 12801 18555 12835
rect 18705 12801 18739 12835
rect 19441 12801 19475 12835
rect 19625 12801 19659 12835
rect 19717 12801 19751 12835
rect 19809 12801 19843 12835
rect 20545 12801 20579 12835
rect 20729 12801 20763 12835
rect 21833 12801 21867 12835
rect 22109 12801 22143 12835
rect 22247 12801 22281 12835
rect 23673 12801 23707 12835
rect 23949 12801 23983 12835
rect 24593 12801 24627 12835
rect 25421 12801 25455 12835
rect 25605 12801 25639 12835
rect 25697 12801 25731 12835
rect 25789 12801 25823 12835
rect 27169 12801 27203 12835
rect 27537 12801 27571 12835
rect 28825 12801 28859 12835
rect 29101 12801 29135 12835
rect 32229 12801 32263 12835
rect 35909 12801 35943 12835
rect 37565 12801 37599 12835
rect 38761 12801 38795 12835
rect 38945 12801 38979 12835
rect 41245 12801 41279 12835
rect 2421 12733 2455 12767
rect 5825 12733 5859 12767
rect 7665 12733 7699 12767
rect 8401 12733 8435 12767
rect 17509 12733 17543 12767
rect 20913 12733 20947 12767
rect 23765 12733 23799 12767
rect 37289 12733 37323 12767
rect 9781 12665 9815 12699
rect 12081 12665 12115 12699
rect 12909 12665 12943 12699
rect 13553 12665 13587 12699
rect 15577 12665 15611 12699
rect 15761 12665 15795 12699
rect 10793 12597 10827 12631
rect 14197 12597 14231 12631
rect 17233 12597 17267 12631
rect 17601 12597 17635 12631
rect 23949 12597 23983 12631
rect 32597 12597 32631 12631
rect 34897 12597 34931 12631
rect 35541 12597 35575 12631
rect 38577 12597 38611 12631
rect 2605 12393 2639 12427
rect 5733 12393 5767 12427
rect 8217 12393 8251 12427
rect 13093 12393 13127 12427
rect 17785 12393 17819 12427
rect 22293 12393 22327 12427
rect 24409 12393 24443 12427
rect 25329 12393 25363 12427
rect 28273 12393 28307 12427
rect 33149 12393 33183 12427
rect 3801 12325 3835 12359
rect 14381 12325 14415 12359
rect 15209 12325 15243 12359
rect 10517 12257 10551 12291
rect 16313 12257 16347 12291
rect 28089 12257 28123 12291
rect 31953 12257 31987 12291
rect 37105 12257 37139 12291
rect 1961 12189 1995 12223
rect 2145 12189 2179 12223
rect 2237 12189 2271 12223
rect 2375 12189 2409 12223
rect 3065 12189 3099 12223
rect 3985 12189 4019 12223
rect 6469 12189 6503 12223
rect 6561 12189 6595 12223
rect 6653 12189 6687 12223
rect 6837 12189 6871 12223
rect 7573 12189 7607 12223
rect 7736 12189 7770 12223
rect 7852 12186 7886 12220
rect 7941 12189 7975 12223
rect 9505 12189 9539 12223
rect 9781 12189 9815 12223
rect 9873 12189 9907 12223
rect 10793 12189 10827 12223
rect 11897 12189 11931 12223
rect 12626 12189 12660 12223
rect 13093 12189 13127 12223
rect 13277 12189 13311 12223
rect 14105 12189 14139 12223
rect 14381 12189 14415 12223
rect 15209 12189 15243 12223
rect 15485 12189 15519 12223
rect 15945 12189 15979 12223
rect 16221 12189 16255 12223
rect 17969 12189 18003 12223
rect 19717 12189 19751 12223
rect 21741 12189 21775 12223
rect 22109 12189 22143 12223
rect 25145 12189 25179 12223
rect 27997 12189 28031 12223
rect 28273 12189 28307 12223
rect 29745 12189 29779 12223
rect 29929 12189 29963 12223
rect 30113 12189 30147 12223
rect 32505 12189 32539 12223
rect 32668 12189 32702 12223
rect 32781 12189 32815 12223
rect 32873 12189 32907 12223
rect 35357 12189 35391 12223
rect 35449 12189 35483 12223
rect 35541 12189 35575 12223
rect 35725 12189 35759 12223
rect 36829 12189 36863 12223
rect 37657 12189 37691 12223
rect 37841 12189 37875 12223
rect 37933 12189 37967 12223
rect 38025 12189 38059 12223
rect 38761 12189 38795 12223
rect 41245 12189 41279 12223
rect 5181 12121 5215 12155
rect 9689 12121 9723 12155
rect 18153 12121 18187 12155
rect 19901 12121 19935 12155
rect 21925 12121 21959 12155
rect 22017 12121 22051 12155
rect 24961 12121 24995 12155
rect 25789 12121 25823 12155
rect 29837 12121 29871 12155
rect 38301 12121 38335 12155
rect 40978 12121 41012 12155
rect 4629 12053 4663 12087
rect 6193 12053 6227 12087
rect 9045 12053 9079 12087
rect 10057 12053 10091 12087
rect 12449 12053 12483 12087
rect 18705 12053 18739 12087
rect 20085 12053 20119 12087
rect 27077 12053 27111 12087
rect 28457 12053 28491 12087
rect 29561 12053 29595 12087
rect 35081 12053 35115 12087
rect 39865 12053 39899 12087
rect 5457 11849 5491 11883
rect 13461 11849 13495 11883
rect 14197 11849 14231 11883
rect 14933 11849 14967 11883
rect 21281 11849 21315 11883
rect 22477 11849 22511 11883
rect 27445 11849 27479 11883
rect 34069 11849 34103 11883
rect 2605 11781 2639 11815
rect 3402 11781 3436 11815
rect 5641 11781 5675 11815
rect 12633 11781 12667 11815
rect 15853 11781 15887 11815
rect 18337 11781 18371 11815
rect 20146 11781 20180 11815
rect 24501 11781 24535 11815
rect 29469 11781 29503 11815
rect 29561 11781 29595 11815
rect 31340 11781 31374 11815
rect 32229 11781 32263 11815
rect 35182 11781 35216 11815
rect 1961 11713 1995 11747
rect 2145 11713 2179 11747
rect 2237 11713 2271 11747
rect 2375 11713 2409 11747
rect 5825 11713 5859 11747
rect 6745 11713 6779 11747
rect 8953 11713 8987 11747
rect 10425 11713 10459 11747
rect 11529 11713 11563 11747
rect 11713 11713 11747 11747
rect 11805 11713 11839 11747
rect 11897 11713 11931 11747
rect 12541 11713 12575 11747
rect 12725 11713 12759 11747
rect 13645 11713 13679 11747
rect 14381 11713 14415 11747
rect 16037 11713 16071 11747
rect 18153 11713 18187 11747
rect 19901 11713 19935 11747
rect 23601 11713 23635 11747
rect 24317 11713 24351 11747
rect 25329 11713 25363 11747
rect 25513 11713 25547 11747
rect 25605 11713 25639 11747
rect 25697 11713 25731 11747
rect 26985 11713 27019 11747
rect 27261 11713 27295 11747
rect 27997 11713 28031 11747
rect 28641 11713 28675 11747
rect 29377 11713 29411 11747
rect 29745 11713 29779 11747
rect 31585 11713 31619 11747
rect 32505 11713 32539 11747
rect 32597 11713 32631 11747
rect 32689 11713 32723 11747
rect 32873 11713 32907 11747
rect 35449 11713 35483 11747
rect 36369 11713 36403 11747
rect 36553 11713 36587 11747
rect 37473 11713 37507 11747
rect 37657 11713 37691 11747
rect 37749 11713 37783 11747
rect 37841 11713 37875 11747
rect 40242 11713 40276 11747
rect 40509 11713 40543 11747
rect 3157 11645 3191 11679
rect 9505 11645 9539 11679
rect 10149 11645 10183 11679
rect 23857 11645 23891 11679
rect 27077 11645 27111 11679
rect 36737 11645 36771 11679
rect 38117 11645 38151 11679
rect 4537 11577 4571 11611
rect 12081 11577 12115 11611
rect 28181 11577 28215 11611
rect 67649 11577 67683 11611
rect 8033 11509 8067 11543
rect 16681 11509 16715 11543
rect 17601 11509 17635 11543
rect 18521 11509 18555 11543
rect 19349 11509 19383 11543
rect 24685 11509 24719 11543
rect 25973 11509 26007 11543
rect 27261 11509 27295 11543
rect 29193 11509 29227 11543
rect 30205 11509 30239 11543
rect 39129 11509 39163 11543
rect 1961 11305 1995 11339
rect 2789 11305 2823 11339
rect 5181 11305 5215 11339
rect 7205 11305 7239 11339
rect 13369 11305 13403 11339
rect 17785 11305 17819 11339
rect 18429 11305 18463 11339
rect 20361 11305 20395 11339
rect 22017 11305 22051 11339
rect 23857 11305 23891 11339
rect 24685 11305 24719 11339
rect 25789 11305 25823 11339
rect 27905 11305 27939 11339
rect 29561 11305 29595 11339
rect 32229 11305 32263 11339
rect 34069 11305 34103 11339
rect 38025 11305 38059 11339
rect 12541 11237 12575 11271
rect 28917 11237 28951 11271
rect 37013 11237 37047 11271
rect 8953 11169 8987 11203
rect 11989 11169 12023 11203
rect 22477 11169 22511 11203
rect 32689 11169 32723 11203
rect 35081 11169 35115 11203
rect 2145 11101 2179 11135
rect 6561 11101 6595 11135
rect 7665 11101 7699 11135
rect 7849 11101 7883 11135
rect 7941 11101 7975 11135
rect 8079 11101 8113 11135
rect 12725 11101 12759 11135
rect 13185 11101 13219 11135
rect 15761 11101 15795 11135
rect 16405 11101 16439 11135
rect 18521 11101 18555 11135
rect 18613 11101 18647 11135
rect 19717 11101 19751 11135
rect 19896 11098 19930 11132
rect 19996 11101 20030 11135
rect 20131 11101 20165 11135
rect 21373 11101 21407 11135
rect 23121 11101 23155 11135
rect 23305 11101 23339 11135
rect 24915 11101 24949 11135
rect 25053 11101 25087 11135
rect 25145 11101 25179 11135
rect 25329 11101 25363 11135
rect 26525 11101 26559 11135
rect 26781 11101 26815 11135
rect 28365 11101 28399 11135
rect 28549 11101 28583 11135
rect 28641 11101 28675 11135
rect 28733 11101 28767 11135
rect 29745 11101 29779 11135
rect 29837 11101 29871 11135
rect 29929 11101 29963 11135
rect 30113 11101 30147 11135
rect 31861 11101 31895 11135
rect 32045 11101 32079 11135
rect 34897 11101 34931 11135
rect 35541 11101 35575 11135
rect 35725 11101 35759 11135
rect 37197 11101 37231 11135
rect 37289 11101 37323 11135
rect 37565 11101 37599 11135
rect 2329 11033 2363 11067
rect 6294 11033 6328 11067
rect 8309 11033 8343 11067
rect 9198 11033 9232 11067
rect 15494 11033 15528 11067
rect 16672 11033 16706 11067
rect 33425 11033 33459 11067
rect 33609 11033 33643 11067
rect 34713 11033 34747 11067
rect 36185 11033 36219 11067
rect 37381 11033 37415 11067
rect 10333 10965 10367 10999
rect 14381 10965 14415 10999
rect 18245 10965 18279 10999
rect 20821 10965 20855 10999
rect 33241 10965 33275 10999
rect 35541 10965 35575 10999
rect 38577 10965 38611 10999
rect 4537 10761 4571 10795
rect 7757 10761 7791 10795
rect 14473 10761 14507 10795
rect 18061 10761 18095 10795
rect 22293 10761 22327 10795
rect 24777 10761 24811 10795
rect 25697 10761 25731 10795
rect 26249 10761 26283 10795
rect 29837 10761 29871 10795
rect 32689 10761 32723 10795
rect 34529 10761 34563 10795
rect 2421 10693 2455 10727
rect 3402 10693 3436 10727
rect 7941 10693 7975 10727
rect 10333 10693 10367 10727
rect 18521 10693 18555 10727
rect 35449 10693 35483 10727
rect 38669 10693 38703 10727
rect 40242 10693 40276 10727
rect 1777 10625 1811 10659
rect 1961 10625 1995 10659
rect 2053 10625 2087 10659
rect 2145 10625 2179 10659
rect 3157 10625 3191 10659
rect 6653 10625 6687 10659
rect 6745 10625 6779 10659
rect 6837 10625 6871 10659
rect 7021 10625 7055 10659
rect 8125 10625 8159 10659
rect 8585 10625 8619 10659
rect 10149 10625 10183 10659
rect 10425 10625 10459 10659
rect 10517 10625 10551 10659
rect 12642 10625 12676 10659
rect 12909 10625 12943 10659
rect 13737 10625 13771 10659
rect 13921 10625 13955 10659
rect 14289 10625 14323 10659
rect 15945 10625 15979 10659
rect 17049 10625 17083 10659
rect 20085 10625 20119 10659
rect 20913 10625 20947 10659
rect 22201 10625 22235 10659
rect 23029 10625 23063 10659
rect 24041 10625 24075 10659
rect 24225 10625 24259 10659
rect 25329 10625 25363 10659
rect 25513 10625 25547 10659
rect 28825 10625 28859 10659
rect 29377 10625 29411 10659
rect 29653 10625 29687 10659
rect 33517 10625 33551 10659
rect 33609 10625 33643 10659
rect 33701 10625 33735 10659
rect 33885 10625 33919 10659
rect 35081 10625 35115 10659
rect 35265 10625 35299 10659
rect 37289 10625 37323 10659
rect 38025 10625 38059 10659
rect 38209 10625 38243 10659
rect 38301 10625 38335 10659
rect 38393 10625 38427 10659
rect 40509 10625 40543 10659
rect 5825 10557 5859 10591
rect 14013 10557 14047 10591
rect 14105 10557 14139 10591
rect 16129 10557 16163 10591
rect 21097 10557 21131 10591
rect 22845 10557 22879 10591
rect 29469 10557 29503 10591
rect 35909 10557 35943 10591
rect 36185 10557 36219 10591
rect 10701 10489 10735 10523
rect 17233 10489 17267 10523
rect 24133 10489 24167 10523
rect 6377 10421 6411 10455
rect 11529 10421 11563 10455
rect 20729 10421 20763 10455
rect 23213 10421 23247 10455
rect 29561 10421 29595 10455
rect 33241 10421 33275 10455
rect 37473 10421 37507 10455
rect 39129 10421 39163 10455
rect 67649 10421 67683 10455
rect 1869 10217 1903 10251
rect 6561 10217 6595 10251
rect 9045 10217 9079 10251
rect 11437 10217 11471 10251
rect 17509 10217 17543 10251
rect 18061 10217 18095 10251
rect 19349 10217 19383 10251
rect 22845 10217 22879 10251
rect 23857 10217 23891 10251
rect 27813 10217 27847 10251
rect 28917 10217 28951 10251
rect 34805 10217 34839 10251
rect 36921 10217 36955 10251
rect 38301 10217 38335 10251
rect 2789 10149 2823 10183
rect 17233 10149 17267 10183
rect 22385 10149 22419 10183
rect 28549 10149 28583 10183
rect 11897 10081 11931 10115
rect 17509 10081 17543 10115
rect 21005 10081 21039 10115
rect 24869 10081 24903 10115
rect 25145 10081 25179 10115
rect 32965 10081 32999 10115
rect 2053 10013 2087 10047
rect 2237 10013 2271 10047
rect 3801 10013 3835 10047
rect 6193 10013 6227 10047
rect 7481 10013 7515 10047
rect 7665 10013 7699 10047
rect 7757 10013 7791 10047
rect 7849 10013 7883 10047
rect 9689 10013 9723 10047
rect 9873 10013 9907 10047
rect 10057 10013 10091 10047
rect 11621 10013 11655 10047
rect 11805 10013 11839 10047
rect 11989 10013 12023 10047
rect 12173 10013 12207 10047
rect 14197 10013 14231 10047
rect 16313 10013 16347 10047
rect 17601 10013 17635 10047
rect 18337 10013 18371 10047
rect 18429 10013 18463 10047
rect 18521 10013 18555 10047
rect 18705 10013 18739 10047
rect 19809 10013 19843 10047
rect 19993 10013 20027 10047
rect 20088 10007 20122 10041
rect 20197 10013 20231 10047
rect 23673 10013 23707 10047
rect 26157 10013 26191 10047
rect 26341 10013 26375 10047
rect 26433 10013 26467 10047
rect 26525 10013 26559 10047
rect 27261 10013 27295 10047
rect 27537 10013 27571 10047
rect 27629 10013 27663 10047
rect 28733 10013 28767 10047
rect 28825 10013 28859 10047
rect 29009 10013 29043 10047
rect 29561 10013 29595 10047
rect 32709 10013 32743 10047
rect 34713 10013 34747 10047
rect 34897 10013 34931 10047
rect 35909 10013 35943 10047
rect 36185 10013 36219 10047
rect 37105 10013 37139 10047
rect 37197 10013 37231 10047
rect 37473 10013 37507 10047
rect 38117 10013 38151 10047
rect 3985 9945 4019 9979
rect 6377 9945 6411 9979
rect 9965 9945 9999 9979
rect 20453 9945 20487 9979
rect 21250 9945 21284 9979
rect 27445 9945 27479 9979
rect 37289 9945 37323 9979
rect 37933 9945 37967 9979
rect 4169 9877 4203 9911
rect 4721 9877 4755 9911
rect 8125 9877 8159 9911
rect 10241 9877 10275 9911
rect 12725 9877 12759 9911
rect 13553 9877 13587 9911
rect 14657 9877 14691 9911
rect 15301 9877 15335 9911
rect 16221 9877 16255 9911
rect 26801 9877 26835 9911
rect 31585 9877 31619 9911
rect 34161 9877 34195 9911
rect 5181 9673 5215 9707
rect 7573 9673 7607 9707
rect 19625 9673 19659 9707
rect 20315 9673 20349 9707
rect 32689 9673 32723 9707
rect 37289 9673 37323 9707
rect 8300 9605 8334 9639
rect 10241 9605 10275 9639
rect 19441 9605 19475 9639
rect 22477 9605 22511 9639
rect 25697 9605 25731 9639
rect 26065 9605 26099 9639
rect 30104 9605 30138 9639
rect 33149 9605 33183 9639
rect 34345 9605 34379 9639
rect 38485 9605 38519 9639
rect 39282 9605 39316 9639
rect 2053 9537 2087 9571
rect 2232 9540 2266 9574
rect 2329 9537 2363 9571
rect 2467 9537 2501 9571
rect 3801 9537 3835 9571
rect 4068 9537 4102 9571
rect 7205 9537 7239 9571
rect 7389 9537 7423 9571
rect 8033 9537 8067 9571
rect 9965 9537 9999 9571
rect 10149 9537 10183 9571
rect 10333 9537 10367 9571
rect 12173 9537 12207 9571
rect 12357 9537 12391 9571
rect 12725 9537 12759 9571
rect 12909 9537 12943 9571
rect 14482 9537 14516 9571
rect 15577 9537 15611 9571
rect 15853 9537 15887 9571
rect 15945 9537 15979 9571
rect 16129 9537 16163 9571
rect 17877 9537 17911 9571
rect 17969 9537 18003 9571
rect 18429 9537 18463 9571
rect 18613 9537 18647 9571
rect 19257 9537 19291 9571
rect 21833 9537 21867 9571
rect 22017 9537 22051 9571
rect 23121 9537 23155 9571
rect 24409 9537 24443 9571
rect 24501 9537 24535 9571
rect 24593 9537 24627 9571
rect 24777 9537 24811 9571
rect 25881 9537 25915 9571
rect 27997 9537 28031 9571
rect 28273 9537 28307 9571
rect 28917 9537 28951 9571
rect 29101 9537 29135 9571
rect 29193 9537 29227 9571
rect 29837 9537 29871 9571
rect 33425 9537 33459 9571
rect 33517 9537 33551 9571
rect 33609 9537 33643 9571
rect 33793 9537 33827 9571
rect 34989 9537 35023 9571
rect 35725 9537 35759 9571
rect 37841 9537 37875 9571
rect 38025 9537 38059 9571
rect 38117 9537 38151 9571
rect 38209 9537 38243 9571
rect 39037 9537 39071 9571
rect 12449 9469 12483 9503
rect 12541 9469 12575 9503
rect 14749 9469 14783 9503
rect 15761 9469 15795 9503
rect 20085 9469 20119 9503
rect 23673 9469 23707 9503
rect 26985 9469 27019 9503
rect 28089 9469 28123 9503
rect 35449 9469 35483 9503
rect 18705 9401 18739 9435
rect 28457 9401 28491 9435
rect 1593 9333 1627 9367
rect 2697 9333 2731 9367
rect 3249 9333 3283 9367
rect 9413 9333 9447 9367
rect 10517 9333 10551 9367
rect 11529 9333 11563 9367
rect 13369 9333 13403 9367
rect 15393 9333 15427 9367
rect 17141 9333 17175 9367
rect 17601 9333 17635 9367
rect 17785 9333 17819 9367
rect 21925 9333 21959 9367
rect 24133 9333 24167 9367
rect 28273 9333 28307 9367
rect 29101 9333 29135 9367
rect 29377 9333 29411 9367
rect 31217 9333 31251 9367
rect 34805 9333 34839 9367
rect 40417 9333 40451 9367
rect 3065 9129 3099 9163
rect 7021 9129 7055 9163
rect 15577 9129 15611 9163
rect 17693 9129 17727 9163
rect 24777 9129 24811 9163
rect 25329 9129 25363 9163
rect 27445 9129 27479 9163
rect 28825 9129 28859 9163
rect 30849 9129 30883 9163
rect 33149 9129 33183 9163
rect 38025 9129 38059 9163
rect 15117 9061 15151 9095
rect 18613 9061 18647 9095
rect 19533 9061 19567 9095
rect 36645 9061 36679 9095
rect 12357 8993 12391 9027
rect 12449 8993 12483 9027
rect 13553 8993 13587 9027
rect 16957 8993 16991 9027
rect 35357 8993 35391 9027
rect 1869 8925 1903 8959
rect 2053 8925 2087 8959
rect 2145 8925 2179 8959
rect 2237 8925 2271 8959
rect 4169 8925 4203 8959
rect 5641 8925 5675 8959
rect 5908 8925 5942 8959
rect 11529 8925 11563 8959
rect 12173 8925 12207 8959
rect 12541 8925 12575 8959
rect 12725 8925 12759 8959
rect 14565 8925 14599 8959
rect 16690 8925 16724 8959
rect 17785 8925 17819 8959
rect 17877 8925 17911 8959
rect 18429 8925 18463 8959
rect 18521 8925 18555 8959
rect 19349 8925 19383 8959
rect 20177 8925 20211 8959
rect 22109 8925 22143 8959
rect 26065 8925 26099 8959
rect 26332 8925 26366 8959
rect 30389 8925 30423 8959
rect 31033 8925 31067 8959
rect 31125 8925 31159 8959
rect 31401 8925 31435 8959
rect 33517 8925 33551 8959
rect 35633 8925 35667 8959
rect 36829 8925 36863 8959
rect 37013 8925 37047 8959
rect 37197 8925 37231 8959
rect 37657 8925 37691 8959
rect 37841 8925 37875 8959
rect 68109 8925 68143 8959
rect 3801 8857 3835 8891
rect 3985 8857 4019 8891
rect 11284 8857 11318 8891
rect 11989 8857 12023 8891
rect 20361 8857 20395 8891
rect 22376 8857 22410 8891
rect 24409 8857 24443 8891
rect 24593 8857 24627 8891
rect 25421 8857 25455 8891
rect 31217 8857 31251 8891
rect 33333 8857 33367 8891
rect 36921 8857 36955 8891
rect 38485 8857 38519 8891
rect 38669 8857 38703 8891
rect 2513 8789 2547 8823
rect 4721 8789 4755 8823
rect 7481 8789 7515 8823
rect 10149 8789 10183 8823
rect 17509 8789 17543 8823
rect 19993 8789 20027 8823
rect 23489 8789 23523 8823
rect 31861 8789 31895 8823
rect 33977 8789 34011 8823
rect 34805 8789 34839 8823
rect 38853 8789 38887 8823
rect 1593 8585 1627 8619
rect 3985 8585 4019 8619
rect 6469 8585 6503 8619
rect 7481 8585 7515 8619
rect 23489 8585 23523 8619
rect 28825 8585 28859 8619
rect 32137 8585 32171 8619
rect 40049 8585 40083 8619
rect 2850 8517 2884 8551
rect 5733 8517 5767 8551
rect 7113 8517 7147 8551
rect 8401 8517 8435 8551
rect 20545 8517 20579 8551
rect 23213 8517 23247 8551
rect 28457 8517 28491 8551
rect 28549 8517 28583 8551
rect 31585 8517 31619 8551
rect 32505 8517 32539 8551
rect 34161 8517 34195 8551
rect 38761 8517 38795 8551
rect 2145 8449 2179 8483
rect 4813 8449 4847 8483
rect 7021 8449 7055 8483
rect 7297 8449 7331 8483
rect 7941 8449 7975 8483
rect 8033 8449 8067 8483
rect 8217 8449 8251 8483
rect 9689 8449 9723 8483
rect 10149 8449 10183 8483
rect 10977 8449 11011 8483
rect 12081 8449 12115 8483
rect 12265 8449 12299 8483
rect 12357 8449 12391 8483
rect 12633 8449 12667 8483
rect 13921 8449 13955 8483
rect 18622 8449 18656 8483
rect 19901 8449 19935 8483
rect 20085 8452 20119 8486
rect 20177 8449 20211 8483
rect 20269 8449 20303 8483
rect 22937 8449 22971 8483
rect 23121 8449 23155 8483
rect 23305 8449 23339 8483
rect 25145 8449 25179 8483
rect 26157 8449 26191 8483
rect 28273 8449 28307 8483
rect 28641 8449 28675 8483
rect 29285 8449 29319 8483
rect 29469 8449 29503 8483
rect 32321 8449 32355 8483
rect 32413 8449 32447 8483
rect 32689 8449 32723 8483
rect 33425 8449 33459 8483
rect 34069 8449 34103 8483
rect 34253 8449 34287 8483
rect 34437 8449 34471 8483
rect 34897 8449 34931 8483
rect 35725 8449 35759 8483
rect 37565 8449 37599 8483
rect 2605 8381 2639 8415
rect 8861 8381 8895 8415
rect 12449 8381 12483 8415
rect 13645 8381 13679 8415
rect 15393 8381 15427 8415
rect 16037 8381 16071 8415
rect 18889 8381 18923 8415
rect 24869 8381 24903 8415
rect 26433 8381 26467 8415
rect 26985 8381 27019 8415
rect 27261 8381 27295 8415
rect 36001 8381 36035 8415
rect 37289 8381 37323 8415
rect 10333 8313 10367 8347
rect 10793 8313 10827 8347
rect 11529 8313 11563 8347
rect 16865 8313 16899 8347
rect 30481 8313 30515 8347
rect 33885 8313 33919 8347
rect 35081 8313 35115 8347
rect 4997 8245 5031 8279
rect 12817 8245 12851 8279
rect 17509 8245 17543 8279
rect 19349 8245 19383 8279
rect 29653 8245 29687 8279
rect 7757 8041 7791 8075
rect 8401 8041 8435 8075
rect 9781 8041 9815 8075
rect 17601 8041 17635 8075
rect 21925 8041 21959 8075
rect 23765 8041 23799 8075
rect 26893 8041 26927 8075
rect 29009 8041 29043 8075
rect 35265 8041 35299 8075
rect 37197 8041 37231 8075
rect 41245 8041 41279 8075
rect 6193 7973 6227 8007
rect 11713 7973 11747 8007
rect 2329 7905 2363 7939
rect 17135 7905 17169 7939
rect 25881 7905 25915 7939
rect 27353 7905 27387 7939
rect 27629 7905 27663 7939
rect 35817 7905 35851 7939
rect 36093 7905 36127 7939
rect 39865 7905 39899 7939
rect 2053 7837 2087 7871
rect 4813 7837 4847 7871
rect 5080 7837 5114 7871
rect 7297 7837 7331 7871
rect 7573 7837 7607 7871
rect 9321 7837 9355 7871
rect 9413 7837 9447 7871
rect 9597 7837 9631 7871
rect 10333 7837 10367 7871
rect 11529 7837 11563 7871
rect 13286 7837 13320 7871
rect 13553 7837 13587 7871
rect 15945 7837 15979 7871
rect 16865 7837 16899 7871
rect 17049 7837 17083 7871
rect 17233 7837 17267 7871
rect 17417 7837 17451 7871
rect 18245 7837 18279 7871
rect 20545 7837 20579 7871
rect 20812 7837 20846 7871
rect 23213 7837 23247 7871
rect 23581 7837 23615 7871
rect 24409 7837 24443 7871
rect 25605 7837 25639 7871
rect 26341 7837 26375 7871
rect 26709 7837 26743 7871
rect 29561 7837 29595 7871
rect 29724 7837 29758 7871
rect 29840 7834 29874 7868
rect 29949 7837 29983 7871
rect 31217 7837 31251 7871
rect 33793 7837 33827 7871
rect 33882 7837 33916 7871
rect 33977 7831 34011 7865
rect 34161 7837 34195 7871
rect 37933 7837 37967 7871
rect 38096 7837 38130 7871
rect 38212 7837 38246 7871
rect 38301 7837 38335 7871
rect 39037 7837 39071 7871
rect 68109 7837 68143 7871
rect 2145 7769 2179 7803
rect 7389 7769 7423 7803
rect 10517 7769 10551 7803
rect 15678 7769 15712 7803
rect 23397 7769 23431 7803
rect 23489 7769 23523 7803
rect 26525 7769 26559 7803
rect 26617 7769 26651 7803
rect 31484 7769 31518 7803
rect 33517 7769 33551 7803
rect 38577 7769 38611 7803
rect 40110 7769 40144 7803
rect 1685 7701 1719 7735
rect 2973 7701 3007 7735
rect 4353 7701 4387 7735
rect 6837 7701 6871 7735
rect 11069 7701 11103 7735
rect 12173 7701 12207 7735
rect 14565 7701 14599 7735
rect 19349 7701 19383 7735
rect 24593 7701 24627 7735
rect 30205 7701 30239 7735
rect 32597 7701 32631 7735
rect 34713 7701 34747 7735
rect 2329 7497 2363 7531
rect 4353 7497 4387 7531
rect 5273 7497 5307 7531
rect 8585 7497 8619 7531
rect 14933 7497 14967 7531
rect 16957 7497 16991 7531
rect 23857 7497 23891 7531
rect 27905 7497 27939 7531
rect 28917 7497 28951 7531
rect 29745 7497 29779 7531
rect 33609 7497 33643 7531
rect 37381 7497 37415 7531
rect 39037 7497 39071 7531
rect 3218 7429 3252 7463
rect 8217 7429 8251 7463
rect 10977 7429 11011 7463
rect 18705 7429 18739 7463
rect 24501 7429 24535 7463
rect 27537 7429 27571 7463
rect 27629 7429 27663 7463
rect 28641 7429 28675 7463
rect 30858 7429 30892 7463
rect 33793 7429 33827 7463
rect 34805 7429 34839 7463
rect 36185 7429 36219 7463
rect 2145 7361 2179 7395
rect 5457 7361 5491 7395
rect 7021 7361 7055 7395
rect 8125 7361 8159 7395
rect 8401 7361 8435 7395
rect 9045 7361 9079 7395
rect 10793 7361 10827 7395
rect 11805 7361 11839 7395
rect 13001 7361 13035 7395
rect 13645 7361 13679 7395
rect 14289 7361 14323 7395
rect 14473 7361 14507 7395
rect 14565 7361 14599 7395
rect 14657 7361 14691 7395
rect 16681 7361 16715 7395
rect 16865 7361 16899 7395
rect 18521 7361 18555 7395
rect 18797 7361 18831 7395
rect 22661 7361 22695 7395
rect 24317 7361 24351 7395
rect 25375 7361 25409 7395
rect 25510 7361 25544 7395
rect 25626 7361 25660 7395
rect 25789 7361 25823 7395
rect 27353 7361 27387 7395
rect 27721 7361 27755 7395
rect 28365 7361 28399 7395
rect 28549 7361 28583 7395
rect 28733 7361 28767 7395
rect 33977 7361 34011 7395
rect 34621 7361 34655 7395
rect 36001 7361 36035 7395
rect 36093 7361 36127 7395
rect 36369 7361 36403 7395
rect 37933 7361 37967 7395
rect 38117 7361 38151 7395
rect 38212 7361 38246 7395
rect 38301 7361 38335 7395
rect 1685 7293 1719 7327
rect 2973 7293 3007 7327
rect 5641 7293 5675 7327
rect 9321 7293 9355 7327
rect 11529 7293 11563 7327
rect 18337 7293 18371 7327
rect 19809 7293 19843 7327
rect 22385 7293 22419 7327
rect 31125 7293 31159 7327
rect 7205 7225 7239 7259
rect 13829 7225 13863 7259
rect 24685 7225 24719 7259
rect 35817 7225 35851 7259
rect 6469 7157 6503 7191
rect 13185 7157 13219 7191
rect 15393 7157 15427 7191
rect 16129 7157 16163 7191
rect 17601 7157 17635 7191
rect 19349 7157 19383 7191
rect 25145 7157 25179 7191
rect 26341 7157 26375 7191
rect 34437 7157 34471 7191
rect 38577 7157 38611 7191
rect 2053 6953 2087 6987
rect 6377 6953 6411 6987
rect 33425 6953 33459 6987
rect 36737 6953 36771 6987
rect 38209 6953 38243 6987
rect 9873 6885 9907 6919
rect 1685 6817 1719 6851
rect 3249 6817 3283 6851
rect 6837 6817 6871 6851
rect 6929 6817 6963 6851
rect 8125 6817 8159 6851
rect 10609 6817 10643 6851
rect 12173 6817 12207 6851
rect 14565 6817 14599 6851
rect 16313 6817 16347 6851
rect 18613 6817 18647 6851
rect 20545 6817 20579 6851
rect 22661 6817 22695 6851
rect 32045 6817 32079 6851
rect 39865 6817 39899 6851
rect 1869 6749 1903 6783
rect 2697 6749 2731 6783
rect 7665 6749 7699 6783
rect 7941 6749 7975 6783
rect 9137 6749 9171 6783
rect 9321 6749 9355 6783
rect 9413 6749 9447 6783
rect 9505 6749 9539 6783
rect 9689 6749 9723 6783
rect 10333 6749 10367 6783
rect 10517 6749 10551 6783
rect 10701 6749 10735 6783
rect 10885 6749 10919 6783
rect 12909 6749 12943 6783
rect 13553 6749 13587 6783
rect 15209 6749 15243 6783
rect 15853 6749 15887 6783
rect 18521 6749 18555 6783
rect 18705 6749 18739 6783
rect 19441 6749 19475 6783
rect 19625 6749 19659 6783
rect 19717 6749 19751 6783
rect 19809 6749 19843 6783
rect 22385 6749 22419 6783
rect 25789 6749 25823 6783
rect 26433 6749 26467 6783
rect 26617 6749 26651 6783
rect 26709 6749 26743 6783
rect 26801 6749 26835 6783
rect 29561 6749 29595 6783
rect 29745 6749 29779 6783
rect 34713 6749 34747 6783
rect 35357 6749 35391 6783
rect 37381 6749 37415 6783
rect 37565 6749 37599 6783
rect 37749 6749 37783 6783
rect 38577 6749 38611 6783
rect 40121 6749 40155 6783
rect 4169 6681 4203 6715
rect 11989 6681 12023 6715
rect 16580 6681 16614 6715
rect 20085 6681 20119 6715
rect 20790 6681 20824 6715
rect 24961 6681 24995 6715
rect 25605 6681 25639 6715
rect 25973 6681 26007 6715
rect 32312 6681 32346 6715
rect 35602 6681 35636 6715
rect 37473 6681 37507 6715
rect 38393 6681 38427 6715
rect 5457 6613 5491 6647
rect 6745 6613 6779 6647
rect 7757 6613 7791 6647
rect 11069 6613 11103 6647
rect 17693 6613 17727 6647
rect 21925 6613 21959 6647
rect 23765 6613 23799 6647
rect 25053 6613 25087 6647
rect 27077 6613 27111 6647
rect 28917 6613 28951 6647
rect 29929 6613 29963 6647
rect 34897 6613 34931 6647
rect 37197 6613 37231 6647
rect 41245 6613 41279 6647
rect 4169 6409 4203 6443
rect 5273 6409 5307 6443
rect 8401 6409 8435 6443
rect 18337 6409 18371 6443
rect 19625 6409 19659 6443
rect 23673 6409 23707 6443
rect 26433 6409 26467 6443
rect 30205 6409 30239 6443
rect 33609 6409 33643 6443
rect 35173 6409 35207 6443
rect 5181 6341 5215 6375
rect 11774 6341 11808 6375
rect 17049 6341 17083 6375
rect 19257 6341 19291 6375
rect 24133 6341 24167 6375
rect 28190 6341 28224 6375
rect 33149 6341 33183 6375
rect 36277 6341 36311 6375
rect 36461 6341 36495 6375
rect 36645 6341 36679 6375
rect 37473 6341 37507 6375
rect 1777 6273 1811 6307
rect 1869 6273 1903 6307
rect 2789 6273 2823 6307
rect 3056 6273 3090 6307
rect 7021 6273 7055 6307
rect 7297 6273 7331 6307
rect 7941 6273 7975 6307
rect 8033 6273 8067 6307
rect 8217 6273 8251 6307
rect 9873 6273 9907 6307
rect 10977 6273 11011 6307
rect 13369 6273 13403 6307
rect 13636 6273 13670 6307
rect 15209 6273 15243 6307
rect 15393 6273 15427 6307
rect 15577 6273 15611 6307
rect 15761 6273 15795 6307
rect 15945 6273 15979 6307
rect 19441 6273 19475 6307
rect 20729 6273 20763 6307
rect 22293 6273 22327 6307
rect 22560 6273 22594 6307
rect 25881 6273 25915 6307
rect 29101 6273 29135 6307
rect 29264 6273 29298 6307
rect 29377 6273 29411 6307
rect 29469 6273 29503 6307
rect 31318 6273 31352 6307
rect 33885 6273 33919 6307
rect 33977 6273 34011 6307
rect 34069 6273 34103 6307
rect 34253 6273 34287 6307
rect 35449 6273 35483 6307
rect 35541 6273 35575 6307
rect 35633 6273 35667 6307
rect 35817 6273 35851 6307
rect 37289 6273 37323 6307
rect 38117 6273 38151 6307
rect 38301 6273 38335 6307
rect 38393 6273 38427 6307
rect 38485 6273 38519 6307
rect 5365 6205 5399 6239
rect 9597 6205 9631 6239
rect 11529 6205 11563 6239
rect 15669 6205 15703 6239
rect 28457 6205 28491 6239
rect 31585 6205 31619 6239
rect 37657 6205 37691 6239
rect 4813 6137 4847 6171
rect 14749 6137 14783 6171
rect 27077 6137 27111 6171
rect 29745 6137 29779 6171
rect 67649 6137 67683 6171
rect 2053 6069 2087 6103
rect 10793 6069 10827 6103
rect 12909 6069 12943 6103
rect 20085 6069 20119 6103
rect 20913 6069 20947 6103
rect 38761 6069 38795 6103
rect 2145 5865 2179 5899
rect 3249 5865 3283 5899
rect 5457 5865 5491 5899
rect 15669 5865 15703 5899
rect 16681 5865 16715 5899
rect 17877 5865 17911 5899
rect 23489 5865 23523 5899
rect 25697 5865 25731 5899
rect 26525 5865 26559 5899
rect 29009 5865 29043 5899
rect 30481 5865 30515 5899
rect 36001 5865 36035 5899
rect 38301 5865 38335 5899
rect 1501 5797 1535 5831
rect 6101 5797 6135 5831
rect 15209 5797 15243 5831
rect 27629 5797 27663 5831
rect 30941 5797 30975 5831
rect 36553 5797 36587 5831
rect 4905 5729 4939 5763
rect 17049 5729 17083 5763
rect 19809 5729 19843 5763
rect 21373 5729 21407 5763
rect 22109 5729 22143 5763
rect 35265 5729 35299 5763
rect 1961 5661 1995 5695
rect 3985 5661 4019 5695
rect 5917 5661 5951 5695
rect 7849 5661 7883 5695
rect 8125 5661 8159 5695
rect 9045 5661 9079 5695
rect 12173 5661 12207 5695
rect 12429 5661 12463 5695
rect 14105 5661 14139 5695
rect 15025 5661 15059 5695
rect 15853 5661 15887 5695
rect 16129 5661 16163 5695
rect 16865 5661 16899 5695
rect 17141 5661 17175 5695
rect 17233 5661 17267 5695
rect 17417 5661 17451 5695
rect 18061 5661 18095 5695
rect 18337 5661 18371 5695
rect 19625 5661 19659 5695
rect 21649 5661 21683 5695
rect 24869 5661 24903 5695
rect 28825 5661 28859 5695
rect 29837 5661 29871 5695
rect 30021 5658 30055 5692
rect 30113 5661 30147 5695
rect 30251 5661 30285 5695
rect 31953 5661 31987 5695
rect 34161 5661 34195 5695
rect 35541 5661 35575 5695
rect 37105 5661 37139 5695
rect 37289 5661 37323 5695
rect 37381 5661 37415 5695
rect 37473 5661 37507 5695
rect 2697 5593 2731 5627
rect 6653 5593 6687 5627
rect 9965 5593 9999 5627
rect 11713 5593 11747 5627
rect 18245 5593 18279 5627
rect 22376 5593 22410 5627
rect 25053 5593 25087 5627
rect 25605 5593 25639 5627
rect 26433 5593 26467 5627
rect 28641 5593 28675 5627
rect 32413 5593 32447 5627
rect 3801 5525 3835 5559
rect 6745 5525 6779 5559
rect 9137 5525 9171 5559
rect 13553 5525 13587 5559
rect 14289 5525 14323 5559
rect 16037 5525 16071 5559
rect 19257 5525 19291 5559
rect 19717 5525 19751 5559
rect 24685 5525 24719 5559
rect 27077 5525 27111 5559
rect 37749 5525 37783 5559
rect 3801 5321 3835 5355
rect 8125 5321 8159 5355
rect 9505 5321 9539 5355
rect 14473 5321 14507 5355
rect 17141 5321 17175 5355
rect 17509 5321 17543 5355
rect 23305 5321 23339 5355
rect 29837 5321 29871 5355
rect 32413 5321 32447 5355
rect 35081 5321 35115 5355
rect 37657 5321 37691 5355
rect 40325 5321 40359 5355
rect 3249 5253 3283 5287
rect 6837 5253 6871 5287
rect 7757 5253 7791 5287
rect 13737 5253 13771 5287
rect 26065 5253 26099 5287
rect 27353 5253 27387 5287
rect 37473 5253 37507 5287
rect 39190 5253 39224 5287
rect 2237 5185 2271 5219
rect 4997 5185 5031 5219
rect 5457 5185 5491 5219
rect 5641 5185 5675 5219
rect 7665 5185 7699 5219
rect 7941 5185 7975 5219
rect 9505 5185 9539 5219
rect 9781 5185 9815 5219
rect 10057 5185 10091 5219
rect 10977 5185 11011 5219
rect 12173 5185 12207 5219
rect 12633 5185 12667 5219
rect 12909 5185 12943 5219
rect 14197 5185 14231 5219
rect 15209 5185 15243 5219
rect 17325 5185 17359 5219
rect 17585 5185 17619 5219
rect 18337 5185 18371 5219
rect 19165 5185 19199 5219
rect 19349 5185 19383 5219
rect 19809 5185 19843 5219
rect 22017 5185 22051 5219
rect 23581 5185 23615 5219
rect 23670 5188 23704 5222
rect 23770 5185 23804 5219
rect 23949 5185 23983 5219
rect 24593 5185 24627 5219
rect 24777 5185 24811 5219
rect 24869 5185 24903 5219
rect 24961 5185 24995 5219
rect 26249 5185 26283 5219
rect 27537 5185 27571 5219
rect 30950 5185 30984 5219
rect 31217 5185 31251 5219
rect 33149 5185 33183 5219
rect 33241 5185 33275 5219
rect 33333 5185 33367 5219
rect 33517 5185 33551 5219
rect 34253 5185 34287 5219
rect 34345 5185 34379 5219
rect 34437 5185 34471 5219
rect 34621 5185 34655 5219
rect 36093 5185 36127 5219
rect 36185 5185 36219 5219
rect 36277 5185 36311 5219
rect 36461 5185 36495 5219
rect 37289 5185 37323 5219
rect 5825 5117 5859 5151
rect 6929 5117 6963 5151
rect 7113 5117 7147 5151
rect 11897 5117 11931 5151
rect 12817 5117 12851 5151
rect 14289 5117 14323 5151
rect 18981 5117 19015 5151
rect 20453 5117 20487 5151
rect 20729 5117 20763 5151
rect 38945 5117 38979 5151
rect 59461 5117 59495 5151
rect 1777 5049 1811 5083
rect 4353 5049 4387 5083
rect 6469 5049 6503 5083
rect 9045 5049 9079 5083
rect 11621 5049 11655 5083
rect 13737 5049 13771 5083
rect 60105 5049 60139 5083
rect 2421 4981 2455 5015
rect 4813 4981 4847 5015
rect 10793 4981 10827 5015
rect 12081 4981 12115 5015
rect 12633 4981 12667 5015
rect 13093 4981 13127 5015
rect 15025 4981 15059 5015
rect 16129 4981 16163 5015
rect 18521 4981 18555 5015
rect 19993 4981 20027 5015
rect 21833 4981 21867 5015
rect 22753 4981 22787 5015
rect 25237 4981 25271 5015
rect 26433 4981 26467 5015
rect 27721 4981 27755 5015
rect 32873 4981 32907 5015
rect 33977 4981 34011 5015
rect 35817 4981 35851 5015
rect 58817 4981 58851 5015
rect 67649 4981 67683 5015
rect 5825 4777 5859 4811
rect 9413 4777 9447 4811
rect 10609 4777 10643 4811
rect 11989 4777 12023 4811
rect 14473 4777 14507 4811
rect 14933 4777 14967 4811
rect 20637 4777 20671 4811
rect 23489 4777 23523 4811
rect 27169 4777 27203 4811
rect 27629 4777 27663 4811
rect 32781 4777 32815 4811
rect 33885 4777 33919 4811
rect 34713 4777 34747 4811
rect 36185 4777 36219 4811
rect 37381 4777 37415 4811
rect 1593 4709 1627 4743
rect 6469 4709 6503 4743
rect 11694 4709 11728 4743
rect 11805 4709 11839 4743
rect 14105 4709 14139 4743
rect 14565 4709 14599 4743
rect 18705 4709 18739 4743
rect 21097 4709 21131 4743
rect 25237 4709 25271 4743
rect 57897 4709 57931 4743
rect 59185 4709 59219 4743
rect 2605 4641 2639 4675
rect 7481 4641 7515 4675
rect 10333 4641 10367 4675
rect 11897 4641 11931 4675
rect 14657 4641 14691 4675
rect 15945 4641 15979 4675
rect 16037 4641 16071 4675
rect 16865 4641 16899 4675
rect 18061 4641 18095 4675
rect 18245 4641 18279 4675
rect 22477 4641 22511 4675
rect 25789 4641 25823 4675
rect 29009 4641 29043 4675
rect 38761 4641 38795 4675
rect 60473 4641 60507 4675
rect 1409 4573 1443 4607
rect 3801 4573 3835 4607
rect 4445 4573 4479 4607
rect 4712 4573 4746 4607
rect 8217 4573 8251 4607
rect 8953 4573 8987 4607
rect 9321 4573 9355 4607
rect 9505 4573 9539 4607
rect 10241 4573 10275 4607
rect 12725 4573 12759 4607
rect 13001 4573 13035 4607
rect 17509 4573 17543 4607
rect 19257 4573 19291 4607
rect 22210 4573 22244 4607
rect 23121 4573 23155 4607
rect 23305 4573 23339 4607
rect 26045 4573 26079 4607
rect 32965 4573 32999 4607
rect 34897 4573 34931 4607
rect 36001 4573 36035 4607
rect 38494 4573 38528 4607
rect 57253 4573 57287 4607
rect 58541 4573 58575 4607
rect 2513 4505 2547 4539
rect 6653 4505 6687 4539
rect 7297 4505 7331 4539
rect 10701 4505 10735 4539
rect 11529 4505 11563 4539
rect 19524 4505 19558 4539
rect 24409 4505 24443 4539
rect 28742 4505 28776 4539
rect 33149 4505 33183 4539
rect 35081 4505 35115 4539
rect 35817 4505 35851 4539
rect 2053 4437 2087 4471
rect 2421 4437 2455 4471
rect 3985 4437 4019 4471
rect 8401 4437 8435 4471
rect 9137 4437 9171 4471
rect 10057 4437 10091 4471
rect 15485 4437 15519 4471
rect 15853 4437 15887 4471
rect 18337 4437 18371 4471
rect 2145 4233 2179 4267
rect 5181 4233 5215 4267
rect 7573 4233 7607 4267
rect 9597 4233 9631 4267
rect 10609 4233 10643 4267
rect 19533 4233 19567 4267
rect 20085 4233 20119 4267
rect 34897 4233 34931 4267
rect 36737 4233 36771 4267
rect 3126 4165 3160 4199
rect 10977 4165 11011 4199
rect 1961 4097 1995 4131
rect 4997 4097 5031 4131
rect 5641 4097 5675 4131
rect 6561 4097 6595 4131
rect 7665 4097 7699 4131
rect 8861 4097 8895 4131
rect 9137 4097 9171 4131
rect 9781 4097 9815 4131
rect 10793 4097 10827 4131
rect 14381 4097 14415 4131
rect 15393 4097 15427 4131
rect 15577 4097 15611 4131
rect 17794 4097 17828 4131
rect 18061 4097 18095 4131
rect 18705 4097 18739 4131
rect 18889 4097 18923 4131
rect 19349 4097 19383 4131
rect 23213 4097 23247 4131
rect 23376 4103 23410 4137
rect 23476 4103 23510 4137
rect 23627 4097 23661 4131
rect 24317 4097 24351 4131
rect 24573 4097 24607 4131
rect 27353 4097 27387 4131
rect 27537 4097 27571 4131
rect 27629 4097 27663 4131
rect 27721 4097 27755 4131
rect 30674 4097 30708 4131
rect 30941 4097 30975 4131
rect 33517 4097 33551 4131
rect 33784 4097 33818 4131
rect 35357 4097 35391 4131
rect 35624 4097 35658 4131
rect 59829 4097 59863 4131
rect 1777 4029 1811 4063
rect 2881 4029 2915 4063
rect 6745 4029 6779 4063
rect 7849 4029 7883 4063
rect 9965 4029 9999 4063
rect 12357 4029 12391 4063
rect 12725 4029 12759 4063
rect 13461 4029 13495 4063
rect 14013 4029 14047 4063
rect 15761 4029 15795 4063
rect 18521 4029 18555 4063
rect 23857 4029 23891 4063
rect 27997 4029 28031 4063
rect 61117 4029 61151 4063
rect 6377 3961 6411 3995
rect 7205 3961 7239 3995
rect 11805 3961 11839 3995
rect 12265 3961 12299 3995
rect 13921 3961 13955 3995
rect 16681 3961 16715 3995
rect 21833 3961 21867 3995
rect 25697 3961 25731 3995
rect 29561 3961 29595 3995
rect 58541 3961 58575 3995
rect 60473 3961 60507 3995
rect 4261 3893 4295 3927
rect 5825 3893 5859 3927
rect 12173 3893 12207 3927
rect 13829 3893 13863 3927
rect 14933 3893 14967 3927
rect 20545 3893 20579 3927
rect 21189 3893 21223 3927
rect 22477 3893 22511 3927
rect 26341 3893 26375 3927
rect 32689 3893 32723 3927
rect 56241 3893 56275 3927
rect 56885 3893 56919 3927
rect 57897 3893 57931 3927
rect 59185 3893 59219 3927
rect 4169 3689 4203 3723
rect 7757 3689 7791 3723
rect 8953 3689 8987 3723
rect 9321 3689 9355 3723
rect 9965 3689 9999 3723
rect 10793 3689 10827 3723
rect 10977 3689 11011 3723
rect 11805 3689 11839 3723
rect 11897 3689 11931 3723
rect 12265 3689 12299 3723
rect 14289 3689 14323 3723
rect 15025 3689 15059 3723
rect 15761 3689 15795 3723
rect 23489 3689 23523 3723
rect 27169 3689 27203 3723
rect 31769 3689 31803 3723
rect 4905 3621 4939 3655
rect 7297 3621 7331 3655
rect 13369 3621 13403 3655
rect 19349 3621 19383 3655
rect 22017 3621 22051 3655
rect 41797 3621 41831 3655
rect 57897 3621 57931 3655
rect 61117 3621 61151 3655
rect 2421 3553 2455 3587
rect 3801 3553 3835 3587
rect 5457 3553 5491 3587
rect 11437 3553 11471 3587
rect 11989 3553 12023 3587
rect 14381 3553 14415 3587
rect 17325 3553 17359 3587
rect 19809 3553 19843 3587
rect 33149 3553 33183 3587
rect 56609 3553 56643 3587
rect 58541 3553 58575 3587
rect 61761 3553 61795 3587
rect 3065 3485 3099 3519
rect 3985 3485 4019 3519
rect 6469 3485 6503 3519
rect 7113 3485 7147 3519
rect 7941 3485 7975 3519
rect 8125 3485 8159 3519
rect 9137 3485 9171 3519
rect 9321 3485 9355 3519
rect 13553 3485 13587 3519
rect 14473 3485 14507 3519
rect 15209 3485 15243 3519
rect 16681 3485 16715 3519
rect 17877 3485 17911 3519
rect 18705 3485 18739 3519
rect 21097 3485 21131 3519
rect 22661 3485 22695 3519
rect 24777 3485 24811 3519
rect 25421 3485 25455 3519
rect 26065 3485 26099 3519
rect 26525 3485 26559 3519
rect 26709 3485 26743 3519
rect 26801 3485 26835 3519
rect 26939 3485 26973 3519
rect 27997 3485 28031 3519
rect 28825 3485 28859 3519
rect 29653 3485 29687 3519
rect 30665 3485 30699 3519
rect 31125 3485 31159 3519
rect 32882 3485 32916 3519
rect 39865 3485 39899 3519
rect 40509 3485 40543 3519
rect 41153 3485 41187 3519
rect 42625 3485 42659 3519
rect 43269 3485 43303 3519
rect 45109 3485 45143 3519
rect 45753 3485 45787 3519
rect 46397 3485 46431 3519
rect 47041 3485 47075 3519
rect 47869 3485 47903 3519
rect 48973 3485 49007 3519
rect 50353 3485 50387 3519
rect 50997 3485 51031 3519
rect 51641 3485 51675 3519
rect 52837 3485 52871 3519
rect 53481 3485 53515 3519
rect 55321 3485 55355 3519
rect 55965 3485 55999 3519
rect 57253 3485 57287 3519
rect 59185 3485 59219 3519
rect 60473 3485 60507 3519
rect 68109 3485 68143 3519
rect 2329 3417 2363 3451
rect 9781 3417 9815 3451
rect 9997 3417 10031 3451
rect 10609 3417 10643 3451
rect 15853 3417 15887 3451
rect 19349 3417 19383 3451
rect 19901 3417 19935 3451
rect 20085 3417 20119 3451
rect 23121 3417 23155 3451
rect 23305 3417 23339 3451
rect 1869 3349 1903 3383
rect 2237 3349 2271 3383
rect 3249 3349 3283 3383
rect 5273 3349 5307 3383
rect 5365 3349 5399 3383
rect 6653 3349 6687 3383
rect 10149 3349 10183 3383
rect 10809 3349 10843 3383
rect 14105 3349 14139 3383
rect 16497 3349 16531 3383
rect 18061 3349 18095 3383
rect 20545 3349 20579 3383
rect 1593 3145 1627 3179
rect 3985 3145 4019 3179
rect 5825 3145 5859 3179
rect 7757 3145 7791 3179
rect 12541 3145 12575 3179
rect 18705 3145 18739 3179
rect 21925 3145 21959 3179
rect 26985 3145 27019 3179
rect 4712 3077 4746 3111
rect 10517 3077 10551 3111
rect 13093 3077 13127 3111
rect 1777 3009 1811 3043
rect 1961 3009 1995 3043
rect 2605 3009 2639 3043
rect 2872 3009 2906 3043
rect 4445 3009 4479 3043
rect 6377 3009 6411 3043
rect 6633 3009 6667 3043
rect 9606 3009 9640 3043
rect 9873 3009 9907 3043
rect 10885 3009 10919 3043
rect 11897 3009 11931 3043
rect 11989 3009 12023 3043
rect 12357 3009 12391 3043
rect 13553 3009 13587 3043
rect 14473 3009 14507 3043
rect 15485 3009 15519 3043
rect 16957 3009 16991 3043
rect 17601 3009 17635 3043
rect 18521 3009 18555 3043
rect 61117 3009 61151 3043
rect 13369 2941 13403 2975
rect 14197 2941 14231 2975
rect 19993 2941 20027 2975
rect 21281 2941 21315 2975
rect 24501 2941 24535 2975
rect 28365 2941 28399 2975
rect 30297 2941 30331 2975
rect 37933 2941 37967 2975
rect 45661 2941 45695 2975
rect 49525 2941 49559 2975
rect 53389 2941 53423 2975
rect 61761 2941 61795 2975
rect 8493 2873 8527 2907
rect 16773 2873 16807 2907
rect 19349 2873 19383 2907
rect 22569 2873 22603 2907
rect 26433 2873 26467 2907
rect 39221 2873 39255 2907
rect 40509 2873 40543 2907
rect 43085 2873 43119 2907
rect 44373 2873 44407 2907
rect 48237 2873 48271 2907
rect 50169 2873 50203 2907
rect 51457 2873 51491 2907
rect 54033 2873 54067 2907
rect 55321 2873 55355 2907
rect 56609 2873 56643 2907
rect 58541 2873 58575 2907
rect 63049 2873 63083 2907
rect 12357 2805 12391 2839
rect 13185 2805 13219 2839
rect 13737 2805 13771 2839
rect 15669 2805 15703 2839
rect 17509 2805 17543 2839
rect 20637 2805 20671 2839
rect 23213 2805 23247 2839
rect 23857 2805 23891 2839
rect 25145 2805 25179 2839
rect 25789 2805 25823 2839
rect 27721 2805 27755 2839
rect 29009 2805 29043 2839
rect 29653 2805 29687 2839
rect 30941 2805 30975 2839
rect 31585 2805 31619 2839
rect 32873 2805 32907 2839
rect 33517 2805 33551 2839
rect 34161 2805 34195 2839
rect 34621 2805 34655 2839
rect 35449 2805 35483 2839
rect 36277 2805 36311 2839
rect 37289 2805 37323 2839
rect 38577 2805 38611 2839
rect 39865 2805 39899 2839
rect 41153 2805 41187 2839
rect 42441 2805 42475 2839
rect 43729 2805 43763 2839
rect 45017 2805 45051 2839
rect 46305 2805 46339 2839
rect 47593 2805 47627 2839
rect 48881 2805 48915 2839
rect 50813 2805 50847 2839
rect 52745 2805 52779 2839
rect 54677 2805 54711 2839
rect 55965 2805 55999 2839
rect 57897 2805 57931 2839
rect 59185 2805 59219 2839
rect 59829 2805 59863 2839
rect 60473 2805 60507 2839
rect 1961 2601 1995 2635
rect 9873 2601 9907 2635
rect 14841 2601 14875 2635
rect 17509 2601 17543 2635
rect 24409 2601 24443 2635
rect 55321 2601 55355 2635
rect 61117 2601 61151 2635
rect 5641 2533 5675 2567
rect 15945 2533 15979 2567
rect 18337 2533 18371 2567
rect 19993 2533 20027 2567
rect 22569 2533 22603 2567
rect 25789 2533 25823 2567
rect 31585 2533 31619 2567
rect 42441 2533 42475 2567
rect 46305 2533 46339 2567
rect 50169 2533 50203 2567
rect 54033 2533 54067 2567
rect 57897 2533 57931 2567
rect 58541 2533 58575 2567
rect 60473 2533 60507 2567
rect 10609 2465 10643 2499
rect 11805 2465 11839 2499
rect 20637 2465 20671 2499
rect 23213 2465 23247 2499
rect 25145 2465 25179 2499
rect 27721 2465 27755 2499
rect 29009 2465 29043 2499
rect 37933 2465 37967 2499
rect 39865 2465 39899 2499
rect 43085 2465 43119 2499
rect 45017 2465 45051 2499
rect 48237 2465 48271 2499
rect 50813 2465 50847 2499
rect 52745 2465 52779 2499
rect 56609 2465 56643 2499
rect 63693 2465 63727 2499
rect 1777 2397 1811 2431
rect 2421 2397 2455 2431
rect 3065 2397 3099 2431
rect 4261 2397 4295 2431
rect 4905 2397 4939 2431
rect 5825 2397 5859 2431
rect 6929 2397 6963 2431
rect 7665 2397 7699 2431
rect 8401 2397 8435 2431
rect 9137 2397 9171 2431
rect 11529 2397 11563 2431
rect 15761 2397 15795 2431
rect 16957 2397 16991 2431
rect 18153 2397 18187 2431
rect 21281 2397 21315 2431
rect 23857 2397 23891 2431
rect 26433 2397 26467 2431
rect 28365 2397 28399 2431
rect 30297 2397 30331 2431
rect 30941 2397 30975 2431
rect 32873 2397 32907 2431
rect 33517 2397 33551 2431
rect 34161 2397 34195 2431
rect 34897 2397 34931 2431
rect 35541 2397 35575 2431
rect 36001 2397 36035 2431
rect 37289 2397 37323 2431
rect 38577 2397 38611 2431
rect 40509 2397 40543 2431
rect 41153 2397 41187 2431
rect 43729 2397 43763 2431
rect 45661 2397 45695 2431
rect 47593 2397 47627 2431
rect 48881 2397 48915 2431
rect 51457 2397 51491 2431
rect 53389 2397 53423 2431
rect 55965 2397 55999 2431
rect 59185 2397 59219 2431
rect 61761 2397 61795 2431
rect 63049 2397 63083 2431
rect 67005 2397 67039 2431
rect 67649 2397 67683 2431
rect 9965 2329 9999 2363
rect 10885 2329 10919 2363
rect 12909 2329 12943 2363
rect 14565 2329 14599 2363
rect 17601 2329 17635 2363
rect 26985 2329 27019 2363
rect 2605 2261 2639 2295
rect 3249 2261 3283 2295
rect 4445 2261 4479 2295
rect 5089 2261 5123 2295
rect 6745 2261 6779 2295
rect 7481 2261 7515 2295
rect 8217 2261 8251 2295
rect 13001 2261 13035 2295
rect 16773 2261 16807 2295
rect 19349 2261 19383 2295
rect 21833 2261 21867 2295
<< metal1 >>
rect 1104 57690 68816 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 68816 57690
rect 1104 57616 68816 57638
rect 5166 57400 5172 57452
rect 5224 57440 5230 57452
rect 5261 57443 5319 57449
rect 5261 57440 5273 57443
rect 5224 57412 5273 57440
rect 5224 57400 5230 57412
rect 5261 57409 5273 57412
rect 5307 57409 5319 57443
rect 15194 57440 15200 57452
rect 15155 57412 15200 57440
rect 5261 57403 5319 57409
rect 15194 57400 15200 57412
rect 15252 57400 15258 57452
rect 25038 57400 25044 57452
rect 25096 57440 25102 57452
rect 25133 57443 25191 57449
rect 25133 57440 25145 57443
rect 25096 57412 25145 57440
rect 25096 57400 25102 57412
rect 25133 57409 25145 57412
rect 25179 57409 25191 57443
rect 25133 57403 25191 57409
rect 34974 57400 34980 57452
rect 35032 57440 35038 57452
rect 35069 57443 35127 57449
rect 35069 57440 35081 57443
rect 35032 57412 35081 57440
rect 35032 57400 35038 57412
rect 35069 57409 35081 57412
rect 35115 57409 35127 57443
rect 35069 57403 35127 57409
rect 44910 57400 44916 57452
rect 44968 57440 44974 57452
rect 45005 57443 45063 57449
rect 45005 57440 45017 57443
rect 44968 57412 45017 57440
rect 44968 57400 44974 57412
rect 45005 57409 45017 57412
rect 45051 57409 45063 57443
rect 45005 57403 45063 57409
rect 54846 57400 54852 57452
rect 54904 57440 54910 57452
rect 55309 57443 55367 57449
rect 55309 57440 55321 57443
rect 54904 57412 55321 57440
rect 54904 57400 54910 57412
rect 55309 57409 55321 57412
rect 55355 57409 55367 57443
rect 55309 57403 55367 57409
rect 64782 57400 64788 57452
rect 64840 57440 64846 57452
rect 64877 57443 64935 57449
rect 64877 57440 64889 57443
rect 64840 57412 64889 57440
rect 64840 57400 64846 57412
rect 64877 57409 64889 57412
rect 64923 57409 64935 57443
rect 66990 57440 66996 57452
rect 66951 57412 66996 57440
rect 64877 57403 64935 57409
rect 66990 57400 66996 57412
rect 67048 57400 67054 57452
rect 67542 57400 67548 57452
rect 67600 57440 67606 57452
rect 67637 57443 67695 57449
rect 67637 57440 67649 57443
rect 67600 57412 67649 57440
rect 67600 57400 67606 57412
rect 67637 57409 67649 57412
rect 67683 57409 67695 57443
rect 67637 57403 67695 57409
rect 1104 57146 68816 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 65654 57146
rect 65706 57094 65718 57146
rect 65770 57094 65782 57146
rect 65834 57094 65846 57146
rect 65898 57094 65910 57146
rect 65962 57094 68816 57146
rect 1104 57072 68816 57094
rect 68094 56828 68100 56840
rect 68055 56800 68100 56828
rect 68094 56788 68100 56800
rect 68152 56788 68158 56840
rect 1104 56602 68816 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 68816 56602
rect 1104 56528 68816 56550
rect 1104 56058 68816 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 65654 56058
rect 65706 56006 65718 56058
rect 65770 56006 65782 56058
rect 65834 56006 65846 56058
rect 65898 56006 65910 56058
rect 65962 56006 68816 56058
rect 1104 55984 68816 56006
rect 1104 55514 68816 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 68816 55514
rect 1104 55440 68816 55462
rect 67634 55128 67640 55140
rect 67595 55100 67640 55128
rect 67634 55088 67640 55100
rect 67692 55088 67698 55140
rect 1104 54970 68816 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 65654 54970
rect 65706 54918 65718 54970
rect 65770 54918 65782 54970
rect 65834 54918 65846 54970
rect 65898 54918 65910 54970
rect 65962 54918 68816 54970
rect 1104 54896 68816 54918
rect 1104 54426 68816 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 68816 54426
rect 1104 54352 68816 54374
rect 67542 53932 67548 53984
rect 67600 53972 67606 53984
rect 67637 53975 67695 53981
rect 67637 53972 67649 53975
rect 67600 53944 67649 53972
rect 67600 53932 67606 53944
rect 67637 53941 67649 53944
rect 67683 53941 67695 53975
rect 67637 53935 67695 53941
rect 1104 53882 68816 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 65654 53882
rect 65706 53830 65718 53882
rect 65770 53830 65782 53882
rect 65834 53830 65846 53882
rect 65898 53830 65910 53882
rect 65962 53830 68816 53882
rect 1104 53808 68816 53830
rect 1104 53338 68816 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 68816 53338
rect 1104 53264 68816 53286
rect 1104 52794 68816 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 65654 52794
rect 65706 52742 65718 52794
rect 65770 52742 65782 52794
rect 65834 52742 65846 52794
rect 65898 52742 65910 52794
rect 65962 52742 68816 52794
rect 1104 52720 68816 52742
rect 68094 52476 68100 52488
rect 68055 52448 68100 52476
rect 68094 52436 68100 52448
rect 68152 52436 68158 52488
rect 1104 52250 68816 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 68816 52250
rect 1104 52176 68816 52198
rect 1104 51706 68816 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 65654 51706
rect 65706 51654 65718 51706
rect 65770 51654 65782 51706
rect 65834 51654 65846 51706
rect 65898 51654 65910 51706
rect 65962 51654 68816 51706
rect 1104 51632 68816 51654
rect 68094 51388 68100 51400
rect 68055 51360 68100 51388
rect 68094 51348 68100 51360
rect 68152 51348 68158 51400
rect 1104 51162 68816 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 68816 51162
rect 1104 51088 68816 51110
rect 1104 50618 68816 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 65654 50618
rect 65706 50566 65718 50618
rect 65770 50566 65782 50618
rect 65834 50566 65846 50618
rect 65898 50566 65910 50618
rect 65962 50566 68816 50618
rect 1104 50544 68816 50566
rect 1104 50074 68816 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 68816 50074
rect 1104 50000 68816 50022
rect 67634 49756 67640 49768
rect 67595 49728 67640 49756
rect 67634 49716 67640 49728
rect 67692 49716 67698 49768
rect 1104 49530 68816 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 65654 49530
rect 65706 49478 65718 49530
rect 65770 49478 65782 49530
rect 65834 49478 65846 49530
rect 65898 49478 65910 49530
rect 65962 49478 68816 49530
rect 1104 49456 68816 49478
rect 1104 48986 68816 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 68816 48986
rect 1104 48912 68816 48934
rect 67634 48532 67640 48544
rect 67595 48504 67640 48532
rect 67634 48492 67640 48504
rect 67692 48492 67698 48544
rect 1104 48442 68816 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 65654 48442
rect 65706 48390 65718 48442
rect 65770 48390 65782 48442
rect 65834 48390 65846 48442
rect 65898 48390 65910 48442
rect 65962 48390 68816 48442
rect 1104 48368 68816 48390
rect 1104 47898 68816 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 68816 47898
rect 1104 47824 68816 47846
rect 1104 47354 68816 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 65654 47354
rect 65706 47302 65718 47354
rect 65770 47302 65782 47354
rect 65834 47302 65846 47354
rect 65898 47302 65910 47354
rect 65962 47302 68816 47354
rect 1104 47280 68816 47302
rect 68094 47036 68100 47048
rect 68055 47008 68100 47036
rect 68094 46996 68100 47008
rect 68152 46996 68158 47048
rect 1104 46810 68816 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 68816 46810
rect 1104 46736 68816 46758
rect 1104 46266 68816 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 65654 46266
rect 65706 46214 65718 46266
rect 65770 46214 65782 46266
rect 65834 46214 65846 46266
rect 65898 46214 65910 46266
rect 65962 46214 68816 46266
rect 1104 46192 68816 46214
rect 68094 45948 68100 45960
rect 68055 45920 68100 45948
rect 68094 45908 68100 45920
rect 68152 45908 68158 45960
rect 1104 45722 68816 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 68816 45722
rect 1104 45648 68816 45670
rect 1104 45178 68816 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 65654 45178
rect 65706 45126 65718 45178
rect 65770 45126 65782 45178
rect 65834 45126 65846 45178
rect 65898 45126 65910 45178
rect 65962 45126 68816 45178
rect 1104 45104 68816 45126
rect 1104 44634 68816 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 68816 44634
rect 1104 44560 68816 44582
rect 67634 44248 67640 44260
rect 67595 44220 67640 44248
rect 67634 44208 67640 44220
rect 67692 44208 67698 44260
rect 1104 44090 68816 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 65654 44090
rect 65706 44038 65718 44090
rect 65770 44038 65782 44090
rect 65834 44038 65846 44090
rect 65898 44038 65910 44090
rect 65962 44038 68816 44090
rect 1104 44016 68816 44038
rect 1104 43546 68816 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 68816 43546
rect 1104 43472 68816 43494
rect 67634 43092 67640 43104
rect 67595 43064 67640 43092
rect 67634 43052 67640 43064
rect 67692 43052 67698 43104
rect 1104 43002 68816 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 65654 43002
rect 65706 42950 65718 43002
rect 65770 42950 65782 43002
rect 65834 42950 65846 43002
rect 65898 42950 65910 43002
rect 65962 42950 68816 43002
rect 1104 42928 68816 42950
rect 1104 42458 68816 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 68816 42458
rect 1104 42384 68816 42406
rect 1104 41914 68816 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 65654 41914
rect 65706 41862 65718 41914
rect 65770 41862 65782 41914
rect 65834 41862 65846 41914
rect 65898 41862 65910 41914
rect 65962 41862 68816 41914
rect 1104 41840 68816 41862
rect 68094 41596 68100 41608
rect 68055 41568 68100 41596
rect 68094 41556 68100 41568
rect 68152 41556 68158 41608
rect 1104 41370 68816 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 68816 41370
rect 1104 41296 68816 41318
rect 1104 40826 68816 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 65654 40826
rect 65706 40774 65718 40826
rect 65770 40774 65782 40826
rect 65834 40774 65846 40826
rect 65898 40774 65910 40826
rect 65962 40774 68816 40826
rect 1104 40752 68816 40774
rect 68094 40508 68100 40520
rect 68055 40480 68100 40508
rect 68094 40468 68100 40480
rect 68152 40468 68158 40520
rect 1104 40282 68816 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 68816 40282
rect 1104 40208 68816 40230
rect 1104 39738 68816 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 65654 39738
rect 65706 39686 65718 39738
rect 65770 39686 65782 39738
rect 65834 39686 65846 39738
rect 65898 39686 65910 39738
rect 65962 39686 68816 39738
rect 1104 39664 68816 39686
rect 1104 39194 68816 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 68816 39194
rect 1104 39120 68816 39142
rect 67634 38808 67640 38820
rect 67595 38780 67640 38808
rect 67634 38768 67640 38780
rect 67692 38768 67698 38820
rect 1104 38650 68816 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 65654 38650
rect 65706 38598 65718 38650
rect 65770 38598 65782 38650
rect 65834 38598 65846 38650
rect 65898 38598 65910 38650
rect 65962 38598 68816 38650
rect 1104 38576 68816 38598
rect 1104 38106 68816 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 68816 38106
rect 1104 38032 68816 38054
rect 67634 37652 67640 37664
rect 67595 37624 67640 37652
rect 67634 37612 67640 37624
rect 67692 37612 67698 37664
rect 1104 37562 68816 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 65654 37562
rect 65706 37510 65718 37562
rect 65770 37510 65782 37562
rect 65834 37510 65846 37562
rect 65898 37510 65910 37562
rect 65962 37510 68816 37562
rect 1104 37488 68816 37510
rect 1104 37018 68816 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 68816 37018
rect 1104 36944 68816 36966
rect 1104 36474 68816 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 65654 36474
rect 65706 36422 65718 36474
rect 65770 36422 65782 36474
rect 65834 36422 65846 36474
rect 65898 36422 65910 36474
rect 65962 36422 68816 36474
rect 1104 36400 68816 36422
rect 68094 36156 68100 36168
rect 68055 36128 68100 36156
rect 68094 36116 68100 36128
rect 68152 36116 68158 36168
rect 1104 35930 68816 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 68816 35930
rect 1104 35856 68816 35878
rect 1104 35386 68816 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 65654 35386
rect 65706 35334 65718 35386
rect 65770 35334 65782 35386
rect 65834 35334 65846 35386
rect 65898 35334 65910 35386
rect 65962 35334 68816 35386
rect 1104 35312 68816 35334
rect 68094 35068 68100 35080
rect 68055 35040 68100 35068
rect 68094 35028 68100 35040
rect 68152 35028 68158 35080
rect 1104 34842 68816 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 68816 34842
rect 1104 34768 68816 34790
rect 1104 34298 68816 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 65654 34298
rect 65706 34246 65718 34298
rect 65770 34246 65782 34298
rect 65834 34246 65846 34298
rect 65898 34246 65910 34298
rect 65962 34246 68816 34298
rect 1104 34224 68816 34246
rect 1104 33754 68816 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 68816 33754
rect 1104 33680 68816 33702
rect 67634 33368 67640 33380
rect 67595 33340 67640 33368
rect 67634 33328 67640 33340
rect 67692 33328 67698 33380
rect 1104 33210 68816 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 65654 33210
rect 65706 33158 65718 33210
rect 65770 33158 65782 33210
rect 65834 33158 65846 33210
rect 65898 33158 65910 33210
rect 65962 33158 68816 33210
rect 1104 33136 68816 33158
rect 1104 32666 68816 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 68816 32666
rect 1104 32592 68816 32614
rect 21358 32172 21364 32224
rect 21416 32212 21422 32224
rect 22462 32212 22468 32224
rect 21416 32184 22468 32212
rect 21416 32172 21422 32184
rect 22462 32172 22468 32184
rect 22520 32172 22526 32224
rect 67634 32212 67640 32224
rect 67595 32184 67640 32212
rect 67634 32172 67640 32184
rect 67692 32172 67698 32224
rect 1104 32122 68816 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 65654 32122
rect 65706 32070 65718 32122
rect 65770 32070 65782 32122
rect 65834 32070 65846 32122
rect 65898 32070 65910 32122
rect 65962 32070 68816 32122
rect 1104 32048 68816 32070
rect 21818 32008 21824 32020
rect 20548 31980 21824 32008
rect 20548 31813 20576 31980
rect 21818 31968 21824 31980
rect 21876 32008 21882 32020
rect 21876 31980 23152 32008
rect 21876 31968 21882 31980
rect 20901 31943 20959 31949
rect 20901 31909 20913 31943
rect 20947 31940 20959 31943
rect 20947 31912 21885 31940
rect 20947 31909 20959 31912
rect 20901 31903 20959 31909
rect 21358 31872 21364 31884
rect 21319 31844 21364 31872
rect 21358 31832 21364 31844
rect 21416 31832 21422 31884
rect 20533 31807 20591 31813
rect 20533 31773 20545 31807
rect 20579 31773 20591 31807
rect 20533 31767 20591 31773
rect 21591 31807 21649 31813
rect 21591 31773 21603 31807
rect 21637 31773 21649 31807
rect 21591 31767 21649 31773
rect 21726 31807 21784 31813
rect 21857 31810 21885 31912
rect 21726 31773 21738 31807
rect 21772 31804 21784 31807
rect 21842 31804 21900 31810
rect 21772 31773 21785 31804
rect 21726 31767 21785 31773
rect 15102 31736 15108 31748
rect 15063 31708 15108 31736
rect 15102 31696 15108 31708
rect 15160 31696 15166 31748
rect 15286 31736 15292 31748
rect 15247 31708 15292 31736
rect 15286 31696 15292 31708
rect 15344 31696 15350 31748
rect 20717 31739 20775 31745
rect 20717 31705 20729 31739
rect 20763 31736 20775 31739
rect 21358 31736 21364 31748
rect 20763 31708 21364 31736
rect 20763 31705 20775 31708
rect 20717 31699 20775 31705
rect 21358 31696 21364 31708
rect 21416 31696 21422 31748
rect 15473 31671 15531 31677
rect 15473 31637 15485 31671
rect 15519 31668 15531 31671
rect 15562 31668 15568 31680
rect 15519 31640 15568 31668
rect 15519 31637 15531 31640
rect 15473 31631 15531 31637
rect 15562 31628 15568 31640
rect 15620 31628 15626 31680
rect 18506 31628 18512 31680
rect 18564 31668 18570 31680
rect 19337 31671 19395 31677
rect 19337 31668 19349 31671
rect 18564 31640 19349 31668
rect 18564 31628 18570 31640
rect 19337 31637 19349 31640
rect 19383 31668 19395 31671
rect 21606 31668 21634 31767
rect 21757 31736 21785 31767
rect 21842 31770 21854 31804
rect 21888 31770 21900 31804
rect 21842 31764 21900 31770
rect 22005 31807 22063 31813
rect 22005 31773 22017 31807
rect 22051 31804 22063 31807
rect 22370 31804 22376 31816
rect 22051 31776 22376 31804
rect 22051 31773 22063 31776
rect 22005 31767 22063 31773
rect 22370 31764 22376 31776
rect 22428 31764 22434 31816
rect 23124 31813 23152 31980
rect 23109 31807 23167 31813
rect 23109 31773 23121 31807
rect 23155 31773 23167 31807
rect 23290 31804 23296 31816
rect 23251 31776 23296 31804
rect 23109 31767 23167 31773
rect 23290 31764 23296 31776
rect 23348 31764 23354 31816
rect 22186 31736 22192 31748
rect 21757 31708 22192 31736
rect 22186 31696 22192 31708
rect 22244 31696 22250 31748
rect 22557 31739 22615 31745
rect 22557 31705 22569 31739
rect 22603 31736 22615 31739
rect 23566 31736 23572 31748
rect 22603 31708 23572 31736
rect 22603 31705 22615 31708
rect 22557 31699 22615 31705
rect 22572 31668 22600 31699
rect 23566 31696 23572 31708
rect 23624 31696 23630 31748
rect 19383 31640 22600 31668
rect 19383 31637 19395 31640
rect 19337 31631 19395 31637
rect 23382 31628 23388 31680
rect 23440 31668 23446 31680
rect 23477 31671 23535 31677
rect 23477 31668 23489 31671
rect 23440 31640 23489 31668
rect 23440 31628 23446 31640
rect 23477 31637 23489 31640
rect 23523 31637 23535 31671
rect 23477 31631 23535 31637
rect 1104 31578 68816 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 68816 31578
rect 1104 31504 68816 31526
rect 12618 31356 12624 31408
rect 12676 31396 12682 31408
rect 12989 31399 13047 31405
rect 12989 31396 13001 31399
rect 12676 31368 13001 31396
rect 12676 31356 12682 31368
rect 12989 31365 13001 31368
rect 13035 31365 13047 31399
rect 15930 31396 15936 31408
rect 12989 31359 13047 31365
rect 15488 31368 15936 31396
rect 3418 31288 3424 31340
rect 3476 31328 3482 31340
rect 3982 31331 4040 31337
rect 3982 31328 3994 31331
rect 3476 31300 3994 31328
rect 3476 31288 3482 31300
rect 3982 31297 3994 31300
rect 4028 31297 4040 31331
rect 3982 31291 4040 31297
rect 12434 31288 12440 31340
rect 12492 31328 12498 31340
rect 12805 31331 12863 31337
rect 12805 31328 12817 31331
rect 12492 31300 12817 31328
rect 12492 31288 12498 31300
rect 12805 31297 12817 31300
rect 12851 31328 12863 31331
rect 15102 31328 15108 31340
rect 12851 31300 15108 31328
rect 12851 31297 12863 31300
rect 12805 31291 12863 31297
rect 15102 31288 15108 31300
rect 15160 31288 15166 31340
rect 15488 31337 15516 31368
rect 15930 31356 15936 31368
rect 15988 31396 15994 31408
rect 15988 31368 19656 31396
rect 15988 31356 15994 31368
rect 15381 31331 15439 31337
rect 15381 31297 15393 31331
rect 15427 31297 15439 31331
rect 15381 31291 15439 31297
rect 15473 31331 15531 31337
rect 15473 31297 15485 31331
rect 15519 31297 15531 31331
rect 15473 31291 15531 31297
rect 4249 31263 4307 31269
rect 4249 31229 4261 31263
rect 4295 31260 4307 31263
rect 4798 31260 4804 31272
rect 4295 31232 4804 31260
rect 4295 31229 4307 31232
rect 4249 31223 4307 31229
rect 4798 31220 4804 31232
rect 4856 31220 4862 31272
rect 15396 31260 15424 31291
rect 15562 31288 15568 31340
rect 15620 31328 15626 31340
rect 15620 31300 15665 31328
rect 15620 31288 15626 31300
rect 15746 31288 15752 31340
rect 15804 31328 15810 31340
rect 17402 31328 17408 31340
rect 15804 31300 15849 31328
rect 17363 31300 17408 31328
rect 15804 31288 15810 31300
rect 17402 31288 17408 31300
rect 17460 31288 17466 31340
rect 17586 31328 17592 31340
rect 17547 31300 17592 31328
rect 17586 31288 17592 31300
rect 17644 31288 17650 31340
rect 18506 31328 18512 31340
rect 18467 31300 18512 31328
rect 18506 31288 18512 31300
rect 18564 31288 18570 31340
rect 18616 31337 18644 31368
rect 18601 31331 18659 31337
rect 18601 31297 18613 31331
rect 18647 31297 18659 31331
rect 18601 31291 18659 31297
rect 18693 31331 18751 31337
rect 18693 31297 18705 31331
rect 18739 31297 18751 31331
rect 18693 31291 18751 31297
rect 18877 31331 18935 31337
rect 18877 31297 18889 31331
rect 18923 31328 18935 31331
rect 19337 31331 19395 31337
rect 19337 31328 19349 31331
rect 18923 31300 19349 31328
rect 18923 31297 18935 31300
rect 18877 31291 18935 31297
rect 19337 31297 19349 31300
rect 19383 31297 19395 31331
rect 19518 31328 19524 31340
rect 19479 31300 19524 31328
rect 19337 31291 19395 31297
rect 17773 31263 17831 31269
rect 15396 31232 16804 31260
rect 15654 31192 15660 31204
rect 12406 31164 15660 31192
rect 2866 31124 2872 31136
rect 2779 31096 2872 31124
rect 2866 31084 2872 31096
rect 2924 31124 2930 31136
rect 12406 31124 12434 31164
rect 15654 31152 15660 31164
rect 15712 31152 15718 31204
rect 16776 31201 16804 31232
rect 17773 31229 17785 31263
rect 17819 31260 17831 31263
rect 18708 31260 18736 31291
rect 17819 31232 18736 31260
rect 19352 31260 19380 31291
rect 19518 31288 19524 31300
rect 19576 31288 19582 31340
rect 19628 31337 19656 31368
rect 19613 31331 19671 31337
rect 19613 31297 19625 31331
rect 19659 31297 19671 31331
rect 19613 31291 19671 31297
rect 19705 31331 19763 31337
rect 19705 31297 19717 31331
rect 19751 31328 19763 31331
rect 22278 31328 22284 31340
rect 19751 31300 22284 31328
rect 19751 31297 19763 31300
rect 19705 31291 19763 31297
rect 22278 31288 22284 31300
rect 22336 31288 22342 31340
rect 22370 31288 22376 31340
rect 22428 31328 22434 31340
rect 23474 31328 23480 31340
rect 22428 31300 23480 31328
rect 22428 31288 22434 31300
rect 23474 31288 23480 31300
rect 23532 31288 23538 31340
rect 23661 31331 23719 31337
rect 23661 31297 23673 31331
rect 23707 31297 23719 31331
rect 23772 31331 23830 31337
rect 23772 31328 23784 31331
rect 23661 31291 23719 31297
rect 23768 31297 23784 31328
rect 23818 31297 23830 31331
rect 23768 31291 23830 31297
rect 23865 31331 23923 31337
rect 23865 31297 23877 31331
rect 23911 31328 23923 31331
rect 23911 31300 23980 31328
rect 23911 31297 23923 31300
rect 23865 31291 23923 31297
rect 20070 31260 20076 31272
rect 19352 31232 20076 31260
rect 17819 31229 17831 31232
rect 17773 31223 17831 31229
rect 20070 31220 20076 31232
rect 20128 31220 20134 31272
rect 23382 31220 23388 31272
rect 23440 31260 23446 31272
rect 23676 31260 23704 31291
rect 23440 31232 23704 31260
rect 23440 31220 23446 31232
rect 16761 31195 16819 31201
rect 16761 31161 16773 31195
rect 16807 31192 16819 31195
rect 16807 31164 22140 31192
rect 16807 31161 16819 31164
rect 16761 31155 16819 31161
rect 2924 31096 12434 31124
rect 13173 31127 13231 31133
rect 2924 31084 2930 31096
rect 13173 31093 13185 31127
rect 13219 31124 13231 31127
rect 13630 31124 13636 31136
rect 13219 31096 13636 31124
rect 13219 31093 13231 31096
rect 13173 31087 13231 31093
rect 13630 31084 13636 31096
rect 13688 31084 13694 31136
rect 15102 31124 15108 31136
rect 15063 31096 15108 31124
rect 15102 31084 15108 31096
rect 15160 31084 15166 31136
rect 15194 31084 15200 31136
rect 15252 31124 15258 31136
rect 17402 31124 17408 31136
rect 15252 31096 17408 31124
rect 15252 31084 15258 31096
rect 17402 31084 17408 31096
rect 17460 31084 17466 31136
rect 18230 31124 18236 31136
rect 18191 31096 18236 31124
rect 18230 31084 18236 31096
rect 18288 31084 18294 31136
rect 19978 31124 19984 31136
rect 19939 31096 19984 31124
rect 19978 31084 19984 31096
rect 20036 31084 20042 31136
rect 22112 31124 22140 31164
rect 22186 31152 22192 31204
rect 22244 31192 22250 31204
rect 23768 31192 23796 31291
rect 22244 31164 23796 31192
rect 22244 31152 22250 31164
rect 23952 31124 23980 31300
rect 24121 31195 24179 31201
rect 24121 31161 24133 31195
rect 24167 31192 24179 31195
rect 25590 31192 25596 31204
rect 24167 31164 25596 31192
rect 24167 31161 24179 31164
rect 24121 31155 24179 31161
rect 25590 31152 25596 31164
rect 25648 31152 25654 31204
rect 24581 31127 24639 31133
rect 24581 31124 24593 31127
rect 22112 31096 24593 31124
rect 24581 31093 24593 31096
rect 24627 31124 24639 31127
rect 24854 31124 24860 31136
rect 24627 31096 24860 31124
rect 24627 31093 24639 31096
rect 24581 31087 24639 31093
rect 24854 31084 24860 31096
rect 24912 31084 24918 31136
rect 1104 31034 68816 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 65654 31034
rect 65706 30982 65718 31034
rect 65770 30982 65782 31034
rect 65834 30982 65846 31034
rect 65898 30982 65910 31034
rect 65962 30982 68816 31034
rect 1104 30960 68816 30982
rect 15286 30880 15292 30932
rect 15344 30920 15350 30932
rect 15473 30923 15531 30929
rect 15473 30920 15485 30923
rect 15344 30892 15485 30920
rect 15344 30880 15350 30892
rect 15473 30889 15485 30892
rect 15519 30889 15531 30923
rect 15473 30883 15531 30889
rect 19518 30880 19524 30932
rect 19576 30920 19582 30932
rect 19613 30923 19671 30929
rect 19613 30920 19625 30923
rect 19576 30892 19625 30920
rect 19576 30880 19582 30892
rect 19613 30889 19625 30892
rect 19659 30889 19671 30923
rect 19613 30883 19671 30889
rect 17402 30744 17408 30796
rect 17460 30784 17466 30796
rect 17460 30756 19288 30784
rect 17460 30744 17466 30756
rect 6730 30716 6736 30728
rect 6691 30688 6736 30716
rect 6730 30676 6736 30688
rect 6788 30676 6794 30728
rect 11054 30676 11060 30728
rect 11112 30716 11118 30728
rect 11425 30719 11483 30725
rect 11425 30716 11437 30719
rect 11112 30688 11437 30716
rect 11112 30676 11118 30688
rect 11425 30685 11437 30688
rect 11471 30685 11483 30719
rect 11425 30679 11483 30685
rect 13814 30676 13820 30728
rect 13872 30716 13878 30728
rect 14093 30719 14151 30725
rect 14093 30716 14105 30719
rect 13872 30688 14105 30716
rect 13872 30676 13878 30688
rect 14093 30685 14105 30688
rect 14139 30716 14151 30719
rect 16393 30719 16451 30725
rect 16393 30716 16405 30719
rect 14139 30688 16405 30716
rect 14139 30685 14151 30688
rect 14093 30679 14151 30685
rect 16393 30685 16405 30688
rect 16439 30685 16451 30719
rect 16393 30679 16451 30685
rect 16660 30719 16718 30725
rect 16660 30685 16672 30719
rect 16706 30716 16718 30719
rect 18230 30716 18236 30728
rect 16706 30688 18236 30716
rect 16706 30685 16718 30688
rect 16660 30679 16718 30685
rect 18230 30676 18236 30688
rect 18288 30676 18294 30728
rect 19260 30725 19288 30756
rect 19245 30719 19303 30725
rect 19245 30685 19257 30719
rect 19291 30685 19303 30719
rect 22462 30716 22468 30728
rect 22520 30725 22526 30728
rect 22432 30688 22468 30716
rect 19245 30679 19303 30685
rect 22462 30676 22468 30688
rect 22520 30679 22532 30725
rect 22741 30719 22799 30725
rect 22741 30685 22753 30719
rect 22787 30716 22799 30719
rect 24026 30716 24032 30728
rect 22787 30688 24032 30716
rect 22787 30685 22799 30688
rect 22741 30679 22799 30685
rect 22520 30676 22526 30679
rect 24026 30676 24032 30688
rect 24084 30676 24090 30728
rect 68094 30716 68100 30728
rect 68055 30688 68100 30716
rect 68094 30676 68100 30688
rect 68152 30676 68158 30728
rect 7000 30651 7058 30657
rect 7000 30617 7012 30651
rect 7046 30648 7058 30651
rect 7098 30648 7104 30660
rect 7046 30620 7104 30648
rect 7046 30617 7058 30620
rect 7000 30611 7058 30617
rect 7098 30608 7104 30620
rect 7156 30608 7162 30660
rect 9214 30608 9220 30660
rect 9272 30648 9278 30660
rect 9493 30651 9551 30657
rect 9493 30648 9505 30651
rect 9272 30620 9505 30648
rect 9272 30608 9278 30620
rect 9493 30617 9505 30620
rect 9539 30617 9551 30651
rect 9493 30611 9551 30617
rect 9677 30651 9735 30657
rect 9677 30617 9689 30651
rect 9723 30648 9735 30651
rect 10962 30648 10968 30660
rect 9723 30620 10968 30648
rect 9723 30617 9735 30620
rect 9677 30611 9735 30617
rect 10962 30608 10968 30620
rect 11020 30608 11026 30660
rect 11692 30651 11750 30657
rect 11692 30617 11704 30651
rect 11738 30648 11750 30651
rect 13170 30648 13176 30660
rect 11738 30620 13176 30648
rect 11738 30617 11750 30620
rect 11692 30611 11750 30617
rect 13170 30608 13176 30620
rect 13228 30608 13234 30660
rect 14360 30651 14418 30657
rect 14360 30617 14372 30651
rect 14406 30648 14418 30651
rect 15102 30648 15108 30660
rect 14406 30620 15108 30648
rect 14406 30617 14418 30620
rect 14360 30611 14418 30617
rect 15102 30608 15108 30620
rect 15160 30608 15166 30660
rect 19426 30648 19432 30660
rect 19387 30620 19432 30648
rect 19426 30608 19432 30620
rect 19484 30608 19490 30660
rect 8110 30580 8116 30592
rect 8071 30552 8116 30580
rect 8110 30540 8116 30552
rect 8168 30540 8174 30592
rect 9766 30540 9772 30592
rect 9824 30580 9830 30592
rect 9861 30583 9919 30589
rect 9861 30580 9873 30583
rect 9824 30552 9873 30580
rect 9824 30540 9830 30552
rect 9861 30549 9873 30552
rect 9907 30549 9919 30583
rect 9861 30543 9919 30549
rect 12618 30540 12624 30592
rect 12676 30580 12682 30592
rect 12805 30583 12863 30589
rect 12805 30580 12817 30583
rect 12676 30552 12817 30580
rect 12676 30540 12682 30552
rect 12805 30549 12817 30552
rect 12851 30549 12863 30583
rect 12805 30543 12863 30549
rect 14090 30540 14096 30592
rect 14148 30580 14154 30592
rect 15746 30580 15752 30592
rect 14148 30552 15752 30580
rect 14148 30540 14154 30552
rect 15746 30540 15752 30552
rect 15804 30540 15810 30592
rect 17402 30540 17408 30592
rect 17460 30580 17466 30592
rect 17586 30580 17592 30592
rect 17460 30552 17592 30580
rect 17460 30540 17466 30552
rect 17586 30540 17592 30552
rect 17644 30580 17650 30592
rect 17773 30583 17831 30589
rect 17773 30580 17785 30583
rect 17644 30552 17785 30580
rect 17644 30540 17650 30552
rect 17773 30549 17785 30552
rect 17819 30549 17831 30583
rect 21358 30580 21364 30592
rect 21319 30552 21364 30580
rect 17773 30543 17831 30549
rect 21358 30540 21364 30552
rect 21416 30540 21422 30592
rect 1104 30490 68816 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 68816 30490
rect 1104 30416 68816 30438
rect 12894 30336 12900 30388
rect 12952 30376 12958 30388
rect 15930 30376 15936 30388
rect 12952 30348 15936 30376
rect 12952 30336 12958 30348
rect 1581 30311 1639 30317
rect 1581 30277 1593 30311
rect 1627 30308 1639 30311
rect 1670 30308 1676 30320
rect 1627 30280 1676 30308
rect 1627 30277 1639 30280
rect 1581 30271 1639 30277
rect 1670 30268 1676 30280
rect 1728 30308 1734 30320
rect 2593 30311 2651 30317
rect 1728 30280 2268 30308
rect 1728 30268 1734 30280
rect 1765 30243 1823 30249
rect 1765 30209 1777 30243
rect 1811 30209 1823 30243
rect 2240 30240 2268 30280
rect 2593 30277 2605 30311
rect 2639 30308 2651 30311
rect 4798 30308 4804 30320
rect 2639 30280 4384 30308
rect 2639 30277 2651 30280
rect 2593 30271 2651 30277
rect 2682 30240 2688 30252
rect 2240 30212 2688 30240
rect 1765 30203 1823 30209
rect 1780 30172 1808 30203
rect 2682 30200 2688 30212
rect 2740 30240 2746 30252
rect 2777 30243 2835 30249
rect 2777 30240 2789 30243
rect 2740 30212 2789 30240
rect 2740 30200 2746 30212
rect 2777 30209 2789 30212
rect 2823 30209 2835 30243
rect 2777 30203 2835 30209
rect 2866 30172 2872 30184
rect 1780 30144 2872 30172
rect 2866 30132 2872 30144
rect 2924 30132 2930 30184
rect 1949 30039 2007 30045
rect 1949 30005 1961 30039
rect 1995 30036 2007 30039
rect 2130 30036 2136 30048
rect 1995 30008 2136 30036
rect 1995 30005 2007 30008
rect 1949 29999 2007 30005
rect 2130 29996 2136 30008
rect 2188 29996 2194 30048
rect 2409 30039 2467 30045
rect 2409 30005 2421 30039
rect 2455 30036 2467 30039
rect 2498 30036 2504 30048
rect 2455 30008 2504 30036
rect 2455 30005 2467 30008
rect 2409 29999 2467 30005
rect 2498 29996 2504 30008
rect 2556 29996 2562 30048
rect 4356 30036 4384 30280
rect 4448 30280 4804 30308
rect 4448 30249 4476 30280
rect 4798 30268 4804 30280
rect 4856 30308 4862 30320
rect 6730 30308 6736 30320
rect 4856 30280 6736 30308
rect 4856 30268 4862 30280
rect 6730 30268 6736 30280
rect 6788 30268 6794 30320
rect 13170 30308 13176 30320
rect 13131 30280 13176 30308
rect 13170 30268 13176 30280
rect 13228 30268 13234 30320
rect 13648 30308 13676 30348
rect 15930 30336 15936 30348
rect 15988 30336 15994 30388
rect 18230 30336 18236 30388
rect 18288 30376 18294 30388
rect 23290 30376 23296 30388
rect 18288 30348 23296 30376
rect 18288 30336 18294 30348
rect 23290 30336 23296 30348
rect 23348 30376 23354 30388
rect 24489 30379 24547 30385
rect 24489 30376 24501 30379
rect 23348 30348 24501 30376
rect 23348 30336 23354 30348
rect 24489 30345 24501 30348
rect 24535 30345 24547 30379
rect 24489 30339 24547 30345
rect 13556 30280 13676 30308
rect 15565 30311 15623 30317
rect 13556 30252 13584 30280
rect 15565 30277 15577 30311
rect 15611 30308 15623 30311
rect 17126 30308 17132 30320
rect 15611 30280 17132 30308
rect 15611 30277 15623 30280
rect 15565 30271 15623 30277
rect 17126 30268 17132 30280
rect 17184 30268 17190 30320
rect 19978 30268 19984 30320
rect 20036 30308 20042 30320
rect 20634 30311 20692 30317
rect 20634 30308 20646 30311
rect 20036 30280 20646 30308
rect 20036 30268 20042 30280
rect 20634 30277 20646 30280
rect 20680 30277 20692 30311
rect 21818 30308 21824 30320
rect 21779 30280 21824 30308
rect 20634 30271 20692 30277
rect 21818 30268 21824 30280
rect 21876 30268 21882 30320
rect 24044 30280 25912 30308
rect 24044 30252 24072 30280
rect 4706 30249 4712 30252
rect 4433 30243 4491 30249
rect 4433 30209 4445 30243
rect 4479 30209 4491 30243
rect 4433 30203 4491 30209
rect 4700 30203 4712 30249
rect 4764 30240 4770 30252
rect 9306 30240 9312 30252
rect 4764 30212 4800 30240
rect 9267 30212 9312 30240
rect 4706 30200 4712 30203
rect 4764 30200 4770 30212
rect 9306 30200 9312 30212
rect 9364 30240 9370 30252
rect 9769 30243 9827 30249
rect 9769 30240 9781 30243
rect 9364 30212 9781 30240
rect 9364 30200 9370 30212
rect 9769 30209 9781 30212
rect 9815 30209 9827 30243
rect 13446 30240 13452 30252
rect 13407 30212 13452 30240
rect 9769 30203 9827 30209
rect 13446 30200 13452 30212
rect 13504 30200 13510 30252
rect 13538 30246 13596 30252
rect 13538 30212 13550 30246
rect 13584 30212 13596 30246
rect 13538 30206 13596 30212
rect 13630 30200 13636 30252
rect 13688 30249 13694 30252
rect 13688 30240 13696 30249
rect 13817 30243 13875 30249
rect 13688 30212 13733 30240
rect 13688 30203 13696 30212
rect 13817 30209 13829 30243
rect 13863 30240 13875 30243
rect 14090 30240 14096 30252
rect 13863 30212 14096 30240
rect 13863 30209 13875 30212
rect 13817 30203 13875 30209
rect 13688 30200 13694 30203
rect 14090 30200 14096 30212
rect 14148 30200 14154 30252
rect 15286 30200 15292 30252
rect 15344 30240 15350 30252
rect 15381 30243 15439 30249
rect 15381 30240 15393 30243
rect 15344 30212 15393 30240
rect 15344 30200 15350 30212
rect 15381 30209 15393 30212
rect 15427 30209 15439 30243
rect 15654 30240 15660 30252
rect 15615 30212 15660 30240
rect 15381 30203 15439 30209
rect 15654 30200 15660 30212
rect 15712 30200 15718 30252
rect 15749 30243 15807 30249
rect 15749 30209 15761 30243
rect 15795 30240 15807 30243
rect 22005 30243 22063 30249
rect 15795 30212 15829 30240
rect 15795 30209 15807 30212
rect 15749 30203 15807 30209
rect 22005 30209 22017 30243
rect 22051 30209 22063 30243
rect 22005 30203 22063 30209
rect 14921 30175 14979 30181
rect 14921 30141 14933 30175
rect 14967 30172 14979 30175
rect 15764 30172 15792 30203
rect 16574 30172 16580 30184
rect 14967 30144 16580 30172
rect 14967 30141 14979 30144
rect 14921 30135 14979 30141
rect 16574 30132 16580 30144
rect 16632 30132 16638 30184
rect 20901 30175 20959 30181
rect 20901 30141 20913 30175
rect 20947 30172 20959 30175
rect 21450 30172 21456 30184
rect 20947 30144 21456 30172
rect 20947 30141 20959 30144
rect 20901 30135 20959 30141
rect 21450 30132 21456 30144
rect 21508 30132 21514 30184
rect 22020 30116 22048 30203
rect 22554 30200 22560 30252
rect 22612 30240 22618 30252
rect 23762 30243 23820 30249
rect 23762 30240 23774 30243
rect 22612 30212 23774 30240
rect 22612 30200 22618 30212
rect 23762 30209 23774 30212
rect 23808 30209 23820 30243
rect 24026 30240 24032 30252
rect 23987 30212 24032 30240
rect 23762 30203 23820 30209
rect 24026 30200 24032 30212
rect 24084 30200 24090 30252
rect 25590 30200 25596 30252
rect 25648 30249 25654 30252
rect 25884 30249 25912 30280
rect 25648 30240 25660 30249
rect 25869 30243 25927 30249
rect 25648 30212 25693 30240
rect 25648 30203 25660 30212
rect 25869 30209 25881 30243
rect 25915 30209 25927 30243
rect 25869 30203 25927 30209
rect 25648 30200 25654 30203
rect 5810 30104 5816 30116
rect 5771 30076 5816 30104
rect 5810 30064 5816 30076
rect 5868 30064 5874 30116
rect 6730 30064 6736 30116
rect 6788 30104 6794 30116
rect 7742 30104 7748 30116
rect 6788 30076 7748 30104
rect 6788 30064 6794 30076
rect 7742 30064 7748 30076
rect 7800 30104 7806 30116
rect 8021 30107 8079 30113
rect 8021 30104 8033 30107
rect 7800 30076 8033 30104
rect 7800 30064 7806 30076
rect 8021 30073 8033 30076
rect 8067 30104 8079 30107
rect 11054 30104 11060 30116
rect 8067 30076 11060 30104
rect 8067 30073 8079 30076
rect 8021 30067 8079 30073
rect 11054 30064 11060 30076
rect 11112 30064 11118 30116
rect 13446 30064 13452 30116
rect 13504 30104 13510 30116
rect 14369 30107 14427 30113
rect 14369 30104 14381 30107
rect 13504 30076 14381 30104
rect 13504 30064 13510 30076
rect 14369 30073 14381 30076
rect 14415 30104 14427 30107
rect 14415 30076 20024 30104
rect 14415 30073 14427 30076
rect 14369 30067 14427 30073
rect 5828 30036 5856 30064
rect 4356 30008 5856 30036
rect 15933 30039 15991 30045
rect 15933 30005 15945 30039
rect 15979 30036 15991 30039
rect 18046 30036 18052 30048
rect 15979 30008 18052 30036
rect 15979 30005 15991 30008
rect 15933 29999 15991 30005
rect 18046 29996 18052 30008
rect 18104 29996 18110 30048
rect 19518 30036 19524 30048
rect 19479 30008 19524 30036
rect 19518 29996 19524 30008
rect 19576 29996 19582 30048
rect 19996 30036 20024 30076
rect 22002 30064 22008 30116
rect 22060 30104 22066 30116
rect 22649 30107 22707 30113
rect 22649 30104 22661 30107
rect 22060 30076 22661 30104
rect 22060 30064 22066 30076
rect 22649 30073 22661 30076
rect 22695 30073 22707 30107
rect 22649 30067 22707 30073
rect 20990 30036 20996 30048
rect 19996 30008 20996 30036
rect 20990 29996 20996 30008
rect 21048 29996 21054 30048
rect 22094 29996 22100 30048
rect 22152 30036 22158 30048
rect 22189 30039 22247 30045
rect 22189 30036 22201 30039
rect 22152 30008 22201 30036
rect 22152 29996 22158 30008
rect 22189 30005 22201 30008
rect 22235 30005 22247 30039
rect 22189 29999 22247 30005
rect 1104 29946 68816 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 65654 29946
rect 65706 29894 65718 29946
rect 65770 29894 65782 29946
rect 65834 29894 65846 29946
rect 65898 29894 65910 29946
rect 65962 29894 68816 29946
rect 1104 29872 68816 29894
rect 2593 29835 2651 29841
rect 2593 29801 2605 29835
rect 2639 29832 2651 29835
rect 3418 29832 3424 29844
rect 2639 29804 3424 29832
rect 2639 29801 2651 29804
rect 2593 29795 2651 29801
rect 3418 29792 3424 29804
rect 3476 29792 3482 29844
rect 10962 29832 10968 29844
rect 10875 29804 10968 29832
rect 10962 29792 10968 29804
rect 11020 29832 11026 29844
rect 19518 29832 19524 29844
rect 11020 29804 17540 29832
rect 11020 29792 11026 29804
rect 1397 29767 1455 29773
rect 1397 29733 1409 29767
rect 1443 29764 1455 29767
rect 2774 29764 2780 29776
rect 1443 29736 2780 29764
rect 1443 29733 1455 29736
rect 1397 29727 1455 29733
rect 1946 29628 1952 29640
rect 1907 29600 1952 29628
rect 1946 29588 1952 29600
rect 2004 29588 2010 29640
rect 2130 29628 2136 29640
rect 2091 29600 2136 29628
rect 2130 29588 2136 29600
rect 2188 29588 2194 29640
rect 2332 29637 2360 29736
rect 2774 29724 2780 29736
rect 2832 29764 2838 29776
rect 9398 29764 9404 29776
rect 2832 29736 9404 29764
rect 2832 29724 2838 29736
rect 9398 29724 9404 29736
rect 9456 29724 9462 29776
rect 12069 29767 12127 29773
rect 12069 29733 12081 29767
rect 12115 29764 12127 29767
rect 13262 29764 13268 29776
rect 12115 29736 13268 29764
rect 12115 29733 12127 29736
rect 12069 29727 12127 29733
rect 13262 29724 13268 29736
rect 13320 29724 13326 29776
rect 12894 29656 12900 29708
rect 12952 29696 12958 29708
rect 12952 29668 13308 29696
rect 12952 29656 12958 29668
rect 2225 29631 2283 29637
rect 2225 29597 2237 29631
rect 2271 29597 2283 29631
rect 2225 29591 2283 29597
rect 2317 29631 2375 29637
rect 2317 29597 2329 29631
rect 2363 29597 2375 29631
rect 7282 29628 7288 29640
rect 7243 29600 7288 29628
rect 2317 29591 2375 29597
rect 2240 29560 2268 29591
rect 7282 29588 7288 29600
rect 7340 29588 7346 29640
rect 7469 29631 7527 29637
rect 7469 29597 7481 29631
rect 7515 29628 7527 29631
rect 9585 29631 9643 29637
rect 7515 29600 8340 29628
rect 7515 29597 7527 29600
rect 7469 29591 7527 29597
rect 2406 29560 2412 29572
rect 2240 29532 2412 29560
rect 2406 29520 2412 29532
rect 2464 29520 2470 29572
rect 2682 29520 2688 29572
rect 2740 29560 2746 29572
rect 3789 29563 3847 29569
rect 3789 29560 3801 29563
rect 2740 29532 3801 29560
rect 2740 29520 2746 29532
rect 3789 29529 3801 29532
rect 3835 29529 3847 29563
rect 3789 29523 3847 29529
rect 3973 29563 4031 29569
rect 3973 29529 3985 29563
rect 4019 29560 4031 29563
rect 5442 29560 5448 29572
rect 4019 29532 5448 29560
rect 4019 29529 4031 29532
rect 3973 29523 4031 29529
rect 5442 29520 5448 29532
rect 5500 29520 5506 29572
rect 6181 29563 6239 29569
rect 6181 29529 6193 29563
rect 6227 29560 6239 29563
rect 7190 29560 7196 29572
rect 6227 29532 7196 29560
rect 6227 29529 6239 29532
rect 6181 29523 6239 29529
rect 7190 29520 7196 29532
rect 7248 29520 7254 29572
rect 8312 29569 8340 29600
rect 9585 29597 9597 29631
rect 9631 29628 9643 29631
rect 11054 29628 11060 29640
rect 9631 29600 11060 29628
rect 9631 29597 9643 29600
rect 9585 29591 9643 29597
rect 11054 29588 11060 29600
rect 11112 29588 11118 29640
rect 12253 29631 12311 29637
rect 12253 29597 12265 29631
rect 12299 29628 12311 29631
rect 12986 29628 12992 29640
rect 12299 29600 12992 29628
rect 12299 29597 12311 29600
rect 12253 29591 12311 29597
rect 12986 29588 12992 29600
rect 13044 29588 13050 29640
rect 13078 29588 13084 29640
rect 13136 29625 13142 29640
rect 13280 29637 13308 29668
rect 13446 29656 13452 29708
rect 13504 29696 13510 29708
rect 14185 29699 14243 29705
rect 14185 29696 14197 29699
rect 13504 29668 14197 29696
rect 13504 29656 13510 29668
rect 14185 29665 14197 29668
rect 14231 29696 14243 29699
rect 17034 29696 17040 29708
rect 14231 29668 17040 29696
rect 14231 29665 14243 29668
rect 14185 29659 14243 29665
rect 17034 29656 17040 29668
rect 17092 29656 17098 29708
rect 13173 29631 13231 29637
rect 13173 29625 13185 29631
rect 13136 29597 13185 29625
rect 13219 29597 13231 29631
rect 13136 29588 13142 29597
rect 13173 29591 13231 29597
rect 13262 29631 13320 29637
rect 13262 29597 13274 29631
rect 13308 29597 13320 29631
rect 13262 29591 13320 29597
rect 13354 29588 13360 29640
rect 13412 29628 13418 29640
rect 13541 29631 13599 29637
rect 13412 29600 13457 29628
rect 13412 29588 13418 29600
rect 13541 29597 13553 29631
rect 13587 29628 13599 29631
rect 14090 29628 14096 29640
rect 13587 29600 14096 29628
rect 13587 29597 13599 29600
rect 13541 29591 13599 29597
rect 14090 29588 14096 29600
rect 14148 29628 14154 29640
rect 14734 29628 14740 29640
rect 14148 29600 14740 29628
rect 14148 29588 14154 29600
rect 14734 29588 14740 29600
rect 14792 29588 14798 29640
rect 17221 29631 17279 29637
rect 17221 29628 17233 29631
rect 16592 29600 17233 29628
rect 8113 29563 8171 29569
rect 8113 29529 8125 29563
rect 8159 29529 8171 29563
rect 8113 29523 8171 29529
rect 8297 29563 8355 29569
rect 8297 29529 8309 29563
rect 8343 29560 8355 29563
rect 9214 29560 9220 29572
rect 8343 29532 9220 29560
rect 8343 29529 8355 29532
rect 8297 29523 8355 29529
rect 4154 29492 4160 29504
rect 4115 29464 4160 29492
rect 4154 29452 4160 29464
rect 4212 29452 4218 29504
rect 6638 29452 6644 29504
rect 6696 29492 6702 29504
rect 7101 29495 7159 29501
rect 7101 29492 7113 29495
rect 6696 29464 7113 29492
rect 6696 29452 6702 29464
rect 7101 29461 7113 29464
rect 7147 29461 7159 29495
rect 7101 29455 7159 29461
rect 7650 29452 7656 29504
rect 7708 29492 7714 29504
rect 7929 29495 7987 29501
rect 7929 29492 7941 29495
rect 7708 29464 7941 29492
rect 7708 29452 7714 29464
rect 7929 29461 7941 29464
rect 7975 29461 7987 29495
rect 8128 29492 8156 29523
rect 9214 29520 9220 29532
rect 9272 29520 9278 29572
rect 9852 29563 9910 29569
rect 9852 29529 9864 29563
rect 9898 29560 9910 29563
rect 10226 29560 10232 29572
rect 9898 29532 10232 29560
rect 9898 29529 9910 29532
rect 9852 29523 9910 29529
rect 10226 29520 10232 29532
rect 10284 29520 10290 29572
rect 12434 29560 12440 29572
rect 12395 29532 12440 29560
rect 12434 29520 12440 29532
rect 12492 29520 12498 29572
rect 16592 29504 16620 29600
rect 17221 29597 17233 29600
rect 17267 29597 17279 29631
rect 17221 29591 17279 29597
rect 17310 29588 17316 29640
rect 17368 29628 17374 29640
rect 17368 29600 17413 29628
rect 17368 29588 17374 29600
rect 17126 29520 17132 29572
rect 17184 29560 17190 29572
rect 17405 29563 17463 29569
rect 17405 29560 17417 29563
rect 17184 29532 17417 29560
rect 17184 29520 17190 29532
rect 17405 29529 17417 29532
rect 17451 29529 17463 29563
rect 17512 29560 17540 29804
rect 17604 29804 19524 29832
rect 17604 29637 17632 29804
rect 19518 29792 19524 29804
rect 19576 29792 19582 29844
rect 22554 29832 22560 29844
rect 22515 29804 22560 29832
rect 22554 29792 22560 29804
rect 22612 29792 22618 29844
rect 22094 29764 22100 29776
rect 22020 29736 22100 29764
rect 21358 29696 21364 29708
rect 18340 29668 19104 29696
rect 17589 29631 17647 29637
rect 17589 29597 17601 29631
rect 17635 29597 17647 29631
rect 18046 29628 18052 29640
rect 18007 29600 18052 29628
rect 17589 29591 17647 29597
rect 18046 29588 18052 29600
rect 18104 29588 18110 29640
rect 18230 29637 18236 29640
rect 18197 29631 18236 29637
rect 18197 29597 18209 29631
rect 18197 29591 18236 29597
rect 18230 29588 18236 29591
rect 18288 29588 18294 29640
rect 18340 29637 18368 29668
rect 18325 29631 18383 29637
rect 18325 29597 18337 29631
rect 18371 29597 18383 29631
rect 18325 29591 18383 29597
rect 18506 29588 18512 29640
rect 18564 29637 18570 29640
rect 18564 29628 18572 29637
rect 18564 29600 18609 29628
rect 18564 29591 18572 29600
rect 18564 29588 18570 29591
rect 19076 29572 19104 29668
rect 19628 29668 21364 29696
rect 19242 29628 19248 29640
rect 19203 29600 19248 29628
rect 19242 29588 19248 29600
rect 19300 29588 19306 29640
rect 19393 29631 19451 29637
rect 19393 29597 19405 29631
rect 19439 29628 19451 29631
rect 19628 29628 19656 29668
rect 21358 29656 21364 29668
rect 21416 29656 21422 29708
rect 19439 29600 19656 29628
rect 19710 29631 19768 29637
rect 19439 29597 19451 29600
rect 19393 29591 19451 29597
rect 19710 29597 19722 29631
rect 19756 29628 19768 29631
rect 21913 29631 21971 29637
rect 19756 29600 19840 29628
rect 19756 29597 19768 29600
rect 19710 29591 19768 29597
rect 18417 29563 18475 29569
rect 18417 29560 18429 29563
rect 17512 29532 18429 29560
rect 17405 29523 17463 29529
rect 18417 29529 18429 29532
rect 18463 29529 18475 29563
rect 18417 29523 18475 29529
rect 19058 29520 19064 29572
rect 19116 29560 19122 29572
rect 19521 29563 19579 29569
rect 19521 29560 19533 29563
rect 19116 29532 19533 29560
rect 19116 29520 19122 29532
rect 19521 29529 19533 29532
rect 19567 29529 19579 29563
rect 19521 29523 19579 29529
rect 19610 29520 19616 29572
rect 19668 29560 19674 29572
rect 19812 29560 19840 29600
rect 21913 29597 21925 29631
rect 21959 29597 21971 29631
rect 22020 29628 22048 29736
rect 22094 29724 22100 29736
rect 22152 29724 22158 29776
rect 22186 29724 22192 29776
rect 22244 29724 22250 29776
rect 22207 29696 22235 29724
rect 22204 29668 22235 29696
rect 22076 29631 22134 29637
rect 22204 29634 22232 29668
rect 22076 29628 22088 29631
rect 22020 29600 22088 29628
rect 21913 29591 21971 29597
rect 22076 29597 22088 29600
rect 22122 29597 22134 29631
rect 22076 29591 22134 29597
rect 22176 29628 22234 29634
rect 22176 29594 22188 29628
rect 22222 29594 22234 29628
rect 20349 29563 20407 29569
rect 20349 29560 20361 29563
rect 19668 29532 19713 29560
rect 19812 29532 20361 29560
rect 19668 29520 19674 29532
rect 9122 29492 9128 29504
rect 8128 29464 9128 29492
rect 7929 29455 7987 29461
rect 9122 29452 9128 29464
rect 9180 29452 9186 29504
rect 12802 29452 12808 29504
rect 12860 29492 12866 29504
rect 12897 29495 12955 29501
rect 12897 29492 12909 29495
rect 12860 29464 12909 29492
rect 12860 29452 12866 29464
rect 12897 29461 12909 29464
rect 12943 29461 12955 29495
rect 16574 29492 16580 29504
rect 16535 29464 16580 29492
rect 12897 29455 12955 29461
rect 16574 29452 16580 29464
rect 16632 29452 16638 29504
rect 17037 29495 17095 29501
rect 17037 29461 17049 29495
rect 17083 29492 17095 29495
rect 18598 29492 18604 29504
rect 17083 29464 18604 29492
rect 17083 29461 17095 29464
rect 17037 29455 17095 29461
rect 18598 29452 18604 29464
rect 18656 29452 18662 29504
rect 18693 29495 18751 29501
rect 18693 29461 18705 29495
rect 18739 29492 18751 29495
rect 19150 29492 19156 29504
rect 18739 29464 19156 29492
rect 18739 29461 18751 29464
rect 18693 29455 18751 29461
rect 19150 29452 19156 29464
rect 19208 29452 19214 29504
rect 19426 29452 19432 29504
rect 19484 29492 19490 29504
rect 19812 29492 19840 29532
rect 20349 29529 20361 29532
rect 20395 29529 20407 29563
rect 20349 29523 20407 29529
rect 19484 29464 19840 29492
rect 19889 29495 19947 29501
rect 19484 29452 19490 29464
rect 19889 29461 19901 29495
rect 19935 29492 19947 29495
rect 20254 29492 20260 29504
rect 19935 29464 20260 29492
rect 19935 29461 19947 29464
rect 19889 29455 19947 29461
rect 20254 29452 20260 29464
rect 20312 29452 20318 29504
rect 21928 29492 21956 29591
rect 22176 29588 22234 29594
rect 22281 29631 22339 29637
rect 22281 29597 22293 29631
rect 22327 29628 22339 29631
rect 22370 29628 22376 29640
rect 22327 29600 22376 29628
rect 22327 29597 22339 29600
rect 22281 29591 22339 29597
rect 22370 29588 22376 29600
rect 22428 29588 22434 29640
rect 26970 29628 26976 29640
rect 26931 29600 26976 29628
rect 26970 29588 26976 29600
rect 27028 29588 27034 29640
rect 68094 29628 68100 29640
rect 68055 29600 68100 29628
rect 68094 29588 68100 29600
rect 68152 29588 68158 29640
rect 26234 29520 26240 29572
rect 26292 29560 26298 29572
rect 26706 29563 26764 29569
rect 26706 29560 26718 29563
rect 26292 29532 26718 29560
rect 26292 29520 26298 29532
rect 26706 29529 26718 29532
rect 26752 29529 26764 29563
rect 26706 29523 26764 29529
rect 23474 29492 23480 29504
rect 21928 29464 23480 29492
rect 23474 29452 23480 29464
rect 23532 29492 23538 29504
rect 25222 29492 25228 29504
rect 23532 29464 25228 29492
rect 23532 29452 23538 29464
rect 25222 29452 25228 29464
rect 25280 29452 25286 29504
rect 25498 29452 25504 29504
rect 25556 29492 25562 29504
rect 25593 29495 25651 29501
rect 25593 29492 25605 29495
rect 25556 29464 25605 29492
rect 25556 29452 25562 29464
rect 25593 29461 25605 29464
rect 25639 29461 25651 29495
rect 25593 29455 25651 29461
rect 1104 29402 68816 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 68816 29402
rect 1104 29328 68816 29350
rect 2406 29248 2412 29300
rect 2464 29248 2470 29300
rect 3053 29291 3111 29297
rect 3053 29257 3065 29291
rect 3099 29288 3111 29291
rect 4706 29288 4712 29300
rect 3099 29260 4712 29288
rect 3099 29257 3111 29260
rect 3053 29251 3111 29257
rect 4706 29248 4712 29260
rect 4764 29248 4770 29300
rect 7098 29288 7104 29300
rect 7059 29260 7104 29288
rect 7098 29248 7104 29260
rect 7156 29248 7162 29300
rect 9950 29288 9956 29300
rect 9876 29260 9956 29288
rect 2424 29220 2452 29248
rect 4798 29220 4804 29232
rect 2424 29192 2728 29220
rect 1946 29112 1952 29164
rect 2004 29152 2010 29164
rect 2409 29155 2467 29161
rect 2409 29152 2421 29155
rect 2004 29124 2421 29152
rect 2004 29112 2010 29124
rect 2409 29121 2421 29124
rect 2455 29121 2467 29155
rect 2409 29115 2467 29121
rect 2424 29084 2452 29115
rect 2498 29112 2504 29164
rect 2556 29152 2562 29164
rect 2700 29161 2728 29192
rect 4080 29192 4804 29220
rect 4080 29161 4108 29192
rect 4798 29180 4804 29192
rect 4856 29180 4862 29232
rect 7190 29220 7196 29232
rect 6472 29192 7196 29220
rect 2593 29155 2651 29161
rect 2593 29152 2605 29155
rect 2556 29124 2605 29152
rect 2556 29112 2562 29124
rect 2593 29121 2605 29124
rect 2639 29121 2651 29155
rect 2593 29115 2651 29121
rect 2685 29155 2743 29161
rect 2685 29121 2697 29155
rect 2731 29121 2743 29155
rect 2685 29115 2743 29121
rect 2777 29155 2835 29161
rect 2777 29121 2789 29155
rect 2823 29152 2835 29155
rect 4065 29155 4123 29161
rect 2823 29124 3648 29152
rect 2823 29121 2835 29124
rect 2777 29115 2835 29121
rect 2424 29056 2636 29084
rect 2608 29028 2636 29056
rect 2590 28976 2596 29028
rect 2648 28976 2654 29028
rect 2682 28976 2688 29028
rect 2740 29016 2746 29028
rect 2774 29016 2780 29028
rect 2740 28988 2780 29016
rect 2740 28976 2746 28988
rect 2774 28976 2780 28988
rect 2832 28976 2838 29028
rect 3620 29025 3648 29124
rect 4065 29121 4077 29155
rect 4111 29121 4123 29155
rect 4065 29115 4123 29121
rect 4332 29155 4390 29161
rect 4332 29121 4344 29155
rect 4378 29152 4390 29155
rect 4614 29152 4620 29164
rect 4378 29124 4620 29152
rect 4378 29121 4390 29124
rect 4332 29115 4390 29121
rect 4614 29112 4620 29124
rect 4672 29112 4678 29164
rect 6472 29161 6500 29192
rect 7190 29180 7196 29192
rect 7248 29180 7254 29232
rect 6457 29155 6515 29161
rect 6457 29121 6469 29155
rect 6503 29121 6515 29155
rect 6638 29152 6644 29164
rect 6599 29124 6644 29152
rect 6457 29115 6515 29121
rect 6638 29112 6644 29124
rect 6696 29112 6702 29164
rect 6733 29155 6791 29161
rect 6733 29121 6745 29155
rect 6779 29121 6791 29155
rect 6733 29115 6791 29121
rect 6748 29084 6776 29115
rect 6822 29112 6828 29164
rect 6880 29152 6886 29164
rect 7742 29152 7748 29164
rect 6880 29124 6925 29152
rect 7703 29124 7748 29152
rect 6880 29112 6886 29124
rect 7742 29112 7748 29124
rect 7800 29112 7806 29164
rect 8018 29161 8024 29164
rect 8012 29115 8024 29161
rect 8076 29152 8082 29164
rect 8076 29124 8112 29152
rect 8018 29112 8024 29115
rect 8076 29112 8082 29124
rect 9490 29112 9496 29164
rect 9548 29152 9554 29164
rect 9585 29155 9643 29161
rect 9585 29152 9597 29155
rect 9548 29124 9597 29152
rect 9548 29112 9554 29124
rect 9585 29121 9597 29124
rect 9631 29121 9643 29155
rect 9766 29152 9772 29164
rect 9727 29124 9772 29152
rect 9585 29115 9643 29121
rect 9766 29112 9772 29124
rect 9824 29112 9830 29164
rect 9876 29161 9904 29260
rect 9950 29248 9956 29260
rect 10008 29248 10014 29300
rect 10226 29288 10232 29300
rect 10187 29260 10232 29288
rect 10226 29248 10232 29260
rect 10284 29248 10290 29300
rect 11517 29291 11575 29297
rect 11517 29257 11529 29291
rect 11563 29288 11575 29291
rect 12986 29288 12992 29300
rect 11563 29260 12992 29288
rect 11563 29257 11575 29260
rect 11517 29251 11575 29257
rect 12986 29248 12992 29260
rect 13044 29248 13050 29300
rect 15194 29248 15200 29300
rect 15252 29288 15258 29300
rect 15381 29291 15439 29297
rect 15381 29288 15393 29291
rect 15252 29260 15393 29288
rect 15252 29248 15258 29260
rect 15381 29257 15393 29260
rect 15427 29257 15439 29291
rect 15930 29288 15936 29300
rect 15891 29260 15936 29288
rect 15381 29251 15439 29257
rect 15930 29248 15936 29260
rect 15988 29248 15994 29300
rect 16853 29291 16911 29297
rect 16853 29257 16865 29291
rect 16899 29288 16911 29291
rect 19242 29288 19248 29300
rect 16899 29260 19248 29288
rect 16899 29257 16911 29260
rect 16853 29251 16911 29257
rect 19242 29248 19248 29260
rect 19300 29248 19306 29300
rect 12526 29220 12532 29232
rect 10152 29192 12532 29220
rect 9861 29155 9919 29161
rect 9861 29121 9873 29155
rect 9907 29121 9919 29155
rect 9861 29115 9919 29121
rect 9953 29155 10011 29161
rect 9953 29121 9965 29155
rect 9999 29152 10011 29155
rect 10042 29152 10048 29164
rect 9999 29124 10048 29152
rect 9999 29121 10011 29124
rect 9953 29115 10011 29121
rect 10042 29112 10048 29124
rect 10100 29112 10106 29164
rect 7374 29084 7380 29096
rect 5276 29056 5672 29084
rect 6748 29056 7380 29084
rect 3605 29019 3663 29025
rect 3605 28985 3617 29019
rect 3651 29016 3663 29019
rect 5276 29016 5304 29056
rect 5442 29016 5448 29028
rect 3651 28988 4108 29016
rect 3651 28985 3663 28988
rect 3605 28979 3663 28985
rect 4080 28948 4108 28988
rect 5000 28988 5304 29016
rect 5403 28988 5448 29016
rect 5000 28948 5028 28988
rect 5442 28976 5448 28988
rect 5500 28976 5506 29028
rect 5644 29016 5672 29056
rect 7374 29044 7380 29056
rect 7432 29044 7438 29096
rect 9306 29044 9312 29096
rect 9364 29084 9370 29096
rect 10152 29084 10180 29192
rect 12526 29180 12532 29192
rect 12584 29220 12590 29232
rect 14277 29223 14335 29229
rect 14277 29220 14289 29223
rect 12584 29192 14289 29220
rect 12584 29180 12590 29192
rect 14277 29189 14289 29192
rect 14323 29220 14335 29223
rect 14458 29220 14464 29232
rect 14323 29192 14464 29220
rect 14323 29189 14335 29192
rect 14277 29183 14335 29189
rect 14458 29180 14464 29192
rect 14516 29180 14522 29232
rect 17218 29220 17224 29232
rect 17131 29192 17224 29220
rect 17218 29180 17224 29192
rect 17276 29220 17282 29232
rect 17494 29220 17500 29232
rect 17276 29192 17500 29220
rect 17276 29180 17282 29192
rect 17494 29180 17500 29192
rect 17552 29180 17558 29232
rect 22002 29220 22008 29232
rect 19168 29192 22008 29220
rect 12641 29155 12699 29161
rect 12641 29121 12653 29155
rect 12687 29152 12699 29155
rect 12802 29152 12808 29164
rect 12687 29124 12808 29152
rect 12687 29121 12699 29124
rect 12641 29115 12699 29121
rect 12802 29112 12808 29124
rect 12860 29112 12866 29164
rect 14642 29112 14648 29164
rect 14700 29152 14706 29164
rect 15197 29155 15255 29161
rect 15197 29152 15209 29155
rect 14700 29124 15209 29152
rect 14700 29112 14706 29124
rect 15197 29121 15209 29124
rect 15243 29121 15255 29155
rect 15197 29115 15255 29121
rect 16025 29155 16083 29161
rect 16025 29121 16037 29155
rect 16071 29152 16083 29155
rect 16298 29152 16304 29164
rect 16071 29124 16304 29152
rect 16071 29121 16083 29124
rect 16025 29115 16083 29121
rect 16298 29112 16304 29124
rect 16356 29112 16362 29164
rect 16574 29112 16580 29164
rect 16632 29152 16638 29164
rect 17037 29155 17095 29161
rect 17037 29152 17049 29155
rect 16632 29124 17049 29152
rect 16632 29112 16638 29124
rect 17037 29121 17049 29124
rect 17083 29121 17095 29155
rect 17037 29115 17095 29121
rect 17126 29112 17132 29164
rect 17184 29152 17190 29164
rect 17402 29152 17408 29164
rect 17184 29124 17229 29152
rect 17363 29124 17408 29152
rect 17184 29112 17190 29124
rect 17402 29112 17408 29124
rect 17460 29112 17466 29164
rect 18598 29112 18604 29164
rect 18656 29152 18662 29164
rect 19168 29161 19196 29192
rect 22002 29180 22008 29192
rect 22060 29180 22066 29232
rect 24026 29180 24032 29232
rect 24084 29220 24090 29232
rect 26970 29220 26976 29232
rect 24084 29192 26976 29220
rect 24084 29180 24090 29192
rect 18969 29155 19027 29161
rect 18969 29152 18981 29155
rect 18656 29124 18981 29152
rect 18656 29112 18662 29124
rect 18969 29121 18981 29124
rect 19015 29121 19027 29155
rect 18969 29115 19027 29121
rect 19117 29155 19196 29161
rect 19117 29121 19129 29155
rect 19163 29124 19196 29155
rect 19245 29155 19303 29161
rect 19163 29121 19175 29124
rect 19117 29115 19175 29121
rect 19245 29121 19257 29155
rect 19291 29121 19303 29155
rect 19245 29115 19303 29121
rect 19337 29155 19395 29161
rect 19337 29121 19349 29155
rect 19383 29121 19395 29155
rect 19337 29115 19395 29121
rect 9364 29056 10180 29084
rect 12897 29087 12955 29093
rect 9364 29044 9370 29056
rect 12897 29053 12909 29087
rect 12943 29084 12955 29087
rect 13814 29084 13820 29096
rect 12943 29056 13820 29084
rect 12943 29053 12955 29056
rect 12897 29047 12955 29053
rect 13814 29044 13820 29056
rect 13872 29044 13878 29096
rect 18874 29044 18880 29096
rect 18932 29084 18938 29096
rect 19260 29084 19288 29115
rect 18932 29056 19288 29084
rect 18932 29044 18938 29056
rect 7006 29016 7012 29028
rect 5644 28988 7012 29016
rect 7006 28976 7012 28988
rect 7064 28976 7070 29028
rect 9122 29016 9128 29028
rect 9035 28988 9128 29016
rect 9122 28976 9128 28988
rect 9180 29016 9186 29028
rect 19352 29016 19380 29115
rect 19426 29112 19432 29164
rect 19484 29161 19490 29164
rect 19484 29152 19492 29161
rect 19484 29124 19577 29152
rect 19484 29115 19492 29124
rect 19484 29112 19490 29115
rect 23842 29112 23848 29164
rect 23900 29152 23906 29164
rect 25148 29161 25176 29192
rect 26970 29180 26976 29192
rect 27028 29220 27034 29232
rect 27341 29223 27399 29229
rect 27341 29220 27353 29223
rect 27028 29192 27353 29220
rect 27028 29180 27034 29192
rect 27341 29189 27353 29192
rect 27387 29189 27399 29223
rect 27341 29183 27399 29189
rect 24866 29155 24924 29161
rect 24866 29152 24878 29155
rect 23900 29124 24878 29152
rect 23900 29112 23906 29124
rect 24866 29121 24878 29124
rect 24912 29121 24924 29155
rect 24866 29115 24924 29121
rect 25133 29155 25191 29161
rect 25133 29121 25145 29155
rect 25179 29121 25191 29155
rect 29086 29152 29092 29164
rect 28999 29124 29092 29152
rect 25133 29115 25191 29121
rect 29086 29112 29092 29124
rect 29144 29152 29150 29164
rect 29549 29155 29607 29161
rect 29549 29152 29561 29155
rect 29144 29124 29561 29152
rect 29144 29112 29150 29124
rect 29549 29121 29561 29124
rect 29595 29121 29607 29155
rect 29549 29115 29607 29121
rect 9180 28988 12020 29016
rect 9180 28976 9186 28988
rect 4080 28920 5028 28948
rect 11992 28948 12020 28988
rect 12912 28988 19380 29016
rect 12912 28948 12940 28988
rect 17954 28948 17960 28960
rect 11992 28920 12940 28948
rect 17915 28920 17960 28948
rect 17954 28908 17960 28920
rect 18012 28948 18018 28960
rect 18417 28951 18475 28957
rect 18417 28948 18429 28951
rect 18012 28920 18429 28948
rect 18012 28908 18018 28920
rect 18417 28917 18429 28920
rect 18463 28948 18475 28951
rect 18506 28948 18512 28960
rect 18463 28920 18512 28948
rect 18463 28917 18475 28920
rect 18417 28911 18475 28917
rect 18506 28908 18512 28920
rect 18564 28948 18570 28960
rect 19444 28948 19472 29112
rect 19613 29019 19671 29025
rect 19613 28985 19625 29019
rect 19659 29016 19671 29019
rect 20162 29016 20168 29028
rect 19659 28988 20168 29016
rect 19659 28985 19671 28988
rect 19613 28979 19671 28985
rect 20162 28976 20168 28988
rect 20220 28976 20226 29028
rect 23750 29016 23756 29028
rect 23711 28988 23756 29016
rect 23750 28976 23756 28988
rect 23808 28976 23814 29028
rect 18564 28920 19472 28948
rect 18564 28908 18570 28920
rect 1104 28858 68816 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 65654 28858
rect 65706 28806 65718 28858
rect 65770 28806 65782 28858
rect 65834 28806 65846 28858
rect 65898 28806 65910 28858
rect 65962 28806 68816 28858
rect 1104 28784 68816 28806
rect 4433 28747 4491 28753
rect 4433 28713 4445 28747
rect 4479 28744 4491 28747
rect 4614 28744 4620 28756
rect 4479 28716 4620 28744
rect 4479 28713 4491 28716
rect 4433 28707 4491 28713
rect 4614 28704 4620 28716
rect 4672 28704 4678 28756
rect 8018 28704 8024 28756
rect 8076 28744 8082 28756
rect 8113 28747 8171 28753
rect 8113 28744 8125 28747
rect 8076 28716 8125 28744
rect 8076 28704 8082 28716
rect 8113 28713 8125 28716
rect 8159 28713 8171 28747
rect 8113 28707 8171 28713
rect 16390 28704 16396 28756
rect 16448 28744 16454 28756
rect 16448 28716 17264 28744
rect 16448 28704 16454 28716
rect 4062 28636 4068 28688
rect 4120 28636 4126 28688
rect 12406 28648 17172 28676
rect 4080 28608 4108 28636
rect 3988 28580 4108 28608
rect 1670 28540 1676 28552
rect 1631 28512 1676 28540
rect 1670 28500 1676 28512
rect 1728 28500 1734 28552
rect 2590 28500 2596 28552
rect 2648 28540 2654 28552
rect 3988 28549 4016 28580
rect 5626 28568 5632 28620
rect 5684 28608 5690 28620
rect 6917 28611 6975 28617
rect 6917 28608 6929 28611
rect 5684 28580 6929 28608
rect 5684 28568 5690 28580
rect 6917 28577 6929 28580
rect 6963 28608 6975 28611
rect 7006 28608 7012 28620
rect 6963 28580 7012 28608
rect 6963 28577 6975 28580
rect 6917 28571 6975 28577
rect 7006 28568 7012 28580
rect 7064 28608 7070 28620
rect 7064 28580 7880 28608
rect 7064 28568 7070 28580
rect 3789 28543 3847 28549
rect 3789 28540 3801 28543
rect 2648 28512 3801 28540
rect 2648 28500 2654 28512
rect 3789 28509 3801 28512
rect 3835 28509 3847 28543
rect 3789 28503 3847 28509
rect 3973 28543 4031 28549
rect 3973 28509 3985 28543
rect 4019 28509 4031 28543
rect 3973 28503 4031 28509
rect 4065 28543 4123 28549
rect 4065 28509 4077 28543
rect 4111 28509 4123 28543
rect 4065 28503 4123 28509
rect 4157 28543 4215 28549
rect 4157 28509 4169 28543
rect 4203 28540 4215 28543
rect 4203 28512 5948 28540
rect 4203 28509 4215 28512
rect 4157 28503 4215 28509
rect 1854 28472 1860 28484
rect 1815 28444 1860 28472
rect 1854 28432 1860 28444
rect 1912 28432 1918 28484
rect 3326 28432 3332 28484
rect 3384 28472 3390 28484
rect 4080 28472 4108 28503
rect 3384 28444 4108 28472
rect 3384 28432 3390 28444
rect 2038 28404 2044 28416
rect 1999 28376 2044 28404
rect 2038 28364 2044 28376
rect 2096 28364 2102 28416
rect 3237 28407 3295 28413
rect 3237 28373 3249 28407
rect 3283 28404 3295 28407
rect 4172 28404 4200 28503
rect 5920 28416 5948 28512
rect 7190 28500 7196 28552
rect 7248 28540 7254 28552
rect 7469 28543 7527 28549
rect 7469 28540 7481 28543
rect 7248 28512 7481 28540
rect 7248 28500 7254 28512
rect 7469 28509 7481 28512
rect 7515 28509 7527 28543
rect 7650 28540 7656 28552
rect 7611 28512 7656 28540
rect 7469 28503 7527 28509
rect 7650 28500 7656 28512
rect 7708 28500 7714 28552
rect 7852 28549 7880 28580
rect 7745 28543 7803 28549
rect 7745 28509 7757 28543
rect 7791 28509 7803 28543
rect 7745 28503 7803 28509
rect 7837 28543 7895 28549
rect 7837 28509 7849 28543
rect 7883 28509 7895 28543
rect 7837 28503 7895 28509
rect 9953 28543 10011 28549
rect 9953 28509 9965 28543
rect 9999 28540 10011 28543
rect 11054 28540 11060 28552
rect 9999 28512 11060 28540
rect 9999 28509 10011 28512
rect 9953 28503 10011 28509
rect 7006 28432 7012 28484
rect 7064 28472 7070 28484
rect 7374 28472 7380 28484
rect 7064 28444 7380 28472
rect 7064 28432 7070 28444
rect 7374 28432 7380 28444
rect 7432 28472 7438 28484
rect 7760 28472 7788 28503
rect 11054 28500 11060 28512
rect 11112 28500 11118 28552
rect 10226 28481 10232 28484
rect 7432 28444 7788 28472
rect 7432 28432 7438 28444
rect 10220 28435 10232 28481
rect 10284 28472 10290 28484
rect 10284 28444 10320 28472
rect 10226 28432 10232 28435
rect 10284 28432 10290 28444
rect 3283 28376 4200 28404
rect 3283 28373 3295 28376
rect 3237 28367 3295 28373
rect 5902 28364 5908 28416
rect 5960 28404 5966 28416
rect 6273 28407 6331 28413
rect 6273 28404 6285 28407
rect 5960 28376 6285 28404
rect 5960 28364 5966 28376
rect 6273 28373 6285 28376
rect 6319 28404 6331 28407
rect 6822 28404 6828 28416
rect 6319 28376 6828 28404
rect 6319 28373 6331 28376
rect 6273 28367 6331 28373
rect 6822 28364 6828 28376
rect 6880 28364 6886 28416
rect 9398 28404 9404 28416
rect 9359 28376 9404 28404
rect 9398 28364 9404 28376
rect 9456 28404 9462 28416
rect 10042 28404 10048 28416
rect 9456 28376 10048 28404
rect 9456 28364 9462 28376
rect 10042 28364 10048 28376
rect 10100 28364 10106 28416
rect 11146 28364 11152 28416
rect 11204 28404 11210 28416
rect 11333 28407 11391 28413
rect 11333 28404 11345 28407
rect 11204 28376 11345 28404
rect 11204 28364 11210 28376
rect 11333 28373 11345 28376
rect 11379 28404 11391 28407
rect 12406 28404 12434 28648
rect 12986 28540 12992 28552
rect 12947 28512 12992 28540
rect 12986 28500 12992 28512
rect 13044 28500 13050 28552
rect 13354 28540 13360 28552
rect 13315 28512 13360 28540
rect 13354 28500 13360 28512
rect 13412 28500 13418 28552
rect 14458 28540 14464 28552
rect 14419 28512 14464 28540
rect 14458 28500 14464 28512
rect 14516 28500 14522 28552
rect 16758 28540 16764 28552
rect 16719 28512 16764 28540
rect 16758 28500 16764 28512
rect 16816 28500 16822 28552
rect 16942 28549 16948 28552
rect 16909 28543 16948 28549
rect 16909 28509 16921 28543
rect 16909 28503 16948 28509
rect 16942 28500 16948 28503
rect 17000 28500 17006 28552
rect 17144 28549 17172 28648
rect 17236 28549 17264 28716
rect 21450 28608 21456 28620
rect 21411 28580 21456 28608
rect 21450 28568 21456 28580
rect 21508 28568 21514 28620
rect 23385 28611 23443 28617
rect 23385 28577 23397 28611
rect 23431 28608 23443 28611
rect 24026 28608 24032 28620
rect 23431 28580 24032 28608
rect 23431 28577 23443 28580
rect 23385 28571 23443 28577
rect 24026 28568 24032 28580
rect 24084 28608 24090 28620
rect 25777 28611 25835 28617
rect 25777 28608 25789 28611
rect 24084 28580 25789 28608
rect 24084 28568 24090 28580
rect 25777 28577 25789 28580
rect 25823 28577 25835 28611
rect 25777 28571 25835 28577
rect 17129 28543 17187 28549
rect 17129 28509 17141 28543
rect 17175 28509 17187 28543
rect 17129 28503 17187 28509
rect 17226 28543 17284 28549
rect 17226 28509 17238 28543
rect 17272 28540 17284 28543
rect 17865 28543 17923 28549
rect 17865 28540 17877 28543
rect 17272 28512 17877 28540
rect 17272 28509 17284 28512
rect 17226 28503 17284 28509
rect 17865 28509 17877 28512
rect 17911 28540 17923 28543
rect 17954 28540 17960 28552
rect 17911 28512 17960 28540
rect 17911 28509 17923 28512
rect 17865 28503 17923 28509
rect 17954 28500 17960 28512
rect 18012 28500 18018 28552
rect 19334 28500 19340 28552
rect 19392 28540 19398 28552
rect 20622 28540 20628 28552
rect 19392 28512 20628 28540
rect 19392 28500 19398 28512
rect 20622 28500 20628 28512
rect 20680 28540 20686 28552
rect 21468 28540 21496 28568
rect 20680 28512 21496 28540
rect 25792 28540 25820 28571
rect 28994 28540 29000 28552
rect 25792 28512 29000 28540
rect 20680 28500 20686 28512
rect 28994 28500 29000 28512
rect 29052 28500 29058 28552
rect 13170 28472 13176 28484
rect 13131 28444 13176 28472
rect 13170 28432 13176 28444
rect 13228 28432 13234 28484
rect 13262 28432 13268 28484
rect 13320 28472 13326 28484
rect 16482 28472 16488 28484
rect 13320 28444 13365 28472
rect 13556 28444 16488 28472
rect 13320 28432 13326 28444
rect 13556 28413 13584 28444
rect 16482 28432 16488 28444
rect 16540 28432 16546 28484
rect 17037 28475 17095 28481
rect 17037 28441 17049 28475
rect 17083 28472 17095 28475
rect 19058 28472 19064 28484
rect 17083 28444 19064 28472
rect 17083 28441 17095 28444
rect 17037 28435 17095 28441
rect 19058 28432 19064 28444
rect 19116 28432 19122 28484
rect 20714 28432 20720 28484
rect 20772 28472 20778 28484
rect 21186 28475 21244 28481
rect 21186 28472 21198 28475
rect 20772 28444 21198 28472
rect 20772 28432 20778 28444
rect 21186 28441 21198 28444
rect 21232 28441 21244 28475
rect 21186 28435 21244 28441
rect 22554 28432 22560 28484
rect 22612 28472 22618 28484
rect 23118 28475 23176 28481
rect 23118 28472 23130 28475
rect 22612 28444 23130 28472
rect 22612 28432 22618 28444
rect 23118 28441 23130 28444
rect 23164 28441 23176 28475
rect 23118 28435 23176 28441
rect 25682 28432 25688 28484
rect 25740 28472 25746 28484
rect 26022 28475 26080 28481
rect 26022 28472 26034 28475
rect 25740 28444 26034 28472
rect 25740 28432 25746 28444
rect 26022 28441 26034 28444
rect 26068 28441 26080 28475
rect 26022 28435 26080 28441
rect 27706 28432 27712 28484
rect 27764 28472 27770 28484
rect 28730 28475 28788 28481
rect 28730 28472 28742 28475
rect 27764 28444 28742 28472
rect 27764 28432 27770 28444
rect 28730 28441 28742 28444
rect 28776 28441 28788 28475
rect 28730 28435 28788 28441
rect 11379 28376 12434 28404
rect 13541 28407 13599 28413
rect 11379 28373 11391 28376
rect 11333 28367 11391 28373
rect 13541 28373 13553 28407
rect 13587 28373 13599 28407
rect 13541 28367 13599 28373
rect 15102 28364 15108 28416
rect 15160 28404 15166 28416
rect 15749 28407 15807 28413
rect 15749 28404 15761 28407
rect 15160 28376 15761 28404
rect 15160 28364 15166 28376
rect 15749 28373 15761 28376
rect 15795 28373 15807 28407
rect 17402 28404 17408 28416
rect 17363 28376 17408 28404
rect 15749 28367 15807 28373
rect 17402 28364 17408 28376
rect 17460 28364 17466 28416
rect 19426 28364 19432 28416
rect 19484 28404 19490 28416
rect 20073 28407 20131 28413
rect 20073 28404 20085 28407
rect 19484 28376 20085 28404
rect 19484 28364 19490 28376
rect 20073 28373 20085 28376
rect 20119 28373 20131 28407
rect 22002 28404 22008 28416
rect 21963 28376 22008 28404
rect 20073 28367 20131 28373
rect 22002 28364 22008 28376
rect 22060 28364 22066 28416
rect 26418 28364 26424 28416
rect 26476 28404 26482 28416
rect 27157 28407 27215 28413
rect 27157 28404 27169 28407
rect 26476 28376 27169 28404
rect 26476 28364 26482 28376
rect 27157 28373 27169 28376
rect 27203 28373 27215 28407
rect 27614 28404 27620 28416
rect 27575 28376 27620 28404
rect 27157 28367 27215 28373
rect 27614 28364 27620 28376
rect 27672 28364 27678 28416
rect 1104 28314 68816 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 68816 28314
rect 1104 28240 68816 28262
rect 1854 28160 1860 28212
rect 1912 28200 1918 28212
rect 6822 28200 6828 28212
rect 1912 28172 6828 28200
rect 1912 28160 1918 28172
rect 6822 28160 6828 28172
rect 6880 28160 6886 28212
rect 10137 28203 10195 28209
rect 10137 28169 10149 28203
rect 10183 28200 10195 28203
rect 10226 28200 10232 28212
rect 10183 28172 10232 28200
rect 10183 28169 10195 28172
rect 10137 28163 10195 28169
rect 10226 28160 10232 28172
rect 10284 28160 10290 28212
rect 13081 28203 13139 28209
rect 13081 28169 13093 28203
rect 13127 28200 13139 28203
rect 16758 28200 16764 28212
rect 13127 28172 16764 28200
rect 13127 28169 13139 28172
rect 13081 28163 13139 28169
rect 16758 28160 16764 28172
rect 16816 28160 16822 28212
rect 20346 28160 20352 28212
rect 20404 28160 20410 28212
rect 20714 28200 20720 28212
rect 20675 28172 20720 28200
rect 20714 28160 20720 28172
rect 20772 28160 20778 28212
rect 22005 28203 22063 28209
rect 22005 28169 22017 28203
rect 22051 28200 22063 28203
rect 22554 28200 22560 28212
rect 22051 28172 22560 28200
rect 22051 28169 22063 28172
rect 22005 28163 22063 28169
rect 22554 28160 22560 28172
rect 22612 28160 22618 28212
rect 25406 28160 25412 28212
rect 25464 28160 25470 28212
rect 25777 28203 25835 28209
rect 25777 28169 25789 28203
rect 25823 28200 25835 28203
rect 26234 28200 26240 28212
rect 25823 28172 26240 28200
rect 25823 28169 25835 28172
rect 25777 28163 25835 28169
rect 26234 28160 26240 28172
rect 26292 28160 26298 28212
rect 2406 28132 2412 28144
rect 2148 28104 2412 28132
rect 1857 28067 1915 28073
rect 1857 28033 1869 28067
rect 1903 28033 1915 28067
rect 2038 28064 2044 28076
rect 1999 28036 2044 28064
rect 1857 28027 1915 28033
rect 1872 27996 1900 28027
rect 2038 28024 2044 28036
rect 2096 28024 2102 28076
rect 2148 28073 2176 28104
rect 2406 28092 2412 28104
rect 2464 28132 2470 28144
rect 3326 28132 3332 28144
rect 2464 28104 3332 28132
rect 2464 28092 2470 28104
rect 3326 28092 3332 28104
rect 3384 28092 3390 28144
rect 5074 28092 5080 28144
rect 5132 28132 5138 28144
rect 5132 28104 9904 28132
rect 5132 28092 5138 28104
rect 2133 28067 2191 28073
rect 2133 28033 2145 28067
rect 2179 28033 2191 28067
rect 2133 28027 2191 28033
rect 2225 28067 2283 28073
rect 2225 28033 2237 28067
rect 2271 28064 2283 28067
rect 2961 28067 3019 28073
rect 2961 28064 2973 28067
rect 2271 28036 2973 28064
rect 2271 28033 2283 28036
rect 2225 28027 2283 28033
rect 2961 28033 2973 28036
rect 3007 28064 3019 28067
rect 3142 28064 3148 28076
rect 3007 28036 3148 28064
rect 3007 28033 3019 28036
rect 2961 28027 3019 28033
rect 3142 28024 3148 28036
rect 3200 28064 3206 28076
rect 7650 28064 7656 28076
rect 3200 28036 7656 28064
rect 3200 28024 3206 28036
rect 7650 28024 7656 28036
rect 7708 28024 7714 28076
rect 9490 28064 9496 28076
rect 9451 28036 9496 28064
rect 9490 28024 9496 28036
rect 9548 28024 9554 28076
rect 9674 28064 9680 28076
rect 9635 28036 9680 28064
rect 9674 28024 9680 28036
rect 9732 28024 9738 28076
rect 9876 28073 9904 28104
rect 12434 28092 12440 28144
rect 12492 28132 12498 28144
rect 12805 28135 12863 28141
rect 12805 28132 12817 28135
rect 12492 28104 12817 28132
rect 12492 28092 12498 28104
rect 12805 28101 12817 28104
rect 12851 28101 12863 28135
rect 12805 28095 12863 28101
rect 13814 28092 13820 28144
rect 13872 28132 13878 28144
rect 15102 28132 15108 28144
rect 13872 28104 15108 28132
rect 13872 28092 13878 28104
rect 15102 28092 15108 28104
rect 15160 28132 15166 28144
rect 15160 28104 15516 28132
rect 15160 28092 15166 28104
rect 9769 28067 9827 28073
rect 9769 28033 9781 28067
rect 9815 28033 9827 28067
rect 9769 28027 9827 28033
rect 9861 28067 9919 28073
rect 9861 28033 9873 28067
rect 9907 28033 9919 28067
rect 9861 28027 9919 28033
rect 12529 28067 12587 28073
rect 12529 28033 12541 28067
rect 12575 28064 12587 28067
rect 12618 28064 12624 28076
rect 12575 28036 12624 28064
rect 12575 28033 12587 28036
rect 12529 28027 12587 28033
rect 2590 27996 2596 28008
rect 1872 27968 2596 27996
rect 2590 27956 2596 27968
rect 2648 27956 2654 28008
rect 7006 27956 7012 28008
rect 7064 27996 7070 28008
rect 7558 27996 7564 28008
rect 7064 27968 7564 27996
rect 7064 27956 7070 27968
rect 7558 27956 7564 27968
rect 7616 27996 7622 28008
rect 9784 27996 9812 28027
rect 12618 28024 12624 28036
rect 12676 28024 12682 28076
rect 12713 28067 12771 28073
rect 12713 28033 12725 28067
rect 12759 28033 12771 28067
rect 12713 28027 12771 28033
rect 12897 28067 12955 28073
rect 12897 28033 12909 28067
rect 12943 28064 12955 28067
rect 13354 28064 13360 28076
rect 12943 28036 13360 28064
rect 12943 28033 12955 28036
rect 12897 28027 12955 28033
rect 9950 27996 9956 28008
rect 7616 27968 9956 27996
rect 7616 27956 7622 27968
rect 9950 27956 9956 27968
rect 10008 27956 10014 28008
rect 12728 27996 12756 28027
rect 13354 28024 13360 28036
rect 13412 28064 13418 28076
rect 13722 28064 13728 28076
rect 13412 28036 13728 28064
rect 13412 28024 13418 28036
rect 13722 28024 13728 28036
rect 13780 28024 13786 28076
rect 15217 28067 15275 28073
rect 15217 28033 15229 28067
rect 15263 28064 15275 28067
rect 15378 28064 15384 28076
rect 15263 28036 15384 28064
rect 15263 28033 15275 28036
rect 15217 28027 15275 28033
rect 15378 28024 15384 28036
rect 15436 28024 15442 28076
rect 15488 28073 15516 28104
rect 16942 28092 16948 28144
rect 17000 28132 17006 28144
rect 19245 28135 19303 28141
rect 17000 28104 19104 28132
rect 17000 28092 17006 28104
rect 15473 28067 15531 28073
rect 15473 28033 15485 28067
rect 15519 28033 15531 28067
rect 15473 28027 15531 28033
rect 18345 28067 18403 28073
rect 18345 28033 18357 28067
rect 18391 28064 18403 28067
rect 18966 28064 18972 28076
rect 18391 28036 18972 28064
rect 18391 28033 18403 28036
rect 18345 28027 18403 28033
rect 18966 28024 18972 28036
rect 19024 28024 19030 28076
rect 19076 28064 19104 28104
rect 19245 28101 19257 28135
rect 19291 28132 19303 28135
rect 19291 28104 20208 28132
rect 19291 28101 19303 28104
rect 19245 28095 19303 28101
rect 19426 28064 19432 28076
rect 19076 28036 19432 28064
rect 19426 28024 19432 28036
rect 19484 28024 19490 28076
rect 19613 28067 19671 28073
rect 19613 28033 19625 28067
rect 19659 28033 19671 28067
rect 20070 28064 20076 28076
rect 20031 28036 20076 28064
rect 19613 28027 19671 28033
rect 13170 27996 13176 28008
rect 12728 27968 13176 27996
rect 13170 27956 13176 27968
rect 13228 27996 13234 28008
rect 18601 27999 18659 28005
rect 13228 27968 13400 27996
rect 13228 27956 13234 27968
rect 13372 27940 13400 27968
rect 18601 27965 18613 27999
rect 18647 27996 18659 27999
rect 19334 27996 19340 28008
rect 18647 27968 19340 27996
rect 18647 27965 18659 27968
rect 18601 27959 18659 27965
rect 19334 27956 19340 27968
rect 19392 27956 19398 28008
rect 19628 27996 19656 28027
rect 20070 28024 20076 28036
rect 20128 28024 20134 28076
rect 20180 28067 20208 28104
rect 20364 28076 20392 28160
rect 20990 28132 20996 28144
rect 20502 28104 20996 28132
rect 20236 28070 20294 28076
rect 20236 28067 20248 28070
rect 20180 28039 20248 28067
rect 20236 28036 20248 28039
rect 20282 28036 20294 28070
rect 20236 28030 20294 28036
rect 20336 28070 20394 28076
rect 20502 28073 20530 28104
rect 20990 28092 20996 28104
rect 21048 28092 21054 28144
rect 22186 28092 22192 28144
rect 22244 28132 22250 28144
rect 22244 28104 22416 28132
rect 22244 28092 22250 28104
rect 20336 28036 20348 28070
rect 20382 28036 20394 28070
rect 20336 28030 20394 28036
rect 20487 28067 20545 28073
rect 20487 28033 20499 28067
rect 20533 28033 20545 28067
rect 21818 28064 21824 28076
rect 20487 28027 20545 28033
rect 20640 28036 21824 28064
rect 20640 27996 20668 28036
rect 21818 28024 21824 28036
rect 21876 28024 21882 28076
rect 22388 28073 22416 28104
rect 25424 28079 25452 28160
rect 28994 28092 29000 28144
rect 29052 28132 29058 28144
rect 30282 28132 30288 28144
rect 29052 28104 30288 28132
rect 29052 28092 29058 28104
rect 30282 28092 30288 28104
rect 30340 28132 30346 28144
rect 30340 28104 30696 28132
rect 30340 28092 30346 28104
rect 22281 28067 22339 28073
rect 22281 28033 22293 28067
rect 22327 28033 22339 28067
rect 22281 28027 22339 28033
rect 22373 28067 22431 28073
rect 22373 28033 22385 28067
rect 22419 28033 22431 28067
rect 22373 28027 22431 28033
rect 21266 27996 21272 28008
rect 19628 27968 20668 27996
rect 21179 27968 21272 27996
rect 21266 27956 21272 27968
rect 21324 27996 21330 28008
rect 22296 27996 22324 28027
rect 22462 28024 22468 28076
rect 22520 28064 22526 28076
rect 22649 28067 22707 28073
rect 22520 28036 22565 28064
rect 22520 28024 22526 28036
rect 22649 28033 22661 28067
rect 22695 28033 22707 28067
rect 25130 28064 25136 28076
rect 25091 28036 25136 28064
rect 22649 28027 22707 28033
rect 22554 27996 22560 28008
rect 21324 27968 22560 27996
rect 21324 27956 21330 27968
rect 22554 27956 22560 27968
rect 22612 27956 22618 28008
rect 13354 27888 13360 27940
rect 13412 27888 13418 27940
rect 20070 27888 20076 27940
rect 20128 27928 20134 27940
rect 20530 27928 20536 27940
rect 20128 27900 20536 27928
rect 20128 27888 20134 27900
rect 20530 27888 20536 27900
rect 20588 27928 20594 27940
rect 22664 27928 22692 28027
rect 25130 28024 25136 28036
rect 25188 28024 25194 28076
rect 25412 28073 25470 28079
rect 25312 28067 25370 28073
rect 25312 28064 25324 28067
rect 25251 28036 25324 28064
rect 20588 27900 22692 27928
rect 25251 27928 25279 28036
rect 25312 28033 25324 28036
rect 25358 28033 25370 28067
rect 25412 28039 25424 28073
rect 25458 28039 25470 28073
rect 25412 28033 25470 28039
rect 25501 28067 25559 28073
rect 25501 28033 25513 28067
rect 25547 28039 25636 28067
rect 25547 28033 25559 28039
rect 25312 28027 25370 28033
rect 25501 28027 25559 28033
rect 25314 27928 25320 27940
rect 25251 27900 25320 27928
rect 20588 27888 20594 27900
rect 25314 27888 25320 27900
rect 25372 27888 25378 27940
rect 2501 27863 2559 27869
rect 2501 27829 2513 27863
rect 2547 27860 2559 27863
rect 2866 27860 2872 27872
rect 2547 27832 2872 27860
rect 2547 27829 2559 27832
rect 2501 27823 2559 27829
rect 2866 27820 2872 27832
rect 2924 27820 2930 27872
rect 7190 27860 7196 27872
rect 7151 27832 7196 27860
rect 7190 27820 7196 27832
rect 7248 27820 7254 27872
rect 13446 27820 13452 27872
rect 13504 27860 13510 27872
rect 13541 27863 13599 27869
rect 13541 27860 13553 27863
rect 13504 27832 13553 27860
rect 13504 27820 13510 27832
rect 13541 27829 13553 27832
rect 13587 27829 13599 27863
rect 14090 27860 14096 27872
rect 14003 27832 14096 27860
rect 13541 27823 13599 27829
rect 14090 27820 14096 27832
rect 14148 27860 14154 27872
rect 14826 27860 14832 27872
rect 14148 27832 14832 27860
rect 14148 27820 14154 27832
rect 14826 27820 14832 27832
rect 14884 27820 14890 27872
rect 15102 27820 15108 27872
rect 15160 27860 15166 27872
rect 15933 27863 15991 27869
rect 15933 27860 15945 27863
rect 15160 27832 15945 27860
rect 15160 27820 15166 27832
rect 15933 27829 15945 27832
rect 15979 27860 15991 27863
rect 16206 27860 16212 27872
rect 15979 27832 16212 27860
rect 15979 27829 15991 27832
rect 15933 27823 15991 27829
rect 16206 27820 16212 27832
rect 16264 27820 16270 27872
rect 16574 27820 16580 27872
rect 16632 27860 16638 27872
rect 16669 27863 16727 27869
rect 16669 27860 16681 27863
rect 16632 27832 16681 27860
rect 16632 27820 16638 27832
rect 16669 27829 16681 27832
rect 16715 27829 16727 27863
rect 16669 27823 16727 27829
rect 17221 27863 17279 27869
rect 17221 27829 17233 27863
rect 17267 27860 17279 27863
rect 17954 27860 17960 27872
rect 17267 27832 17960 27860
rect 17267 27829 17279 27832
rect 17221 27823 17279 27829
rect 17954 27820 17960 27832
rect 18012 27820 18018 27872
rect 19886 27820 19892 27872
rect 19944 27860 19950 27872
rect 21266 27860 21272 27872
rect 19944 27832 21272 27860
rect 19944 27820 19950 27832
rect 21266 27820 21272 27832
rect 21324 27820 21330 27872
rect 22554 27820 22560 27872
rect 22612 27860 22618 27872
rect 23201 27863 23259 27869
rect 23201 27860 23213 27863
rect 22612 27832 23213 27860
rect 22612 27820 22618 27832
rect 23201 27829 23213 27832
rect 23247 27860 23259 27863
rect 23566 27860 23572 27872
rect 23247 27832 23572 27860
rect 23247 27829 23259 27832
rect 23201 27823 23259 27829
rect 23566 27820 23572 27832
rect 23624 27820 23630 27872
rect 24670 27820 24676 27872
rect 24728 27860 24734 27872
rect 25608 27860 25636 28039
rect 29178 28024 29184 28076
rect 29236 28064 29242 28076
rect 30668 28073 30696 28104
rect 30386 28067 30444 28073
rect 30386 28064 30398 28067
rect 29236 28036 30398 28064
rect 29236 28024 29242 28036
rect 30386 28033 30398 28036
rect 30432 28033 30444 28067
rect 30386 28027 30444 28033
rect 30653 28067 30711 28073
rect 30653 28033 30665 28067
rect 30699 28033 30711 28067
rect 30653 28027 30711 28033
rect 67634 27928 67640 27940
rect 67595 27900 67640 27928
rect 67634 27888 67640 27900
rect 67692 27888 67698 27940
rect 26237 27863 26295 27869
rect 26237 27860 26249 27863
rect 24728 27832 26249 27860
rect 24728 27820 24734 27832
rect 26237 27829 26249 27832
rect 26283 27860 26295 27863
rect 26326 27860 26332 27872
rect 26283 27832 26332 27860
rect 26283 27829 26295 27832
rect 26237 27823 26295 27829
rect 26326 27820 26332 27832
rect 26384 27820 26390 27872
rect 29270 27860 29276 27872
rect 29231 27832 29276 27860
rect 29270 27820 29276 27832
rect 29328 27820 29334 27872
rect 1104 27770 68816 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 65654 27770
rect 65706 27718 65718 27770
rect 65770 27718 65782 27770
rect 65834 27718 65846 27770
rect 65898 27718 65910 27770
rect 65962 27718 68816 27770
rect 1104 27696 68816 27718
rect 2866 27616 2872 27668
rect 2924 27656 2930 27668
rect 2924 27628 5488 27656
rect 2924 27616 2930 27628
rect 3326 27480 3332 27532
rect 3384 27520 3390 27532
rect 5460 27520 5488 27628
rect 9674 27616 9680 27668
rect 9732 27656 9738 27668
rect 10045 27659 10103 27665
rect 10045 27656 10057 27659
rect 9732 27628 10057 27656
rect 9732 27616 9738 27628
rect 10045 27625 10057 27628
rect 10091 27625 10103 27659
rect 10045 27619 10103 27625
rect 13446 27616 13452 27668
rect 13504 27656 13510 27668
rect 13504 27628 14228 27656
rect 13504 27616 13510 27628
rect 14093 27591 14151 27597
rect 14093 27588 14105 27591
rect 12406 27560 14105 27588
rect 7742 27520 7748 27532
rect 3384 27492 4108 27520
rect 5460 27492 5580 27520
rect 3384 27480 3390 27492
rect 1670 27412 1676 27464
rect 1728 27412 1734 27464
rect 2225 27455 2283 27461
rect 2225 27421 2237 27455
rect 2271 27452 2283 27455
rect 2314 27452 2320 27464
rect 2271 27424 2320 27452
rect 2271 27421 2283 27424
rect 2225 27415 2283 27421
rect 2314 27412 2320 27424
rect 2372 27412 2378 27464
rect 2590 27412 2596 27464
rect 2648 27452 2654 27464
rect 4080 27461 4108 27492
rect 3789 27455 3847 27461
rect 3789 27452 3801 27455
rect 2648 27424 3801 27452
rect 2648 27412 2654 27424
rect 3789 27421 3801 27424
rect 3835 27421 3847 27455
rect 3789 27415 3847 27421
rect 3973 27455 4031 27461
rect 3973 27421 3985 27455
rect 4019 27421 4031 27455
rect 3973 27415 4031 27421
rect 4065 27455 4123 27461
rect 4065 27421 4077 27455
rect 4111 27421 4123 27455
rect 4065 27415 4123 27421
rect 4157 27455 4215 27461
rect 4157 27421 4169 27455
rect 4203 27452 4215 27455
rect 5074 27452 5080 27464
rect 4203 27424 5080 27452
rect 4203 27421 4215 27424
rect 4157 27415 4215 27421
rect 1688 27384 1716 27412
rect 2130 27384 2136 27396
rect 1688 27356 2136 27384
rect 2130 27344 2136 27356
rect 2188 27384 2194 27396
rect 2869 27387 2927 27393
rect 2869 27384 2881 27387
rect 2188 27356 2881 27384
rect 2188 27344 2194 27356
rect 2869 27353 2881 27356
rect 2915 27353 2927 27387
rect 3050 27384 3056 27396
rect 3011 27356 3056 27384
rect 2869 27347 2927 27353
rect 3050 27344 3056 27356
rect 3108 27344 3114 27396
rect 3237 27387 3295 27393
rect 3237 27353 3249 27387
rect 3283 27384 3295 27387
rect 3988 27384 4016 27415
rect 5074 27412 5080 27424
rect 5132 27412 5138 27464
rect 5442 27452 5448 27464
rect 5403 27424 5448 27452
rect 5442 27412 5448 27424
rect 5500 27412 5506 27464
rect 5552 27452 5580 27492
rect 7300 27492 7748 27520
rect 7300 27461 7328 27492
rect 7742 27480 7748 27492
rect 7800 27520 7806 27532
rect 9490 27520 9496 27532
rect 7800 27492 9496 27520
rect 7800 27480 7806 27492
rect 9490 27480 9496 27492
rect 9548 27480 9554 27532
rect 11054 27520 11060 27532
rect 11015 27492 11060 27520
rect 11054 27480 11060 27492
rect 11112 27480 11118 27532
rect 5701 27455 5759 27461
rect 5701 27452 5713 27455
rect 5552 27424 5713 27452
rect 5701 27421 5713 27424
rect 5747 27421 5759 27455
rect 5701 27415 5759 27421
rect 7285 27455 7343 27461
rect 7285 27421 7297 27455
rect 7331 27421 7343 27455
rect 7466 27452 7472 27464
rect 7427 27424 7472 27452
rect 7285 27415 7343 27421
rect 7466 27412 7472 27424
rect 7524 27412 7530 27464
rect 7564 27449 7622 27455
rect 7564 27440 7576 27449
rect 7610 27440 7622 27449
rect 7558 27388 7564 27440
rect 7616 27388 7622 27440
rect 7650 27412 7656 27464
rect 7708 27452 7714 27464
rect 9861 27455 9919 27461
rect 7708 27424 7753 27452
rect 7852 27424 9812 27452
rect 7708 27412 7714 27424
rect 7852 27384 7880 27424
rect 3283 27356 4016 27384
rect 7760 27356 7880 27384
rect 3283 27353 3295 27356
rect 3237 27347 3295 27353
rect 1670 27276 1676 27328
rect 1728 27316 1734 27328
rect 2041 27319 2099 27325
rect 2041 27316 2053 27319
rect 1728 27288 2053 27316
rect 1728 27276 1734 27288
rect 2041 27285 2053 27288
rect 2087 27285 2099 27319
rect 4430 27316 4436 27328
rect 4391 27288 4436 27316
rect 2041 27279 2099 27285
rect 4430 27276 4436 27288
rect 4488 27276 4494 27328
rect 6822 27316 6828 27328
rect 6735 27288 6828 27316
rect 6822 27276 6828 27288
rect 6880 27316 6886 27328
rect 7760 27316 7788 27356
rect 9214 27344 9220 27396
rect 9272 27384 9278 27396
rect 9677 27387 9735 27393
rect 9677 27384 9689 27387
rect 9272 27356 9689 27384
rect 9272 27344 9278 27356
rect 9677 27353 9689 27356
rect 9723 27353 9735 27387
rect 9784 27384 9812 27424
rect 9861 27421 9873 27455
rect 9907 27452 9919 27455
rect 11146 27452 11152 27464
rect 9907 27424 11152 27452
rect 9907 27421 9919 27424
rect 9861 27415 9919 27421
rect 11146 27412 11152 27424
rect 11204 27412 11210 27464
rect 11324 27455 11382 27461
rect 11324 27421 11336 27455
rect 11370 27452 11382 27455
rect 12406 27452 12434 27560
rect 14093 27557 14105 27560
rect 14139 27557 14151 27591
rect 14093 27551 14151 27557
rect 11370 27424 12434 27452
rect 13357 27455 13415 27461
rect 11370 27421 11382 27424
rect 11324 27415 11382 27421
rect 13357 27421 13369 27455
rect 13403 27452 13415 27455
rect 14090 27452 14096 27464
rect 13403 27424 14096 27452
rect 13403 27421 13415 27424
rect 13357 27415 13415 27421
rect 14090 27412 14096 27424
rect 14148 27412 14154 27464
rect 14200 27452 14228 27628
rect 17034 27616 17040 27668
rect 17092 27656 17098 27668
rect 17678 27656 17684 27668
rect 17092 27628 17684 27656
rect 17092 27616 17098 27628
rect 17678 27616 17684 27628
rect 17736 27656 17742 27668
rect 19886 27656 19892 27668
rect 17736 27628 19892 27656
rect 17736 27616 17742 27628
rect 19886 27616 19892 27628
rect 19944 27616 19950 27668
rect 20990 27616 20996 27668
rect 21048 27656 21054 27668
rect 21453 27659 21511 27665
rect 21453 27656 21465 27659
rect 21048 27628 21465 27656
rect 21048 27616 21054 27628
rect 21453 27625 21465 27628
rect 21499 27656 21511 27659
rect 24670 27656 24676 27668
rect 21499 27628 24676 27656
rect 21499 27625 21511 27628
rect 21453 27619 21511 27625
rect 24670 27616 24676 27628
rect 24728 27616 24734 27668
rect 25682 27656 25688 27668
rect 25251 27628 25543 27656
rect 25643 27628 25688 27656
rect 22002 27588 22008 27600
rect 17052 27560 22008 27588
rect 16298 27520 16304 27532
rect 14476 27492 15056 27520
rect 16259 27492 16304 27520
rect 14476 27461 14504 27492
rect 15028 27464 15056 27492
rect 16298 27480 16304 27492
rect 16356 27480 16362 27532
rect 14369 27455 14427 27461
rect 14369 27452 14381 27455
rect 14200 27424 14381 27452
rect 14369 27421 14381 27424
rect 14415 27421 14427 27455
rect 14369 27415 14427 27421
rect 14461 27455 14519 27461
rect 14461 27421 14473 27455
rect 14507 27421 14519 27455
rect 14461 27415 14519 27421
rect 14550 27412 14556 27464
rect 14608 27452 14614 27464
rect 14608 27424 14653 27452
rect 14608 27412 14614 27424
rect 14734 27412 14740 27464
rect 14792 27452 14798 27464
rect 14792 27424 14837 27452
rect 14792 27412 14798 27424
rect 15010 27412 15016 27464
rect 15068 27452 15074 27464
rect 16025 27455 16083 27461
rect 16025 27452 16037 27455
rect 15068 27424 16037 27452
rect 15068 27412 15074 27424
rect 16025 27421 16037 27424
rect 16071 27421 16083 27455
rect 16025 27415 16083 27421
rect 16482 27412 16488 27464
rect 16540 27452 16546 27464
rect 16761 27455 16819 27461
rect 16761 27452 16773 27455
rect 16540 27424 16773 27452
rect 16540 27412 16546 27424
rect 16761 27421 16773 27424
rect 16807 27421 16819 27455
rect 16761 27415 16819 27421
rect 16909 27455 16967 27461
rect 16909 27421 16921 27455
rect 16955 27452 16967 27455
rect 17052 27452 17080 27560
rect 22002 27548 22008 27560
rect 22060 27588 22066 27600
rect 23842 27588 23848 27600
rect 22060 27560 22324 27588
rect 22060 27548 22066 27560
rect 19334 27520 19340 27532
rect 19247 27492 19340 27520
rect 19334 27480 19340 27492
rect 19392 27520 19398 27532
rect 20165 27523 20223 27529
rect 20165 27520 20177 27523
rect 19392 27492 20177 27520
rect 19392 27480 19398 27492
rect 20165 27489 20177 27492
rect 20211 27489 20223 27523
rect 20165 27483 20223 27489
rect 20346 27480 20352 27532
rect 20404 27520 20410 27532
rect 20441 27523 20499 27529
rect 20441 27520 20453 27523
rect 20404 27492 20453 27520
rect 20404 27480 20410 27492
rect 20441 27489 20453 27492
rect 20487 27520 20499 27523
rect 22186 27520 22192 27532
rect 20487 27492 22192 27520
rect 20487 27489 20499 27492
rect 20441 27483 20499 27489
rect 22186 27480 22192 27492
rect 22244 27480 22250 27532
rect 17218 27452 17224 27464
rect 17276 27461 17282 27464
rect 16955 27424 17080 27452
rect 17184 27424 17224 27452
rect 16955 27421 16967 27424
rect 16909 27415 16967 27421
rect 17218 27412 17224 27424
rect 17276 27415 17284 27461
rect 17276 27412 17282 27415
rect 18138 27412 18144 27464
rect 18196 27452 18202 27464
rect 19058 27452 19064 27464
rect 18196 27424 19064 27452
rect 18196 27412 18202 27424
rect 19058 27412 19064 27424
rect 19116 27452 19122 27464
rect 19245 27455 19303 27461
rect 19245 27452 19257 27455
rect 19116 27424 19257 27452
rect 19116 27412 19122 27424
rect 19245 27421 19257 27424
rect 19291 27421 19303 27455
rect 19245 27415 19303 27421
rect 19429 27455 19487 27461
rect 19429 27421 19441 27455
rect 19475 27421 19487 27455
rect 19429 27415 19487 27421
rect 13262 27384 13268 27396
rect 9784 27356 13268 27384
rect 9677 27347 9735 27353
rect 13262 27344 13268 27356
rect 13320 27344 13326 27396
rect 13541 27387 13599 27393
rect 13541 27353 13553 27387
rect 13587 27384 13599 27387
rect 14642 27384 14648 27396
rect 13587 27356 14648 27384
rect 13587 27353 13599 27356
rect 13541 27347 13599 27353
rect 14642 27344 14648 27356
rect 14700 27344 14706 27396
rect 17034 27384 17040 27396
rect 16995 27356 17040 27384
rect 17034 27344 17040 27356
rect 17092 27344 17098 27396
rect 17126 27344 17132 27396
rect 17184 27384 17190 27396
rect 17957 27387 18015 27393
rect 17957 27384 17969 27387
rect 17184 27356 17229 27384
rect 17328 27356 17969 27384
rect 17184 27344 17190 27356
rect 7926 27316 7932 27328
rect 6880 27288 7788 27316
rect 7887 27288 7932 27316
rect 6880 27276 6886 27288
rect 7926 27276 7932 27288
rect 7984 27276 7990 27328
rect 12437 27319 12495 27325
rect 12437 27285 12449 27319
rect 12483 27316 12495 27319
rect 12618 27316 12624 27328
rect 12483 27288 12624 27316
rect 12483 27285 12495 27288
rect 12437 27279 12495 27285
rect 12618 27276 12624 27288
rect 12676 27276 12682 27328
rect 13173 27319 13231 27325
rect 13173 27285 13185 27319
rect 13219 27316 13231 27319
rect 15930 27316 15936 27328
rect 13219 27288 15936 27316
rect 13219 27285 13231 27288
rect 13173 27279 13231 27285
rect 15930 27276 15936 27288
rect 15988 27276 15994 27328
rect 16022 27276 16028 27328
rect 16080 27316 16086 27328
rect 17328 27316 17356 27356
rect 17957 27353 17969 27356
rect 18003 27353 18015 27387
rect 17957 27347 18015 27353
rect 16080 27288 17356 27316
rect 17405 27319 17463 27325
rect 16080 27276 16086 27288
rect 17405 27285 17417 27319
rect 17451 27316 17463 27319
rect 17770 27316 17776 27328
rect 17451 27288 17776 27316
rect 17451 27285 17463 27288
rect 17405 27279 17463 27285
rect 17770 27276 17776 27288
rect 17828 27276 17834 27328
rect 17972 27316 18000 27347
rect 18046 27344 18052 27396
rect 18104 27384 18110 27396
rect 19444 27384 19472 27415
rect 21818 27412 21824 27464
rect 21876 27452 21882 27464
rect 22296 27461 22324 27560
rect 23492 27560 23612 27588
rect 23803 27560 23848 27588
rect 22462 27520 22468 27532
rect 22423 27492 22468 27520
rect 22462 27480 22468 27492
rect 22520 27480 22526 27532
rect 22097 27455 22155 27461
rect 22097 27452 22109 27455
rect 21876 27424 22109 27452
rect 21876 27412 21882 27424
rect 22097 27421 22109 27424
rect 22143 27421 22155 27455
rect 22097 27415 22155 27421
rect 22281 27455 22339 27461
rect 22281 27421 22293 27455
rect 22327 27421 22339 27455
rect 23198 27452 23204 27464
rect 23159 27424 23204 27452
rect 22281 27415 22339 27421
rect 23198 27412 23204 27424
rect 23256 27412 23262 27464
rect 23492 27461 23520 27560
rect 23584 27520 23612 27560
rect 23842 27548 23848 27560
rect 23900 27548 23906 27600
rect 24581 27591 24639 27597
rect 24581 27557 24593 27591
rect 24627 27588 24639 27591
rect 24854 27588 24860 27600
rect 24627 27560 24860 27588
rect 24627 27557 24639 27560
rect 24581 27551 24639 27557
rect 24854 27548 24860 27560
rect 24912 27588 24918 27600
rect 25251 27588 25279 27628
rect 25406 27588 25412 27600
rect 24912 27560 25279 27588
rect 25332 27560 25412 27588
rect 24912 27548 24918 27560
rect 24946 27520 24952 27532
rect 23584 27492 24952 27520
rect 24946 27480 24952 27492
rect 25004 27520 25010 27532
rect 25332 27520 25360 27560
rect 25406 27548 25412 27560
rect 25464 27548 25470 27600
rect 25004 27492 25360 27520
rect 25004 27480 25010 27492
rect 23364 27455 23422 27461
rect 23364 27452 23376 27455
rect 23308 27424 23376 27452
rect 18104 27356 19472 27384
rect 18104 27344 18110 27356
rect 18598 27316 18604 27328
rect 17972 27288 18604 27316
rect 18598 27276 18604 27288
rect 18656 27276 18662 27328
rect 23308 27316 23336 27424
rect 23364 27421 23376 27424
rect 23410 27421 23422 27455
rect 23364 27415 23422 27421
rect 23464 27455 23522 27461
rect 23464 27421 23476 27455
rect 23510 27421 23522 27455
rect 23464 27415 23522 27421
rect 23566 27412 23572 27464
rect 23624 27452 23630 27464
rect 23624 27424 23669 27452
rect 23624 27412 23630 27424
rect 24210 27412 24216 27464
rect 24268 27452 24274 27464
rect 25041 27455 25099 27461
rect 25041 27452 25053 27455
rect 24268 27424 25053 27452
rect 24268 27412 24274 27424
rect 25041 27421 25053 27424
rect 25087 27452 25099 27455
rect 25130 27452 25136 27464
rect 25087 27424 25136 27452
rect 25087 27421 25099 27424
rect 25041 27415 25099 27421
rect 25130 27412 25136 27424
rect 25188 27412 25194 27464
rect 25332 27461 25360 27492
rect 25225 27455 25283 27461
rect 25225 27421 25237 27455
rect 25271 27421 25283 27455
rect 25225 27415 25283 27421
rect 25317 27455 25375 27461
rect 25317 27421 25329 27455
rect 25363 27421 25375 27455
rect 25317 27415 25375 27421
rect 25409 27455 25467 27461
rect 25409 27421 25421 27455
rect 25455 27452 25467 27455
rect 25515 27452 25543 27628
rect 25682 27616 25688 27628
rect 25740 27616 25746 27668
rect 28261 27591 28319 27597
rect 28261 27557 28273 27591
rect 28307 27588 28319 27591
rect 29178 27588 29184 27600
rect 28307 27560 29184 27588
rect 28307 27557 28319 27560
rect 28261 27551 28319 27557
rect 29178 27548 29184 27560
rect 29236 27548 29242 27600
rect 27430 27480 27436 27532
rect 27488 27520 27494 27532
rect 27488 27492 27927 27520
rect 27488 27480 27494 27492
rect 26050 27452 26056 27464
rect 25455 27424 26056 27452
rect 25455 27421 25467 27424
rect 25409 27415 25467 27421
rect 25235 27384 25263 27415
rect 26050 27412 26056 27424
rect 26108 27412 26114 27464
rect 26786 27412 26792 27464
rect 26844 27452 26850 27464
rect 27899 27461 27927 27492
rect 27617 27455 27675 27461
rect 27617 27452 27629 27455
rect 26844 27424 27629 27452
rect 26844 27412 26850 27424
rect 27617 27421 27629 27424
rect 27663 27421 27675 27455
rect 27780 27455 27838 27461
rect 27780 27452 27792 27455
rect 27617 27415 27675 27421
rect 27724 27424 27792 27452
rect 26142 27384 26148 27396
rect 25235 27356 25543 27384
rect 26103 27356 26148 27384
rect 23474 27316 23480 27328
rect 23308 27288 23480 27316
rect 23474 27276 23480 27288
rect 23532 27276 23538 27328
rect 25515 27316 25543 27356
rect 26142 27344 26148 27356
rect 26200 27344 26206 27396
rect 26329 27387 26387 27393
rect 26329 27353 26341 27387
rect 26375 27384 26387 27387
rect 26418 27384 26424 27396
rect 26375 27356 26424 27384
rect 26375 27353 26387 27356
rect 26329 27347 26387 27353
rect 26418 27344 26424 27356
rect 26476 27344 26482 27396
rect 27522 27344 27528 27396
rect 27580 27384 27586 27396
rect 27724 27384 27752 27424
rect 27780 27421 27792 27424
rect 27826 27421 27838 27455
rect 27780 27415 27838 27421
rect 27880 27455 27938 27461
rect 27880 27421 27892 27455
rect 27926 27421 27938 27455
rect 27880 27415 27938 27421
rect 27985 27455 28043 27461
rect 27985 27421 27997 27455
rect 28031 27421 28043 27455
rect 27985 27415 28043 27421
rect 27580 27356 27752 27384
rect 27580 27344 27586 27356
rect 26513 27319 26571 27325
rect 26513 27316 26525 27319
rect 25515 27288 26525 27316
rect 26513 27285 26525 27288
rect 26559 27285 26571 27319
rect 26513 27279 26571 27285
rect 26878 27276 26884 27328
rect 26936 27316 26942 27328
rect 27065 27319 27123 27325
rect 27065 27316 27077 27319
rect 26936 27288 27077 27316
rect 26936 27276 26942 27288
rect 27065 27285 27077 27288
rect 27111 27316 27123 27319
rect 28000 27316 28028 27415
rect 27111 27288 28028 27316
rect 27111 27285 27123 27288
rect 27065 27279 27123 27285
rect 1104 27226 68816 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 68816 27226
rect 1104 27152 68816 27174
rect 2130 27112 2136 27124
rect 2091 27084 2136 27112
rect 2130 27072 2136 27084
rect 2188 27072 2194 27124
rect 2314 27072 2320 27124
rect 2372 27112 2378 27124
rect 2372 27084 2774 27112
rect 2372 27072 2378 27084
rect 2746 27044 2774 27084
rect 3050 27072 3056 27124
rect 3108 27112 3114 27124
rect 5445 27115 5503 27121
rect 5445 27112 5457 27115
rect 3108 27084 5457 27112
rect 3108 27072 3114 27084
rect 5445 27081 5457 27084
rect 5491 27112 5503 27115
rect 5491 27084 7052 27112
rect 5491 27081 5503 27084
rect 5445 27075 5503 27081
rect 4332 27047 4390 27053
rect 2746 27016 4292 27044
rect 2314 26976 2320 26988
rect 2275 26948 2320 26976
rect 2314 26936 2320 26948
rect 2372 26936 2378 26988
rect 3326 26976 3332 26988
rect 3287 26948 3332 26976
rect 3326 26936 3332 26948
rect 3384 26936 3390 26988
rect 4264 26976 4292 27016
rect 4332 27013 4344 27047
rect 4378 27044 4390 27047
rect 4430 27044 4436 27056
rect 4378 27016 4436 27044
rect 4378 27013 4390 27016
rect 4332 27007 4390 27013
rect 4430 27004 4436 27016
rect 4488 27004 4494 27056
rect 5350 26976 5356 26988
rect 4264 26948 5356 26976
rect 5350 26936 5356 26948
rect 5408 26936 5414 26988
rect 6917 26979 6975 26985
rect 6917 26945 6929 26979
rect 6963 26945 6975 26979
rect 7024 26976 7052 27084
rect 7466 27072 7472 27124
rect 7524 27112 7530 27124
rect 9401 27115 9459 27121
rect 9401 27112 9413 27115
rect 7524 27084 9413 27112
rect 7524 27072 7530 27084
rect 9401 27081 9413 27084
rect 9447 27081 9459 27115
rect 9401 27075 9459 27081
rect 12805 27115 12863 27121
rect 12805 27081 12817 27115
rect 12851 27112 12863 27115
rect 14550 27112 14556 27124
rect 12851 27084 14556 27112
rect 12851 27081 12863 27084
rect 12805 27075 12863 27081
rect 14550 27072 14556 27084
rect 14608 27072 14614 27124
rect 14642 27072 14648 27124
rect 14700 27112 14706 27124
rect 14700 27084 14745 27112
rect 14936 27084 15240 27112
rect 14700 27072 14706 27084
rect 7828 27047 7886 27053
rect 7828 27013 7840 27047
rect 7874 27044 7886 27047
rect 7926 27044 7932 27056
rect 7874 27016 7932 27044
rect 7874 27013 7886 27016
rect 7828 27007 7886 27013
rect 7926 27004 7932 27016
rect 7984 27004 7990 27056
rect 12342 27044 12348 27056
rect 8036 27016 12348 27044
rect 8036 26976 8064 27016
rect 12342 27004 12348 27016
rect 12400 27004 12406 27056
rect 12618 27044 12624 27056
rect 12579 27016 12624 27044
rect 12618 27004 12624 27016
rect 12676 27044 12682 27056
rect 12676 27016 13308 27044
rect 12676 27004 12682 27016
rect 9582 26976 9588 26988
rect 7024 26948 8064 26976
rect 9543 26948 9588 26976
rect 6917 26939 6975 26945
rect 3602 26908 3608 26920
rect 3563 26880 3608 26908
rect 3602 26868 3608 26880
rect 3660 26868 3666 26920
rect 4062 26908 4068 26920
rect 4023 26880 4068 26908
rect 4062 26868 4068 26880
rect 4120 26868 4126 26920
rect 6932 26908 6960 26939
rect 9582 26936 9588 26948
rect 9640 26936 9646 26988
rect 9769 26979 9827 26985
rect 9769 26945 9781 26979
rect 9815 26945 9827 26979
rect 9769 26939 9827 26945
rect 12437 26979 12495 26985
rect 12437 26945 12449 26979
rect 12483 26976 12495 26979
rect 12986 26976 12992 26988
rect 12483 26948 12992 26976
rect 12483 26945 12495 26948
rect 12437 26939 12495 26945
rect 7098 26908 7104 26920
rect 6932 26880 7104 26908
rect 7098 26868 7104 26880
rect 7156 26868 7162 26920
rect 7561 26911 7619 26917
rect 7561 26877 7573 26911
rect 7607 26877 7619 26911
rect 7561 26871 7619 26877
rect 7101 26775 7159 26781
rect 7101 26741 7113 26775
rect 7147 26772 7159 26775
rect 7466 26772 7472 26784
rect 7147 26744 7472 26772
rect 7147 26741 7159 26744
rect 7101 26735 7159 26741
rect 7466 26732 7472 26744
rect 7524 26732 7530 26784
rect 7576 26772 7604 26871
rect 9214 26868 9220 26920
rect 9272 26908 9278 26920
rect 9784 26908 9812 26939
rect 12986 26936 12992 26948
rect 13044 26936 13050 26988
rect 13280 26985 13308 27016
rect 13354 27004 13360 27056
rect 13412 27044 13418 27056
rect 13449 27047 13507 27053
rect 13449 27044 13461 27047
rect 13412 27016 13461 27044
rect 13412 27004 13418 27016
rect 13449 27013 13461 27016
rect 13495 27044 13507 27047
rect 14274 27044 14280 27056
rect 13495 27016 14280 27044
rect 13495 27013 13507 27016
rect 13449 27007 13507 27013
rect 14274 27004 14280 27016
rect 14332 27004 14338 27056
rect 13265 26979 13323 26985
rect 13265 26945 13277 26979
rect 13311 26945 13323 26979
rect 13541 26979 13599 26985
rect 13541 26976 13553 26979
rect 13265 26939 13323 26945
rect 13372 26948 13553 26976
rect 9272 26880 9812 26908
rect 9272 26868 9278 26880
rect 8941 26843 8999 26849
rect 8941 26809 8953 26843
rect 8987 26840 8999 26843
rect 9582 26840 9588 26852
rect 8987 26812 9588 26840
rect 8987 26809 8999 26812
rect 8941 26803 8999 26809
rect 9582 26800 9588 26812
rect 9640 26800 9646 26852
rect 9674 26800 9680 26852
rect 9732 26840 9738 26852
rect 13372 26840 13400 26948
rect 13541 26945 13553 26948
rect 13587 26945 13599 26979
rect 13541 26939 13599 26945
rect 13633 26979 13691 26985
rect 13633 26945 13645 26979
rect 13679 26976 13691 26979
rect 13722 26976 13728 26988
rect 13679 26948 13728 26976
rect 13679 26945 13691 26948
rect 13633 26939 13691 26945
rect 13722 26936 13728 26948
rect 13780 26936 13786 26988
rect 14829 26979 14887 26985
rect 14829 26945 14841 26979
rect 14875 26976 14887 26979
rect 14936 26976 14964 27084
rect 15212 27044 15240 27084
rect 15378 27072 15384 27124
rect 15436 27112 15442 27124
rect 15473 27115 15531 27121
rect 15473 27112 15485 27115
rect 15436 27084 15485 27112
rect 15436 27072 15442 27084
rect 15473 27081 15485 27084
rect 15519 27081 15531 27115
rect 17494 27112 17500 27124
rect 15473 27075 15531 27081
rect 15580 27084 17500 27112
rect 15580 27056 15608 27084
rect 17494 27072 17500 27084
rect 17552 27072 17558 27124
rect 18966 27112 18972 27124
rect 18927 27084 18972 27112
rect 18966 27072 18972 27084
rect 19024 27072 19030 27124
rect 19058 27072 19064 27124
rect 19116 27112 19122 27124
rect 21177 27115 21235 27121
rect 19116 27084 20208 27112
rect 19116 27072 19122 27084
rect 15562 27044 15568 27056
rect 15212 27016 15568 27044
rect 15562 27004 15568 27016
rect 15620 27004 15626 27056
rect 16298 27044 16304 27056
rect 15856 27016 16304 27044
rect 14875 26948 14964 26976
rect 15013 26979 15071 26985
rect 14875 26945 14887 26948
rect 14829 26939 14887 26945
rect 15013 26945 15025 26979
rect 15059 26976 15071 26979
rect 15102 26976 15108 26988
rect 15059 26948 15108 26976
rect 15059 26945 15071 26948
rect 15013 26939 15071 26945
rect 15102 26936 15108 26948
rect 15160 26936 15166 26988
rect 15746 26976 15752 26988
rect 15707 26948 15752 26976
rect 15746 26936 15752 26948
rect 15804 26936 15810 26988
rect 15856 26985 15884 27016
rect 16298 27004 16304 27016
rect 16356 27044 16362 27056
rect 17589 27047 17647 27053
rect 17589 27044 17601 27047
rect 16356 27016 17601 27044
rect 16356 27004 16362 27016
rect 17589 27013 17601 27016
rect 17635 27013 17647 27047
rect 17589 27007 17647 27013
rect 17954 27004 17960 27056
rect 18012 27044 18018 27056
rect 20180 27053 20208 27084
rect 21177 27081 21189 27115
rect 21223 27112 21235 27115
rect 21818 27112 21824 27124
rect 21223 27084 21824 27112
rect 21223 27081 21235 27084
rect 21177 27075 21235 27081
rect 21818 27072 21824 27084
rect 21876 27072 21882 27124
rect 23474 27112 23480 27124
rect 23435 27084 23480 27112
rect 23474 27072 23480 27084
rect 23532 27072 23538 27124
rect 25041 27115 25099 27121
rect 25041 27081 25053 27115
rect 25087 27112 25099 27115
rect 25314 27112 25320 27124
rect 25087 27084 25320 27112
rect 25087 27081 25099 27084
rect 25041 27075 25099 27081
rect 25314 27072 25320 27084
rect 25372 27072 25378 27124
rect 26326 27112 26332 27124
rect 26287 27084 26332 27112
rect 26326 27072 26332 27084
rect 26384 27072 26390 27124
rect 27522 27072 27528 27124
rect 27580 27072 27586 27124
rect 27617 27115 27675 27121
rect 27617 27081 27629 27115
rect 27663 27112 27675 27115
rect 27706 27112 27712 27124
rect 27663 27084 27712 27112
rect 27663 27081 27675 27084
rect 27617 27075 27675 27081
rect 27706 27072 27712 27084
rect 27764 27072 27770 27124
rect 28445 27115 28503 27121
rect 28445 27081 28457 27115
rect 28491 27081 28503 27115
rect 28445 27075 28503 27081
rect 18325 27047 18383 27053
rect 18325 27044 18337 27047
rect 18012 27016 18337 27044
rect 18012 27004 18018 27016
rect 18325 27013 18337 27016
rect 18371 27013 18383 27047
rect 18325 27007 18383 27013
rect 18509 27047 18567 27053
rect 18509 27013 18521 27047
rect 18555 27044 18567 27047
rect 20165 27047 20223 27053
rect 18555 27016 19472 27044
rect 18555 27013 18567 27016
rect 18509 27007 18567 27013
rect 15841 26979 15899 26985
rect 15841 26945 15853 26979
rect 15887 26945 15899 26979
rect 15841 26939 15899 26945
rect 15930 26936 15936 26988
rect 15988 26976 15994 26988
rect 15988 26948 16033 26976
rect 15988 26936 15994 26948
rect 16114 26936 16120 26988
rect 16172 26976 16178 26988
rect 16666 26976 16672 26988
rect 16172 26948 16217 26976
rect 16627 26948 16672 26976
rect 16172 26936 16178 26948
rect 16666 26936 16672 26948
rect 16724 26936 16730 26988
rect 16853 26979 16911 26985
rect 16853 26945 16865 26979
rect 16899 26945 16911 26979
rect 17494 26976 17500 26988
rect 17455 26948 17500 26976
rect 16853 26939 16911 26945
rect 15194 26868 15200 26920
rect 15252 26908 15258 26920
rect 16868 26908 16896 26939
rect 17494 26936 17500 26948
rect 17552 26936 17558 26988
rect 17681 26979 17739 26985
rect 17681 26945 17693 26979
rect 17727 26976 17739 26979
rect 18046 26976 18052 26988
rect 17727 26948 18052 26976
rect 17727 26945 17739 26948
rect 17681 26939 17739 26945
rect 18046 26936 18052 26948
rect 18104 26936 18110 26988
rect 18141 26979 18199 26985
rect 18141 26945 18153 26979
rect 18187 26945 18199 26979
rect 18141 26939 18199 26945
rect 15252 26880 16896 26908
rect 18156 26908 18184 26939
rect 18598 26936 18604 26988
rect 18656 26976 18662 26988
rect 19199 26979 19257 26985
rect 19199 26976 19211 26979
rect 18656 26948 19211 26976
rect 18656 26936 18662 26948
rect 19199 26945 19211 26948
rect 19245 26945 19257 26979
rect 19334 26976 19340 26988
rect 19295 26948 19340 26976
rect 19199 26939 19257 26945
rect 19334 26936 19340 26948
rect 19392 26936 19398 26988
rect 19444 26985 19472 27016
rect 20165 27013 20177 27047
rect 20211 27013 20223 27047
rect 20165 27007 20223 27013
rect 22554 27004 22560 27056
rect 22612 27044 22618 27056
rect 23293 27047 23351 27053
rect 23293 27044 23305 27047
rect 22612 27016 23305 27044
rect 22612 27004 22618 27016
rect 23293 27013 23305 27016
rect 23339 27044 23351 27047
rect 23750 27044 23756 27056
rect 23339 27016 23756 27044
rect 23339 27013 23351 27016
rect 23293 27007 23351 27013
rect 23750 27004 23756 27016
rect 23808 27004 23814 27056
rect 24673 27047 24731 27053
rect 24673 27013 24685 27047
rect 24719 27013 24731 27047
rect 26344 27044 26372 27072
rect 27540 27044 27568 27072
rect 28460 27044 28488 27075
rect 26344 27016 27384 27044
rect 27540 27016 28488 27044
rect 24673 27007 24731 27013
rect 19429 26979 19487 26985
rect 19429 26945 19441 26979
rect 19475 26945 19487 26979
rect 19429 26939 19487 26945
rect 19613 26979 19671 26985
rect 19613 26945 19625 26979
rect 19659 26976 19671 26979
rect 19978 26976 19984 26988
rect 19659 26948 19984 26976
rect 19659 26945 19671 26948
rect 19613 26939 19671 26945
rect 19978 26936 19984 26948
rect 20036 26936 20042 26988
rect 20346 26976 20352 26988
rect 20307 26948 20352 26976
rect 20346 26936 20352 26948
rect 20404 26936 20410 26988
rect 20993 26979 21051 26985
rect 20993 26945 21005 26979
rect 21039 26945 21051 26979
rect 20993 26939 21051 26945
rect 23109 26979 23167 26985
rect 23109 26945 23121 26979
rect 23155 26976 23167 26979
rect 23198 26976 23204 26988
rect 23155 26948 23204 26976
rect 23155 26945 23167 26948
rect 23109 26939 23167 26945
rect 21008 26908 21036 26939
rect 23198 26936 23204 26948
rect 23256 26976 23262 26988
rect 24688 26976 24716 27007
rect 27356 26988 27384 27016
rect 23256 26948 24716 26976
rect 23256 26936 23262 26948
rect 18156 26880 21036 26908
rect 24688 26908 24716 26948
rect 24857 26979 24915 26985
rect 24857 26945 24869 26979
rect 24903 26976 24915 26979
rect 25498 26976 25504 26988
rect 24903 26948 25504 26976
rect 24903 26945 24915 26948
rect 24857 26939 24915 26945
rect 25498 26936 25504 26948
rect 25556 26936 25562 26988
rect 26786 26936 26792 26988
rect 26844 26976 26850 26988
rect 26973 26979 27031 26985
rect 26973 26976 26985 26979
rect 26844 26948 26985 26976
rect 26844 26936 26850 26948
rect 26973 26945 26985 26948
rect 27019 26945 27031 26979
rect 27136 26979 27194 26985
rect 27136 26976 27148 26979
rect 26973 26939 27031 26945
rect 27080 26948 27148 26976
rect 26142 26908 26148 26920
rect 24688 26880 26148 26908
rect 15252 26868 15258 26880
rect 19260 26852 19288 26880
rect 26142 26868 26148 26880
rect 26200 26868 26206 26920
rect 27080 26852 27108 26948
rect 27136 26945 27148 26948
rect 27182 26945 27194 26979
rect 27136 26939 27194 26945
rect 27249 26979 27307 26985
rect 27249 26945 27261 26979
rect 27295 26945 27307 26979
rect 27249 26939 27307 26945
rect 27264 26908 27292 26939
rect 27338 26936 27344 26988
rect 27396 26976 27402 26988
rect 27396 26948 27489 26976
rect 27396 26936 27402 26948
rect 27522 26936 27528 26988
rect 27580 26976 27586 26988
rect 28077 26979 28135 26985
rect 28077 26976 28089 26979
rect 27580 26948 28089 26976
rect 27580 26936 27586 26948
rect 28077 26945 28089 26948
rect 28123 26945 28135 26979
rect 28077 26939 28135 26945
rect 28261 26979 28319 26985
rect 28261 26945 28273 26979
rect 28307 26976 28319 26979
rect 29178 26976 29184 26988
rect 28307 26948 29184 26976
rect 28307 26945 28319 26948
rect 28261 26939 28319 26945
rect 29178 26936 29184 26948
rect 29236 26936 29242 26988
rect 27430 26908 27436 26920
rect 27264 26880 27436 26908
rect 27430 26868 27436 26880
rect 27488 26868 27494 26920
rect 9732 26812 13400 26840
rect 13817 26843 13875 26849
rect 9732 26800 9738 26812
rect 13817 26809 13829 26843
rect 13863 26840 13875 26843
rect 16942 26840 16948 26852
rect 13863 26812 16948 26840
rect 13863 26809 13875 26812
rect 13817 26803 13875 26809
rect 16942 26800 16948 26812
rect 17000 26800 17006 26852
rect 19242 26800 19248 26852
rect 19300 26800 19306 26852
rect 20533 26843 20591 26849
rect 20533 26809 20545 26843
rect 20579 26840 20591 26843
rect 22002 26840 22008 26852
rect 20579 26812 22008 26840
rect 20579 26809 20591 26812
rect 20533 26803 20591 26809
rect 22002 26800 22008 26812
rect 22060 26800 22066 26852
rect 23566 26800 23572 26852
rect 23624 26840 23630 26852
rect 26326 26840 26332 26852
rect 23624 26812 26332 26840
rect 23624 26800 23630 26812
rect 26326 26800 26332 26812
rect 26384 26800 26390 26852
rect 27062 26800 27068 26852
rect 27120 26800 27126 26852
rect 8202 26772 8208 26784
rect 7576 26744 8208 26772
rect 8202 26732 8208 26744
rect 8260 26732 8266 26784
rect 13906 26732 13912 26784
rect 13964 26772 13970 26784
rect 15470 26772 15476 26784
rect 13964 26744 15476 26772
rect 13964 26732 13970 26744
rect 15470 26732 15476 26744
rect 15528 26732 15534 26784
rect 15654 26732 15660 26784
rect 15712 26772 15718 26784
rect 17037 26775 17095 26781
rect 17037 26772 17049 26775
rect 15712 26744 17049 26772
rect 15712 26732 15718 26744
rect 17037 26741 17049 26744
rect 17083 26741 17095 26775
rect 17037 26735 17095 26741
rect 17402 26732 17408 26784
rect 17460 26772 17466 26784
rect 18414 26772 18420 26784
rect 17460 26744 18420 26772
rect 17460 26732 17466 26744
rect 18414 26732 18420 26744
rect 18472 26732 18478 26784
rect 67634 26772 67640 26784
rect 67595 26744 67640 26772
rect 67634 26732 67640 26744
rect 67692 26732 67698 26784
rect 1104 26682 68816 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 65654 26682
rect 65706 26630 65718 26682
rect 65770 26630 65782 26682
rect 65834 26630 65846 26682
rect 65898 26630 65910 26682
rect 65962 26630 68816 26682
rect 1104 26608 68816 26630
rect 5810 26568 5816 26580
rect 5723 26540 5816 26568
rect 5810 26528 5816 26540
rect 5868 26568 5874 26580
rect 9674 26568 9680 26580
rect 5868 26540 9680 26568
rect 5868 26528 5874 26540
rect 9674 26528 9680 26540
rect 9732 26528 9738 26580
rect 14090 26528 14096 26580
rect 14148 26568 14154 26580
rect 15194 26568 15200 26580
rect 14148 26540 15200 26568
rect 14148 26528 14154 26540
rect 15194 26528 15200 26540
rect 15252 26528 15258 26580
rect 15470 26528 15476 26580
rect 15528 26568 15534 26580
rect 16114 26568 16120 26580
rect 15528 26540 16120 26568
rect 15528 26528 15534 26540
rect 16114 26528 16120 26540
rect 16172 26528 16178 26580
rect 26881 26571 26939 26577
rect 26881 26537 26893 26571
rect 26927 26568 26939 26571
rect 27062 26568 27068 26580
rect 26927 26540 27068 26568
rect 26927 26537 26939 26540
rect 26881 26531 26939 26537
rect 27062 26528 27068 26540
rect 27120 26528 27126 26580
rect 14645 26503 14703 26509
rect 14645 26469 14657 26503
rect 14691 26469 14703 26503
rect 14645 26463 14703 26469
rect 2590 26432 2596 26444
rect 2551 26404 2596 26432
rect 2590 26392 2596 26404
rect 2648 26392 2654 26444
rect 7006 26432 7012 26444
rect 6967 26404 7012 26432
rect 7006 26392 7012 26404
rect 7064 26392 7070 26444
rect 7466 26392 7472 26444
rect 7524 26432 7530 26444
rect 9214 26432 9220 26444
rect 7524 26404 9220 26432
rect 7524 26392 7530 26404
rect 9214 26392 9220 26404
rect 9272 26392 9278 26444
rect 13722 26392 13728 26444
rect 13780 26432 13786 26444
rect 14660 26432 14688 26463
rect 14918 26460 14924 26512
rect 14976 26500 14982 26512
rect 16666 26500 16672 26512
rect 14976 26472 16672 26500
rect 14976 26460 14982 26472
rect 16666 26460 16672 26472
rect 16724 26460 16730 26512
rect 17402 26500 17408 26512
rect 17363 26472 17408 26500
rect 17402 26460 17408 26472
rect 17460 26460 17466 26512
rect 20346 26500 20352 26512
rect 19260 26472 20352 26500
rect 19260 26432 19288 26472
rect 20346 26460 20352 26472
rect 20404 26500 20410 26512
rect 21361 26503 21419 26509
rect 21361 26500 21373 26503
rect 20404 26472 21373 26500
rect 20404 26460 20410 26472
rect 21361 26469 21373 26472
rect 21407 26469 21419 26503
rect 21361 26463 21419 26469
rect 13780 26404 14504 26432
rect 14660 26404 16804 26432
rect 13780 26392 13786 26404
rect 2869 26367 2927 26373
rect 2869 26333 2881 26367
rect 2915 26364 2927 26367
rect 3878 26364 3884 26376
rect 2915 26336 3884 26364
rect 2915 26333 2927 26336
rect 2869 26327 2927 26333
rect 3878 26324 3884 26336
rect 3936 26324 3942 26376
rect 4246 26324 4252 26376
rect 4304 26364 4310 26376
rect 4433 26367 4491 26373
rect 4433 26364 4445 26367
rect 4304 26336 4445 26364
rect 4304 26324 4310 26336
rect 4433 26333 4445 26336
rect 4479 26364 4491 26367
rect 5442 26364 5448 26376
rect 4479 26336 5448 26364
rect 4479 26333 4491 26336
rect 4433 26327 4491 26333
rect 5442 26324 5448 26336
rect 5500 26324 5506 26376
rect 7282 26364 7288 26376
rect 7243 26336 7288 26364
rect 7282 26324 7288 26336
rect 7340 26324 7346 26376
rect 7926 26364 7932 26376
rect 7839 26336 7932 26364
rect 7926 26324 7932 26336
rect 7984 26364 7990 26376
rect 8113 26367 8171 26373
rect 7984 26336 8064 26364
rect 7984 26324 7990 26336
rect 3050 26256 3056 26308
rect 3108 26296 3114 26308
rect 4678 26299 4736 26305
rect 4678 26296 4690 26299
rect 3108 26268 4690 26296
rect 3108 26256 3114 26268
rect 4678 26265 4690 26268
rect 4724 26265 4736 26299
rect 8036 26296 8064 26336
rect 8113 26333 8125 26367
rect 8159 26364 8171 26367
rect 8846 26364 8852 26376
rect 8159 26336 8852 26364
rect 8159 26333 8171 26336
rect 8113 26327 8171 26333
rect 8846 26324 8852 26336
rect 8904 26324 8910 26376
rect 11790 26364 11796 26376
rect 11703 26336 11796 26364
rect 11790 26324 11796 26336
rect 11848 26364 11854 26376
rect 13814 26364 13820 26376
rect 11848 26336 13820 26364
rect 11848 26324 11854 26336
rect 13814 26324 13820 26336
rect 13872 26324 13878 26376
rect 14090 26364 14096 26376
rect 14051 26336 14096 26364
rect 14090 26324 14096 26336
rect 14148 26324 14154 26376
rect 14476 26373 14504 26404
rect 14461 26367 14519 26373
rect 14461 26333 14473 26367
rect 14507 26333 14519 26367
rect 14461 26327 14519 26333
rect 14734 26324 14740 26376
rect 14792 26364 14798 26376
rect 15102 26364 15108 26376
rect 14792 26336 15108 26364
rect 14792 26324 14798 26336
rect 15102 26324 15108 26336
rect 15160 26324 15166 26376
rect 15378 26324 15384 26376
rect 15436 26364 15442 26376
rect 15473 26367 15531 26373
rect 15473 26364 15485 26367
rect 15436 26336 15485 26364
rect 15436 26324 15442 26336
rect 15473 26333 15485 26336
rect 15519 26333 15531 26367
rect 15473 26327 15531 26333
rect 15565 26367 15623 26373
rect 15565 26333 15577 26367
rect 15611 26333 15623 26367
rect 15565 26327 15623 26333
rect 8036 26268 8156 26296
rect 4678 26259 4736 26265
rect 7466 26188 7472 26240
rect 7524 26228 7530 26240
rect 7745 26231 7803 26237
rect 7745 26228 7757 26231
rect 7524 26200 7757 26228
rect 7524 26188 7530 26200
rect 7745 26197 7757 26200
rect 7791 26197 7803 26231
rect 8128 26228 8156 26268
rect 8386 26256 8392 26308
rect 8444 26296 8450 26308
rect 8941 26299 8999 26305
rect 8941 26296 8953 26299
rect 8444 26268 8953 26296
rect 8444 26256 8450 26268
rect 8941 26265 8953 26268
rect 8987 26296 8999 26299
rect 9306 26296 9312 26308
rect 8987 26268 9312 26296
rect 8987 26265 8999 26268
rect 8941 26259 8999 26265
rect 9306 26256 9312 26268
rect 9364 26256 9370 26308
rect 11548 26299 11606 26305
rect 11548 26265 11560 26299
rect 11594 26296 11606 26299
rect 12894 26296 12900 26308
rect 11594 26268 12900 26296
rect 11594 26265 11606 26268
rect 11548 26259 11606 26265
rect 12894 26256 12900 26268
rect 12952 26256 12958 26308
rect 12986 26256 12992 26308
rect 13044 26296 13050 26308
rect 14274 26296 14280 26308
rect 13044 26268 13860 26296
rect 14235 26268 14280 26296
rect 13044 26256 13050 26268
rect 13832 26240 13860 26268
rect 14274 26256 14280 26268
rect 14332 26256 14338 26308
rect 14366 26256 14372 26308
rect 14424 26296 14430 26308
rect 14424 26268 14469 26296
rect 14424 26256 14430 26268
rect 15010 26256 15016 26308
rect 15068 26296 15074 26308
rect 15580 26296 15608 26327
rect 15654 26324 15660 26376
rect 15712 26364 15718 26376
rect 16776 26373 16804 26404
rect 16960 26404 19288 26432
rect 16960 26373 16988 26404
rect 19334 26392 19340 26444
rect 19392 26432 19398 26444
rect 19981 26435 20039 26441
rect 19981 26432 19993 26435
rect 19392 26404 19993 26432
rect 19392 26392 19398 26404
rect 19981 26401 19993 26404
rect 20027 26401 20039 26435
rect 19981 26395 20039 26401
rect 30282 26392 30288 26444
rect 30340 26432 30346 26444
rect 30377 26435 30435 26441
rect 30377 26432 30389 26435
rect 30340 26404 30389 26432
rect 30340 26392 30346 26404
rect 30377 26401 30389 26404
rect 30423 26401 30435 26435
rect 30377 26395 30435 26401
rect 15841 26367 15899 26373
rect 15712 26336 15757 26364
rect 15712 26324 15718 26336
rect 15841 26333 15853 26367
rect 15887 26333 15899 26367
rect 15841 26327 15899 26333
rect 16761 26367 16819 26373
rect 16761 26333 16773 26367
rect 16807 26333 16819 26367
rect 16761 26327 16819 26333
rect 16909 26367 16988 26373
rect 16909 26333 16921 26367
rect 16955 26336 16988 26367
rect 16955 26333 16967 26336
rect 16909 26327 16967 26333
rect 15856 26296 15884 26327
rect 17034 26324 17040 26376
rect 17092 26364 17098 26376
rect 17092 26336 17137 26364
rect 17092 26324 17098 26336
rect 17218 26324 17224 26376
rect 17276 26373 17282 26376
rect 17276 26364 17284 26373
rect 17770 26364 17776 26376
rect 17276 26336 17321 26364
rect 17420 26336 17776 26364
rect 17276 26327 17284 26336
rect 17276 26324 17282 26327
rect 15068 26268 15608 26296
rect 15672 26268 15884 26296
rect 15068 26256 15074 26268
rect 8478 26228 8484 26240
rect 8128 26200 8484 26228
rect 7745 26191 7803 26197
rect 8478 26188 8484 26200
rect 8536 26188 8542 26240
rect 10410 26228 10416 26240
rect 10371 26200 10416 26228
rect 10410 26188 10416 26200
rect 10468 26188 10474 26240
rect 13814 26228 13820 26240
rect 13727 26200 13820 26228
rect 13814 26188 13820 26200
rect 13872 26228 13878 26240
rect 14734 26228 14740 26240
rect 13872 26200 14740 26228
rect 13872 26188 13878 26200
rect 14734 26188 14740 26200
rect 14792 26228 14798 26240
rect 14918 26228 14924 26240
rect 14792 26200 14924 26228
rect 14792 26188 14798 26200
rect 14918 26188 14924 26200
rect 14976 26188 14982 26240
rect 15194 26228 15200 26240
rect 15155 26200 15200 26228
rect 15194 26188 15200 26200
rect 15252 26188 15258 26240
rect 15286 26188 15292 26240
rect 15344 26228 15350 26240
rect 15672 26228 15700 26268
rect 17126 26256 17132 26308
rect 17184 26296 17190 26308
rect 17184 26268 17229 26296
rect 17184 26256 17190 26268
rect 15344 26200 15700 26228
rect 15344 26188 15350 26200
rect 16666 26188 16672 26240
rect 16724 26228 16730 26240
rect 17420 26228 17448 26336
rect 17770 26324 17776 26336
rect 17828 26364 17834 26376
rect 17865 26367 17923 26373
rect 17865 26364 17877 26367
rect 17828 26336 17877 26364
rect 17828 26324 17834 26336
rect 17865 26333 17877 26336
rect 17911 26333 17923 26367
rect 18138 26364 18144 26376
rect 18099 26336 18144 26364
rect 17865 26327 17923 26333
rect 18138 26324 18144 26336
rect 18196 26324 18202 26376
rect 19242 26324 19248 26376
rect 19300 26364 19306 26376
rect 19429 26367 19487 26373
rect 19429 26364 19441 26367
rect 19300 26336 19441 26364
rect 19300 26324 19306 26336
rect 19429 26333 19441 26336
rect 19475 26333 19487 26367
rect 19429 26327 19487 26333
rect 20257 26367 20315 26373
rect 20257 26333 20269 26367
rect 20303 26364 20315 26367
rect 20346 26364 20352 26376
rect 20303 26336 20352 26364
rect 20303 26333 20315 26336
rect 20257 26327 20315 26333
rect 20346 26324 20352 26336
rect 20404 26324 20410 26376
rect 22738 26364 22744 26376
rect 22699 26336 22744 26364
rect 22738 26324 22744 26336
rect 22796 26364 22802 26376
rect 26053 26367 26111 26373
rect 26053 26364 26065 26367
rect 22796 26336 26065 26364
rect 22796 26324 22802 26336
rect 26053 26333 26065 26336
rect 26099 26364 26111 26367
rect 26234 26364 26240 26376
rect 26099 26336 26240 26364
rect 26099 26333 26111 26336
rect 26053 26327 26111 26333
rect 26234 26324 26240 26336
rect 26292 26324 26298 26376
rect 26697 26367 26755 26373
rect 26697 26364 26709 26367
rect 26436 26336 26709 26364
rect 22462 26296 22468 26308
rect 22520 26305 22526 26308
rect 22432 26268 22468 26296
rect 22462 26256 22468 26268
rect 22520 26259 22532 26305
rect 22520 26256 22526 26259
rect 23198 26256 23204 26308
rect 23256 26296 23262 26308
rect 23477 26299 23535 26305
rect 23477 26296 23489 26299
rect 23256 26268 23489 26296
rect 23256 26256 23262 26268
rect 23477 26265 23489 26268
rect 23523 26265 23535 26299
rect 23477 26259 23535 26265
rect 23566 26256 23572 26308
rect 23624 26296 23630 26308
rect 23661 26299 23719 26305
rect 23661 26296 23673 26299
rect 23624 26268 23673 26296
rect 23624 26256 23630 26268
rect 23661 26265 23673 26268
rect 23707 26296 23719 26299
rect 23707 26268 24716 26296
rect 23707 26265 23719 26268
rect 23661 26259 23719 26265
rect 16724 26200 17448 26228
rect 16724 26188 16730 26200
rect 18690 26188 18696 26240
rect 18748 26228 18754 26240
rect 19058 26228 19064 26240
rect 18748 26200 19064 26228
rect 18748 26188 18754 26200
rect 19058 26188 19064 26200
rect 19116 26228 19122 26240
rect 19245 26231 19303 26237
rect 19245 26228 19257 26231
rect 19116 26200 19257 26228
rect 19116 26188 19122 26200
rect 19245 26197 19257 26200
rect 19291 26197 19303 26231
rect 23842 26228 23848 26240
rect 23803 26200 23848 26228
rect 19245 26191 19303 26197
rect 23842 26188 23848 26200
rect 23900 26188 23906 26240
rect 24688 26237 24716 26268
rect 24854 26256 24860 26308
rect 24912 26296 24918 26308
rect 25786 26299 25844 26305
rect 25786 26296 25798 26299
rect 24912 26268 25798 26296
rect 24912 26256 24918 26268
rect 25786 26265 25798 26268
rect 25832 26265 25844 26299
rect 25786 26259 25844 26265
rect 25958 26256 25964 26308
rect 26016 26296 26022 26308
rect 26436 26296 26464 26336
rect 26697 26333 26709 26336
rect 26743 26364 26755 26367
rect 27614 26364 27620 26376
rect 26743 26336 27620 26364
rect 26743 26333 26755 26336
rect 26697 26327 26755 26333
rect 27614 26324 27620 26336
rect 27672 26324 27678 26376
rect 26016 26268 26464 26296
rect 26513 26299 26571 26305
rect 26016 26256 26022 26268
rect 26513 26265 26525 26299
rect 26559 26296 26571 26299
rect 26970 26296 26976 26308
rect 26559 26268 26976 26296
rect 26559 26265 26571 26268
rect 26513 26259 26571 26265
rect 26970 26256 26976 26268
rect 27028 26296 27034 26308
rect 27522 26296 27528 26308
rect 27028 26268 27528 26296
rect 27028 26256 27034 26268
rect 27522 26256 27528 26268
rect 27580 26256 27586 26308
rect 30644 26299 30702 26305
rect 30644 26265 30656 26299
rect 30690 26296 30702 26299
rect 30742 26296 30748 26308
rect 30690 26268 30748 26296
rect 30690 26265 30702 26268
rect 30644 26259 30702 26265
rect 30742 26256 30748 26268
rect 30800 26256 30806 26308
rect 24673 26231 24731 26237
rect 24673 26197 24685 26231
rect 24719 26197 24731 26231
rect 24673 26191 24731 26197
rect 31570 26188 31576 26240
rect 31628 26228 31634 26240
rect 31757 26231 31815 26237
rect 31757 26228 31769 26231
rect 31628 26200 31769 26228
rect 31628 26188 31634 26200
rect 31757 26197 31769 26200
rect 31803 26197 31815 26231
rect 31757 26191 31815 26197
rect 1104 26138 68816 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 68816 26138
rect 1104 26064 68816 26086
rect 13173 26027 13231 26033
rect 13173 25993 13185 26027
rect 13219 26024 13231 26027
rect 14090 26024 14096 26036
rect 13219 25996 14096 26024
rect 13219 25993 13231 25996
rect 13173 25987 13231 25993
rect 14090 25984 14096 25996
rect 14148 25984 14154 26036
rect 14458 25984 14464 26036
rect 14516 26024 14522 26036
rect 18141 26027 18199 26033
rect 18141 26024 18153 26027
rect 14516 25996 18153 26024
rect 14516 25984 14522 25996
rect 18141 25993 18153 25996
rect 18187 25993 18199 26027
rect 18141 25987 18199 25993
rect 2041 25959 2099 25965
rect 2041 25925 2053 25959
rect 2087 25956 2099 25959
rect 5810 25956 5816 25968
rect 2087 25928 5816 25956
rect 2087 25925 2099 25928
rect 2041 25919 2099 25925
rect 5810 25916 5816 25928
rect 5868 25916 5874 25968
rect 6733 25959 6791 25965
rect 6733 25925 6745 25959
rect 6779 25956 6791 25959
rect 8386 25956 8392 25968
rect 6779 25928 8392 25956
rect 6779 25925 6791 25928
rect 6733 25919 6791 25925
rect 8386 25916 8392 25928
rect 8444 25916 8450 25968
rect 9398 25956 9404 25968
rect 8956 25928 9404 25956
rect 1670 25848 1676 25900
rect 1728 25888 1734 25900
rect 1857 25891 1915 25897
rect 1857 25888 1869 25891
rect 1728 25860 1869 25888
rect 1728 25848 1734 25860
rect 1857 25857 1869 25860
rect 1903 25857 1915 25891
rect 1857 25851 1915 25857
rect 2958 25848 2964 25900
rect 3016 25888 3022 25900
rect 3982 25891 4040 25897
rect 3982 25888 3994 25891
rect 3016 25860 3994 25888
rect 3016 25848 3022 25860
rect 3982 25857 3994 25860
rect 4028 25857 4040 25891
rect 4246 25888 4252 25900
rect 4207 25860 4252 25888
rect 3982 25851 4040 25857
rect 4246 25848 4252 25860
rect 4304 25848 4310 25900
rect 8294 25848 8300 25900
rect 8352 25888 8358 25900
rect 8956 25897 8984 25928
rect 9398 25916 9404 25928
rect 9456 25916 9462 25968
rect 12060 25959 12118 25965
rect 12060 25925 12072 25959
rect 12106 25956 12118 25959
rect 15194 25956 15200 25968
rect 12106 25928 15200 25956
rect 12106 25925 12118 25928
rect 12060 25919 12118 25925
rect 15194 25916 15200 25928
rect 15252 25916 15258 25968
rect 18156 25956 18184 25987
rect 20622 25984 20628 26036
rect 20680 26024 20686 26036
rect 20809 26027 20867 26033
rect 20809 26024 20821 26027
rect 20680 25996 20821 26024
rect 20680 25984 20686 25996
rect 20809 25993 20821 25996
rect 20855 25993 20867 26027
rect 22462 26024 22468 26036
rect 22423 25996 22468 26024
rect 20809 25987 20867 25993
rect 22462 25984 22468 25996
rect 22520 25984 22526 26036
rect 24854 26024 24860 26036
rect 24815 25996 24860 26024
rect 24854 25984 24860 25996
rect 24912 25984 24918 26036
rect 26050 25984 26056 26036
rect 26108 26024 26114 26036
rect 26329 26027 26387 26033
rect 26329 26024 26341 26027
rect 26108 25996 26341 26024
rect 26108 25984 26114 25996
rect 26329 25993 26341 25996
rect 26375 26024 26387 26027
rect 26375 25996 27287 26024
rect 26375 25993 26387 25996
rect 26329 25987 26387 25993
rect 19521 25959 19579 25965
rect 19521 25956 19533 25959
rect 18156 25928 19533 25956
rect 19521 25925 19533 25928
rect 19567 25925 19579 25959
rect 19521 25919 19579 25925
rect 20346 25916 20352 25968
rect 20404 25956 20410 25968
rect 20404 25928 22140 25956
rect 20404 25916 20410 25928
rect 8481 25891 8539 25897
rect 8481 25888 8493 25891
rect 8352 25860 8493 25888
rect 8352 25848 8358 25860
rect 8481 25857 8493 25860
rect 8527 25888 8539 25891
rect 8941 25891 8999 25897
rect 8941 25888 8953 25891
rect 8527 25860 8953 25888
rect 8527 25857 8539 25860
rect 8481 25851 8539 25857
rect 8941 25857 8953 25860
rect 8987 25857 8999 25891
rect 8941 25851 8999 25857
rect 9030 25848 9036 25900
rect 9088 25888 9094 25900
rect 9197 25891 9255 25897
rect 9197 25888 9209 25891
rect 9088 25860 9209 25888
rect 9088 25848 9094 25860
rect 9197 25857 9209 25860
rect 9243 25857 9255 25891
rect 11790 25888 11796 25900
rect 11751 25860 11796 25888
rect 9197 25851 9255 25857
rect 11790 25848 11796 25860
rect 11848 25848 11854 25900
rect 14642 25888 14648 25900
rect 14603 25860 14648 25888
rect 14642 25848 14648 25860
rect 14700 25848 14706 25900
rect 15562 25888 15568 25900
rect 15523 25860 15568 25888
rect 15562 25848 15568 25860
rect 15620 25848 15626 25900
rect 16945 25891 17003 25897
rect 16945 25857 16957 25891
rect 16991 25888 17003 25891
rect 17034 25888 17040 25900
rect 16991 25860 17040 25888
rect 16991 25857 17003 25860
rect 16945 25851 17003 25857
rect 17034 25848 17040 25860
rect 17092 25888 17098 25900
rect 17310 25888 17316 25900
rect 17092 25860 17316 25888
rect 17092 25848 17098 25860
rect 17310 25848 17316 25860
rect 17368 25848 17374 25900
rect 18138 25848 18144 25900
rect 18196 25888 18202 25900
rect 18690 25888 18696 25900
rect 18196 25860 18696 25888
rect 18196 25848 18202 25860
rect 18690 25848 18696 25860
rect 18748 25848 18754 25900
rect 18874 25888 18880 25900
rect 18835 25860 18880 25888
rect 18874 25848 18880 25860
rect 18932 25848 18938 25900
rect 20530 25848 20536 25900
rect 20588 25888 20594 25900
rect 21821 25891 21879 25897
rect 21821 25888 21833 25891
rect 20588 25860 21833 25888
rect 20588 25848 20594 25860
rect 21821 25857 21833 25860
rect 21867 25857 21879 25891
rect 22002 25888 22008 25900
rect 21963 25860 22008 25888
rect 21821 25851 21879 25857
rect 22002 25848 22008 25860
rect 22060 25848 22066 25900
rect 22112 25897 22140 25928
rect 23842 25916 23848 25968
rect 23900 25956 23906 25968
rect 27259 25956 27287 25996
rect 30282 25984 30288 26036
rect 30340 25984 30346 26036
rect 30742 26024 30748 26036
rect 30703 25996 30748 26024
rect 30742 25984 30748 25996
rect 30800 25984 30806 26036
rect 27709 25959 27767 25965
rect 23900 25928 24348 25956
rect 27259 25928 27476 25956
rect 23900 25916 23906 25928
rect 22097 25891 22155 25897
rect 22097 25857 22109 25891
rect 22143 25857 22155 25891
rect 22097 25851 22155 25857
rect 22186 25848 22192 25900
rect 22244 25888 22250 25900
rect 22925 25891 22983 25897
rect 22925 25888 22937 25891
rect 22244 25860 22937 25888
rect 22244 25848 22250 25860
rect 22925 25857 22937 25860
rect 22971 25857 22983 25891
rect 24210 25888 24216 25900
rect 24171 25860 24216 25888
rect 22925 25851 22983 25857
rect 24210 25848 24216 25860
rect 24268 25848 24274 25900
rect 24320 25888 24348 25928
rect 24376 25891 24434 25897
rect 24376 25888 24388 25891
rect 24320 25860 24388 25888
rect 24376 25857 24388 25860
rect 24422 25857 24434 25891
rect 24376 25851 24434 25857
rect 24492 25891 24550 25897
rect 24492 25857 24504 25891
rect 24538 25857 24550 25891
rect 24492 25851 24550 25857
rect 14090 25780 14096 25832
rect 14148 25820 14154 25832
rect 14918 25820 14924 25832
rect 14148 25792 14924 25820
rect 14148 25780 14154 25792
rect 14918 25780 14924 25792
rect 14976 25820 14982 25832
rect 15289 25823 15347 25829
rect 15289 25820 15301 25823
rect 14976 25792 15301 25820
rect 14976 25780 14982 25792
rect 15289 25789 15301 25792
rect 15335 25789 15347 25823
rect 16666 25820 16672 25832
rect 16627 25792 16672 25820
rect 15289 25783 15347 25789
rect 16666 25780 16672 25792
rect 16724 25780 16730 25832
rect 23750 25780 23756 25832
rect 23808 25820 23814 25832
rect 24507 25820 24535 25851
rect 24578 25848 24584 25900
rect 24636 25897 24642 25900
rect 24636 25891 24659 25897
rect 24647 25857 24659 25891
rect 24636 25851 24659 25857
rect 24636 25848 24642 25851
rect 25406 25848 25412 25900
rect 25464 25888 25470 25900
rect 26786 25888 26792 25900
rect 25464 25860 26792 25888
rect 25464 25848 25470 25860
rect 26786 25848 26792 25860
rect 26844 25888 26850 25900
rect 27065 25891 27123 25897
rect 27065 25888 27077 25891
rect 26844 25860 27077 25888
rect 26844 25848 26850 25860
rect 27065 25857 27077 25860
rect 27111 25857 27123 25891
rect 27246 25888 27252 25900
rect 27207 25860 27252 25888
rect 27065 25851 27123 25857
rect 27246 25848 27252 25860
rect 27304 25848 27310 25900
rect 27448 25897 27476 25928
rect 27709 25925 27721 25959
rect 27755 25956 27767 25959
rect 29282 25959 29340 25965
rect 29282 25956 29294 25959
rect 27755 25928 29294 25956
rect 27755 25925 27767 25928
rect 27709 25919 27767 25925
rect 29282 25925 29294 25928
rect 29328 25925 29340 25959
rect 30300 25956 30328 25984
rect 29282 25919 29340 25925
rect 29564 25928 30328 25956
rect 31389 25959 31447 25965
rect 27341 25891 27399 25897
rect 27341 25857 27353 25891
rect 27387 25857 27399 25891
rect 27341 25851 27399 25857
rect 27433 25891 27491 25897
rect 27433 25857 27445 25891
rect 27479 25888 27491 25891
rect 27522 25888 27528 25900
rect 27479 25860 27528 25888
rect 27479 25857 27491 25860
rect 27433 25851 27491 25857
rect 24946 25820 24952 25832
rect 23808 25792 24952 25820
rect 23808 25780 23814 25792
rect 24946 25780 24952 25792
rect 25004 25780 25010 25832
rect 27356 25820 27384 25851
rect 27522 25848 27528 25860
rect 27580 25848 27586 25900
rect 29564 25897 29592 25928
rect 31389 25925 31401 25959
rect 31435 25956 31447 25959
rect 31570 25956 31576 25968
rect 31435 25928 31576 25956
rect 31435 25925 31447 25928
rect 31389 25919 31447 25925
rect 31570 25916 31576 25928
rect 31628 25916 31634 25968
rect 29549 25891 29607 25897
rect 29549 25857 29561 25891
rect 29595 25857 29607 25891
rect 30098 25888 30104 25900
rect 30059 25860 30104 25888
rect 29549 25851 29607 25857
rect 30098 25848 30104 25860
rect 30156 25848 30162 25900
rect 30282 25888 30288 25900
rect 30243 25860 30288 25888
rect 30282 25848 30288 25860
rect 30340 25848 30346 25900
rect 30558 25897 30564 25900
rect 30380 25891 30438 25897
rect 30380 25857 30392 25891
rect 30426 25857 30438 25891
rect 30380 25851 30438 25857
rect 30515 25891 30564 25897
rect 30515 25857 30527 25891
rect 30561 25857 30564 25891
rect 30515 25851 30564 25857
rect 27356 25792 27476 25820
rect 27448 25764 27476 25792
rect 17126 25752 17132 25764
rect 13096 25724 17132 25752
rect 2225 25687 2283 25693
rect 2225 25653 2237 25687
rect 2271 25684 2283 25687
rect 2406 25684 2412 25696
rect 2271 25656 2412 25684
rect 2271 25653 2283 25656
rect 2225 25647 2283 25653
rect 2406 25644 2412 25656
rect 2464 25644 2470 25696
rect 2866 25684 2872 25696
rect 2827 25656 2872 25684
rect 2866 25644 2872 25656
rect 2924 25644 2930 25696
rect 9122 25644 9128 25696
rect 9180 25684 9186 25696
rect 10321 25687 10379 25693
rect 10321 25684 10333 25687
rect 9180 25656 10333 25684
rect 9180 25644 9186 25656
rect 10321 25653 10333 25656
rect 10367 25684 10379 25687
rect 13096 25684 13124 25724
rect 17126 25712 17132 25724
rect 17184 25712 17190 25764
rect 27430 25712 27436 25764
rect 27488 25712 27494 25764
rect 29822 25712 29828 25764
rect 29880 25752 29886 25764
rect 30395 25752 30423 25851
rect 30558 25848 30564 25851
rect 30616 25848 30622 25900
rect 31018 25848 31024 25900
rect 31076 25888 31082 25900
rect 31205 25891 31263 25897
rect 31205 25888 31217 25891
rect 31076 25860 31217 25888
rect 31076 25848 31082 25860
rect 31205 25857 31217 25860
rect 31251 25857 31263 25891
rect 31205 25851 31263 25857
rect 29880 25724 30423 25752
rect 29880 25712 29886 25724
rect 10367 25656 13124 25684
rect 10367 25653 10379 25656
rect 10321 25647 10379 25653
rect 13170 25644 13176 25696
rect 13228 25684 13234 25696
rect 13633 25687 13691 25693
rect 13633 25684 13645 25687
rect 13228 25656 13645 25684
rect 13228 25644 13234 25656
rect 13633 25653 13645 25656
rect 13679 25653 13691 25687
rect 13633 25647 13691 25653
rect 14734 25644 14740 25696
rect 14792 25684 14798 25696
rect 14829 25687 14887 25693
rect 14829 25684 14841 25687
rect 14792 25656 14841 25684
rect 14792 25644 14798 25656
rect 14829 25653 14841 25656
rect 14875 25653 14887 25687
rect 14829 25647 14887 25653
rect 19061 25687 19119 25693
rect 19061 25653 19073 25687
rect 19107 25684 19119 25687
rect 19702 25684 19708 25696
rect 19107 25656 19708 25684
rect 19107 25653 19119 25656
rect 19061 25647 19119 25653
rect 19702 25644 19708 25656
rect 19760 25644 19766 25696
rect 21726 25644 21732 25696
rect 21784 25684 21790 25696
rect 23658 25684 23664 25696
rect 21784 25656 23664 25684
rect 21784 25644 21790 25656
rect 23658 25644 23664 25656
rect 23716 25684 23722 25696
rect 24578 25684 24584 25696
rect 23716 25656 24584 25684
rect 23716 25644 23722 25656
rect 24578 25644 24584 25656
rect 24636 25684 24642 25696
rect 26878 25684 26884 25696
rect 24636 25656 26884 25684
rect 24636 25644 24642 25656
rect 26878 25644 26884 25656
rect 26936 25644 26942 25696
rect 27154 25644 27160 25696
rect 27212 25684 27218 25696
rect 28169 25687 28227 25693
rect 28169 25684 28181 25687
rect 27212 25656 28181 25684
rect 27212 25644 27218 25656
rect 28169 25653 28181 25656
rect 28215 25653 28227 25687
rect 28169 25647 28227 25653
rect 30282 25644 30288 25696
rect 30340 25684 30346 25696
rect 31573 25687 31631 25693
rect 31573 25684 31585 25687
rect 30340 25656 31585 25684
rect 30340 25644 30346 25656
rect 31573 25653 31585 25656
rect 31619 25653 31631 25687
rect 31573 25647 31631 25653
rect 1104 25594 68816 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 65654 25594
rect 65706 25542 65718 25594
rect 65770 25542 65782 25594
rect 65834 25542 65846 25594
rect 65898 25542 65910 25594
rect 65962 25542 68816 25594
rect 1104 25520 68816 25542
rect 2958 25480 2964 25492
rect 2919 25452 2964 25480
rect 2958 25440 2964 25452
rect 3016 25440 3022 25492
rect 6733 25483 6791 25489
rect 5368 25452 6316 25480
rect 2866 25412 2872 25424
rect 1688 25384 2872 25412
rect 1688 25285 1716 25384
rect 2866 25372 2872 25384
rect 2924 25412 2930 25424
rect 5368 25412 5396 25452
rect 2924 25384 5396 25412
rect 6288 25412 6316 25452
rect 6733 25449 6745 25483
rect 6779 25480 6791 25483
rect 7926 25480 7932 25492
rect 6779 25452 7932 25480
rect 6779 25449 6791 25452
rect 6733 25443 6791 25449
rect 7926 25440 7932 25452
rect 7984 25440 7990 25492
rect 8389 25483 8447 25489
rect 8389 25449 8401 25483
rect 8435 25480 8447 25483
rect 9030 25480 9036 25492
rect 8435 25452 9036 25480
rect 8435 25449 8447 25452
rect 8389 25443 8447 25449
rect 9030 25440 9036 25452
rect 9088 25440 9094 25492
rect 12894 25480 12900 25492
rect 12855 25452 12900 25480
rect 12894 25440 12900 25452
rect 12952 25440 12958 25492
rect 18874 25480 18880 25492
rect 17144 25452 18880 25480
rect 14366 25412 14372 25424
rect 6288 25384 14372 25412
rect 2924 25372 2930 25384
rect 14366 25372 14372 25384
rect 14424 25372 14430 25424
rect 1857 25347 1915 25353
rect 1857 25313 1869 25347
rect 1903 25344 1915 25347
rect 8294 25344 8300 25356
rect 1903 25316 2544 25344
rect 1903 25313 1915 25316
rect 1857 25307 1915 25313
rect 1673 25279 1731 25285
rect 1673 25245 1685 25279
rect 1719 25245 1731 25279
rect 2314 25276 2320 25288
rect 2275 25248 2320 25276
rect 1673 25239 1731 25245
rect 2314 25236 2320 25248
rect 2372 25236 2378 25288
rect 2516 25285 2544 25316
rect 6748 25316 8300 25344
rect 2501 25279 2559 25285
rect 2501 25245 2513 25279
rect 2547 25245 2559 25279
rect 2501 25239 2559 25245
rect 2593 25279 2651 25285
rect 2593 25245 2605 25279
rect 2639 25245 2651 25279
rect 2593 25239 2651 25245
rect 2685 25279 2743 25285
rect 2685 25245 2697 25279
rect 2731 25276 2743 25279
rect 5353 25279 5411 25285
rect 2731 25248 3924 25276
rect 2731 25245 2743 25248
rect 2685 25239 2743 25245
rect 1489 25211 1547 25217
rect 1489 25177 1501 25211
rect 1535 25177 1547 25211
rect 2608 25208 2636 25239
rect 1489 25171 1547 25177
rect 2516 25180 2636 25208
rect 1504 25140 1532 25171
rect 2516 25152 2544 25180
rect 1670 25140 1676 25152
rect 1504 25112 1676 25140
rect 1670 25100 1676 25112
rect 1728 25100 1734 25152
rect 2498 25100 2504 25152
rect 2556 25100 2562 25152
rect 3896 25149 3924 25248
rect 5353 25245 5365 25279
rect 5399 25276 5411 25279
rect 5442 25276 5448 25288
rect 5399 25248 5448 25276
rect 5399 25245 5411 25248
rect 5353 25239 5411 25245
rect 5442 25236 5448 25248
rect 5500 25276 5506 25288
rect 6748 25276 6776 25316
rect 8294 25304 8300 25316
rect 8352 25304 8358 25356
rect 14090 25344 14096 25356
rect 14051 25316 14096 25344
rect 14090 25304 14096 25316
rect 14148 25304 14154 25356
rect 5500 25248 6776 25276
rect 7285 25279 7343 25285
rect 5500 25236 5506 25248
rect 7285 25245 7297 25279
rect 7331 25276 7343 25279
rect 7558 25276 7564 25288
rect 7331 25248 7564 25276
rect 7331 25245 7343 25248
rect 7285 25239 7343 25245
rect 5620 25211 5678 25217
rect 5620 25177 5632 25211
rect 5666 25208 5678 25211
rect 7006 25208 7012 25220
rect 5666 25180 7012 25208
rect 5666 25177 5678 25180
rect 5620 25171 5678 25177
rect 7006 25168 7012 25180
rect 7064 25168 7070 25220
rect 3881 25143 3939 25149
rect 3881 25109 3893 25143
rect 3927 25140 3939 25143
rect 7300 25140 7328 25239
rect 7558 25236 7564 25248
rect 7616 25236 7622 25288
rect 7742 25276 7748 25288
rect 7703 25248 7748 25276
rect 7742 25236 7748 25248
rect 7800 25236 7806 25288
rect 7906 25276 7912 25288
rect 7867 25248 7912 25276
rect 7906 25236 7912 25248
rect 7964 25236 7970 25288
rect 8202 25285 8208 25288
rect 8005 25233 8011 25285
rect 8063 25273 8069 25285
rect 8159 25279 8208 25285
rect 8063 25245 8108 25273
rect 8159 25245 8171 25279
rect 8205 25245 8208 25279
rect 8063 25233 8069 25245
rect 8159 25239 8208 25245
rect 8202 25236 8208 25239
rect 8260 25236 8266 25288
rect 8846 25236 8852 25288
rect 8904 25276 8910 25288
rect 8941 25279 8999 25285
rect 8941 25276 8953 25279
rect 8904 25248 8953 25276
rect 8904 25236 8910 25248
rect 8941 25245 8953 25248
rect 8987 25245 8999 25279
rect 9122 25276 9128 25288
rect 9083 25248 9128 25276
rect 8941 25239 8999 25245
rect 9122 25236 9128 25248
rect 9180 25236 9186 25288
rect 13170 25285 13176 25288
rect 13153 25279 13176 25285
rect 13153 25245 13165 25279
rect 13153 25239 13176 25245
rect 13170 25236 13176 25239
rect 13228 25236 13234 25288
rect 13262 25279 13320 25285
rect 13262 25245 13274 25279
rect 13308 25245 13320 25279
rect 13262 25239 13320 25245
rect 8478 25168 8484 25220
rect 8536 25208 8542 25220
rect 12986 25208 12992 25220
rect 8536 25180 12992 25208
rect 8536 25168 8542 25180
rect 12986 25168 12992 25180
rect 13044 25168 13050 25220
rect 13280 25208 13308 25239
rect 13354 25236 13360 25288
rect 13412 25285 13418 25288
rect 13412 25276 13420 25285
rect 13541 25279 13599 25285
rect 13412 25248 13457 25276
rect 13412 25239 13420 25248
rect 13541 25245 13553 25279
rect 13587 25276 13599 25279
rect 13906 25276 13912 25288
rect 13587 25248 13912 25276
rect 13587 25245 13599 25248
rect 13541 25239 13599 25245
rect 13412 25236 13418 25239
rect 13906 25236 13912 25248
rect 13964 25236 13970 25288
rect 14366 25276 14372 25288
rect 14327 25248 14372 25276
rect 14366 25236 14372 25248
rect 14424 25236 14430 25288
rect 16942 25236 16948 25288
rect 17000 25276 17006 25288
rect 17144 25285 17172 25452
rect 18874 25440 18880 25452
rect 18932 25480 18938 25492
rect 20625 25483 20683 25489
rect 20625 25480 20637 25483
rect 18932 25452 20637 25480
rect 18932 25440 18938 25452
rect 20625 25449 20637 25452
rect 20671 25449 20683 25483
rect 20625 25443 20683 25449
rect 27246 25440 27252 25492
rect 27304 25480 27310 25492
rect 27341 25483 27399 25489
rect 27341 25480 27353 25483
rect 27304 25452 27353 25480
rect 27304 25440 27310 25452
rect 27341 25449 27353 25452
rect 27387 25449 27399 25483
rect 27341 25443 27399 25449
rect 27522 25440 27528 25492
rect 27580 25480 27586 25492
rect 29917 25483 29975 25489
rect 29917 25480 29929 25483
rect 27580 25452 29929 25480
rect 27580 25440 27586 25452
rect 29917 25449 29929 25452
rect 29963 25480 29975 25483
rect 30558 25480 30564 25492
rect 29963 25452 30564 25480
rect 29963 25449 29975 25452
rect 29917 25443 29975 25449
rect 30558 25440 30564 25452
rect 30616 25440 30622 25492
rect 18325 25415 18383 25421
rect 18325 25381 18337 25415
rect 18371 25412 18383 25415
rect 19242 25412 19248 25424
rect 18371 25384 19248 25412
rect 18371 25381 18383 25384
rect 18325 25375 18383 25381
rect 19242 25372 19248 25384
rect 19300 25372 19306 25424
rect 20530 25412 20536 25424
rect 19536 25384 20536 25412
rect 17218 25304 17224 25356
rect 17276 25344 17282 25356
rect 17276 25316 17545 25344
rect 17276 25304 17282 25316
rect 17037 25279 17095 25285
rect 17037 25276 17049 25279
rect 17000 25248 17049 25276
rect 17000 25236 17006 25248
rect 17037 25245 17049 25248
rect 17083 25245 17095 25279
rect 17037 25239 17095 25245
rect 17130 25279 17188 25285
rect 17130 25245 17142 25279
rect 17176 25245 17188 25279
rect 17310 25276 17316 25288
rect 17271 25248 17316 25276
rect 17130 25239 17188 25245
rect 17310 25236 17316 25248
rect 17368 25236 17374 25288
rect 17517 25285 17545 25316
rect 17770 25304 17776 25356
rect 17828 25344 17834 25356
rect 17828 25316 18552 25344
rect 17828 25304 17834 25316
rect 18524 25285 18552 25316
rect 17517 25279 17579 25285
rect 17517 25248 17533 25279
rect 17521 25245 17533 25248
rect 17567 25245 17579 25279
rect 17521 25239 17579 25245
rect 18509 25279 18567 25285
rect 18509 25245 18521 25279
rect 18555 25245 18567 25279
rect 18509 25239 18567 25245
rect 18598 25236 18604 25288
rect 18656 25276 18662 25288
rect 18656 25248 18701 25276
rect 18656 25236 18662 25248
rect 19426 25236 19432 25288
rect 19484 25276 19490 25288
rect 19536 25285 19564 25384
rect 20530 25372 20536 25384
rect 20588 25372 20594 25424
rect 26878 25372 26884 25424
rect 26936 25412 26942 25424
rect 30377 25415 30435 25421
rect 30377 25412 30389 25415
rect 26936 25384 30389 25412
rect 26936 25372 26942 25384
rect 30377 25381 30389 25384
rect 30423 25412 30435 25415
rect 30423 25384 31319 25412
rect 30423 25381 30435 25384
rect 30377 25375 30435 25381
rect 20346 25344 20352 25356
rect 19812 25316 20352 25344
rect 19521 25279 19579 25285
rect 19521 25276 19533 25279
rect 19484 25248 19533 25276
rect 19484 25236 19490 25248
rect 19521 25245 19533 25248
rect 19567 25245 19579 25279
rect 19702 25276 19708 25288
rect 19663 25248 19708 25276
rect 19521 25239 19579 25245
rect 19702 25236 19708 25248
rect 19760 25236 19766 25288
rect 19812 25285 19840 25316
rect 20346 25304 20352 25316
rect 20404 25304 20410 25356
rect 31291 25344 31319 25384
rect 31291 25316 31340 25344
rect 19797 25279 19855 25285
rect 19797 25245 19809 25279
rect 19843 25245 19855 25279
rect 19797 25239 19855 25245
rect 19889 25279 19947 25285
rect 19889 25245 19901 25279
rect 19935 25276 19947 25279
rect 20530 25276 20536 25288
rect 19935 25248 20536 25276
rect 19935 25245 19947 25248
rect 19889 25239 19947 25245
rect 20530 25236 20536 25248
rect 20588 25236 20594 25288
rect 22005 25279 22063 25285
rect 22005 25245 22017 25279
rect 22051 25276 22063 25279
rect 22738 25276 22744 25288
rect 22051 25248 22744 25276
rect 22051 25245 22063 25248
rect 22005 25239 22063 25245
rect 22738 25236 22744 25248
rect 22796 25276 22802 25288
rect 23845 25279 23903 25285
rect 23845 25276 23857 25279
rect 22796 25248 23857 25276
rect 22796 25236 22802 25248
rect 23845 25245 23857 25248
rect 23891 25245 23903 25279
rect 23845 25239 23903 25245
rect 25409 25279 25467 25285
rect 25409 25245 25421 25279
rect 25455 25276 25467 25279
rect 25455 25248 26648 25276
rect 25455 25245 25467 25248
rect 25409 25239 25467 25245
rect 15010 25208 15016 25220
rect 13280 25180 15016 25208
rect 15010 25168 15016 25180
rect 15068 25168 15074 25220
rect 17402 25208 17408 25220
rect 17363 25180 17408 25208
rect 17402 25168 17408 25180
rect 17460 25168 17466 25220
rect 20165 25211 20223 25217
rect 20165 25177 20177 25211
rect 20211 25208 20223 25211
rect 21738 25211 21796 25217
rect 21738 25208 21750 25211
rect 20211 25180 21750 25208
rect 20211 25177 20223 25180
rect 20165 25171 20223 25177
rect 21738 25177 21750 25180
rect 21784 25177 21796 25211
rect 21738 25171 21796 25177
rect 23474 25168 23480 25220
rect 23532 25208 23538 25220
rect 23578 25211 23636 25217
rect 23578 25208 23590 25211
rect 23532 25180 23590 25208
rect 23532 25168 23538 25180
rect 23578 25177 23590 25180
rect 23624 25177 23636 25211
rect 23578 25171 23636 25177
rect 25593 25211 25651 25217
rect 25593 25177 25605 25211
rect 25639 25208 25651 25211
rect 26142 25208 26148 25220
rect 25639 25180 26148 25208
rect 25639 25177 25651 25180
rect 25593 25171 25651 25177
rect 26142 25168 26148 25180
rect 26200 25168 26206 25220
rect 26620 25208 26648 25248
rect 26694 25236 26700 25288
rect 26752 25276 26758 25288
rect 27154 25276 27160 25288
rect 26752 25248 27160 25276
rect 26752 25236 26758 25248
rect 27154 25236 27160 25248
rect 27212 25236 27218 25288
rect 29454 25236 29460 25288
rect 29512 25276 29518 25288
rect 30098 25276 30104 25288
rect 29512 25248 30104 25276
rect 29512 25236 29518 25248
rect 30098 25236 30104 25248
rect 30156 25276 30162 25288
rect 31312 25285 31340 25316
rect 30929 25279 30987 25285
rect 31208 25279 31266 25285
rect 30929 25276 30941 25279
rect 30156 25248 30941 25276
rect 30156 25236 30162 25248
rect 30929 25245 30941 25248
rect 30975 25245 30987 25279
rect 30929 25239 30987 25245
rect 31113 25273 31171 25279
rect 31113 25239 31125 25273
rect 31159 25239 31171 25273
rect 31208 25245 31220 25279
rect 31254 25245 31266 25279
rect 31208 25239 31266 25245
rect 31297 25279 31355 25285
rect 31297 25245 31309 25279
rect 31343 25245 31355 25279
rect 31297 25239 31355 25245
rect 33413 25279 33471 25285
rect 33413 25245 33425 25279
rect 33459 25276 33471 25279
rect 33962 25276 33968 25288
rect 33459 25248 33968 25276
rect 33459 25245 33471 25248
rect 33413 25239 33471 25245
rect 31113 25233 31171 25239
rect 26970 25208 26976 25220
rect 26620 25180 26976 25208
rect 26970 25168 26976 25180
rect 27028 25168 27034 25220
rect 31128 25152 31156 25233
rect 31211 25208 31239 25239
rect 33962 25236 33968 25248
rect 34020 25236 34026 25288
rect 68094 25276 68100 25288
rect 68055 25248 68100 25276
rect 68094 25236 68100 25248
rect 68152 25236 68158 25288
rect 31386 25208 31392 25220
rect 31211 25180 31392 25208
rect 31386 25168 31392 25180
rect 31444 25168 31450 25220
rect 31573 25211 31631 25217
rect 31573 25177 31585 25211
rect 31619 25208 31631 25211
rect 33146 25211 33204 25217
rect 33146 25208 33158 25211
rect 31619 25180 33158 25208
rect 31619 25177 31631 25180
rect 31573 25171 31631 25177
rect 33146 25177 33158 25180
rect 33192 25177 33204 25211
rect 33146 25171 33204 25177
rect 3927 25112 7328 25140
rect 3927 25109 3939 25112
rect 3881 25103 3939 25109
rect 7926 25100 7932 25152
rect 7984 25140 7990 25152
rect 9309 25143 9367 25149
rect 9309 25140 9321 25143
rect 7984 25112 9321 25140
rect 7984 25100 7990 25112
rect 9309 25109 9321 25112
rect 9355 25109 9367 25143
rect 9858 25140 9864 25152
rect 9819 25112 9864 25140
rect 9309 25103 9367 25109
rect 9858 25100 9864 25112
rect 9916 25100 9922 25152
rect 15378 25100 15384 25152
rect 15436 25140 15442 25152
rect 15930 25140 15936 25152
rect 15436 25112 15936 25140
rect 15436 25100 15442 25112
rect 15930 25100 15936 25112
rect 15988 25100 15994 25152
rect 17678 25140 17684 25152
rect 17639 25112 17684 25140
rect 17678 25100 17684 25112
rect 17736 25100 17742 25152
rect 22465 25143 22523 25149
rect 22465 25109 22477 25143
rect 22511 25140 22523 25143
rect 23290 25140 23296 25152
rect 22511 25112 23296 25140
rect 22511 25109 22523 25112
rect 22465 25103 22523 25109
rect 23290 25100 23296 25112
rect 23348 25100 23354 25152
rect 25682 25100 25688 25152
rect 25740 25140 25746 25152
rect 25777 25143 25835 25149
rect 25777 25140 25789 25143
rect 25740 25112 25789 25140
rect 25740 25100 25746 25112
rect 25777 25109 25789 25112
rect 25823 25109 25835 25143
rect 26326 25140 26332 25152
rect 26287 25112 26332 25140
rect 25777 25103 25835 25109
rect 26326 25100 26332 25112
rect 26384 25100 26390 25152
rect 31110 25100 31116 25152
rect 31168 25100 31174 25152
rect 31662 25100 31668 25152
rect 31720 25140 31726 25152
rect 32033 25143 32091 25149
rect 32033 25140 32045 25143
rect 31720 25112 32045 25140
rect 31720 25100 31726 25112
rect 32033 25109 32045 25112
rect 32079 25109 32091 25143
rect 32033 25103 32091 25109
rect 1104 25050 68816 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 68816 25050
rect 1104 24976 68816 24998
rect 7558 24896 7564 24948
rect 7616 24936 7622 24948
rect 8202 24936 8208 24948
rect 7616 24908 8208 24936
rect 7616 24896 7622 24908
rect 8202 24896 8208 24908
rect 8260 24896 8266 24948
rect 9858 24896 9864 24948
rect 9916 24896 9922 24948
rect 12618 24936 12624 24948
rect 12579 24908 12624 24936
rect 12618 24896 12624 24908
rect 12676 24896 12682 24948
rect 15930 24896 15936 24948
rect 15988 24936 15994 24948
rect 16114 24936 16120 24948
rect 15988 24908 16120 24936
rect 15988 24896 15994 24908
rect 16114 24896 16120 24908
rect 16172 24936 16178 24948
rect 22186 24936 22192 24948
rect 16172 24908 22192 24936
rect 16172 24896 16178 24908
rect 22186 24896 22192 24908
rect 22244 24896 22250 24948
rect 23474 24936 23480 24948
rect 23435 24908 23480 24936
rect 23474 24896 23480 24908
rect 23532 24896 23538 24948
rect 24949 24939 25007 24945
rect 24949 24905 24961 24939
rect 24995 24936 25007 24939
rect 26050 24936 26056 24948
rect 24995 24908 26056 24936
rect 24995 24905 25007 24908
rect 24949 24899 25007 24905
rect 26050 24896 26056 24908
rect 26108 24896 26114 24948
rect 31110 24936 31116 24948
rect 31071 24908 31116 24936
rect 31110 24896 31116 24908
rect 31168 24896 31174 24948
rect 1397 24871 1455 24877
rect 1397 24837 1409 24871
rect 1443 24868 1455 24871
rect 1670 24868 1676 24880
rect 1443 24840 1676 24868
rect 1443 24837 1455 24840
rect 1397 24831 1455 24837
rect 1670 24828 1676 24840
rect 1728 24828 1734 24880
rect 1765 24871 1823 24877
rect 1765 24837 1777 24871
rect 1811 24868 1823 24871
rect 3234 24868 3240 24880
rect 1811 24840 3240 24868
rect 1811 24837 1823 24840
rect 1765 24831 1823 24837
rect 3234 24828 3240 24840
rect 3292 24828 3298 24880
rect 5442 24868 5448 24880
rect 3988 24840 5448 24868
rect 1581 24803 1639 24809
rect 1581 24769 1593 24803
rect 1627 24769 1639 24803
rect 1581 24763 1639 24769
rect 2225 24803 2283 24809
rect 2225 24769 2237 24803
rect 2271 24769 2283 24803
rect 2406 24800 2412 24812
rect 2367 24772 2412 24800
rect 2225 24763 2283 24769
rect 1596 24664 1624 24763
rect 2240 24732 2268 24763
rect 2406 24760 2412 24772
rect 2464 24760 2470 24812
rect 2498 24760 2504 24812
rect 2556 24800 2562 24812
rect 2639 24803 2697 24809
rect 2556 24772 2601 24800
rect 2556 24760 2562 24772
rect 2639 24769 2651 24803
rect 2685 24800 2697 24803
rect 3694 24800 3700 24812
rect 2685 24772 3700 24800
rect 2685 24769 2697 24772
rect 2639 24763 2697 24769
rect 3694 24760 3700 24772
rect 3752 24760 3758 24812
rect 3789 24803 3847 24809
rect 3789 24769 3801 24803
rect 3835 24800 3847 24803
rect 3988 24800 4016 24840
rect 5442 24828 5448 24840
rect 5500 24828 5506 24880
rect 5534 24828 5540 24880
rect 5592 24868 5598 24880
rect 9876 24868 9904 24896
rect 5592 24840 9904 24868
rect 12176 24840 12388 24868
rect 5592 24828 5598 24840
rect 4062 24809 4068 24812
rect 3835 24772 4016 24800
rect 3835 24769 3847 24772
rect 3789 24763 3847 24769
rect 4056 24763 4068 24809
rect 4120 24800 4126 24812
rect 7101 24803 7159 24809
rect 4120 24772 4156 24800
rect 4062 24760 4068 24763
rect 4120 24760 4126 24772
rect 7101 24769 7113 24803
rect 7147 24800 7159 24803
rect 7742 24800 7748 24812
rect 7147 24772 7748 24800
rect 7147 24769 7159 24772
rect 7101 24763 7159 24769
rect 7742 24760 7748 24772
rect 7800 24760 7806 24812
rect 8478 24800 8484 24812
rect 8439 24772 8484 24800
rect 8478 24760 8484 24772
rect 8536 24760 8542 24812
rect 8662 24800 8668 24812
rect 8623 24772 8668 24800
rect 8662 24760 8668 24772
rect 8720 24760 8726 24812
rect 8864 24809 8892 24840
rect 8757 24803 8815 24809
rect 8757 24769 8769 24803
rect 8803 24769 8815 24803
rect 8757 24763 8815 24769
rect 8849 24803 8907 24809
rect 8849 24769 8861 24803
rect 8895 24769 8907 24803
rect 9841 24803 9899 24809
rect 9841 24800 9853 24803
rect 8849 24763 8907 24769
rect 9140 24772 9853 24800
rect 2314 24732 2320 24744
rect 2240 24704 2320 24732
rect 2314 24692 2320 24704
rect 2372 24692 2378 24744
rect 2869 24735 2927 24741
rect 2700 24704 2820 24732
rect 2700 24664 2728 24704
rect 1596 24636 2728 24664
rect 2792 24596 2820 24704
rect 2869 24701 2881 24735
rect 2915 24732 2927 24735
rect 3050 24732 3056 24744
rect 2915 24704 3056 24732
rect 2915 24701 2927 24704
rect 2869 24695 2927 24701
rect 3050 24692 3056 24704
rect 3108 24692 3114 24744
rect 6270 24692 6276 24744
rect 6328 24732 6334 24744
rect 6825 24735 6883 24741
rect 6825 24732 6837 24735
rect 6328 24704 6837 24732
rect 6328 24692 6334 24704
rect 6825 24701 6837 24704
rect 6871 24701 6883 24735
rect 6825 24695 6883 24701
rect 8018 24692 8024 24744
rect 8076 24732 8082 24744
rect 8570 24732 8576 24744
rect 8076 24704 8576 24732
rect 8076 24692 8082 24704
rect 8570 24692 8576 24704
rect 8628 24732 8634 24744
rect 8772 24732 8800 24763
rect 9140 24741 9168 24772
rect 9841 24769 9853 24772
rect 9887 24769 9899 24803
rect 9841 24763 9899 24769
rect 10410 24760 10416 24812
rect 10468 24800 10474 24812
rect 12066 24800 12072 24812
rect 10468 24772 12072 24800
rect 10468 24760 10474 24772
rect 12066 24760 12072 24772
rect 12124 24760 12130 24812
rect 8628 24704 8800 24732
rect 9125 24735 9183 24741
rect 8628 24692 8634 24704
rect 9125 24701 9137 24735
rect 9171 24701 9183 24735
rect 9125 24695 9183 24701
rect 9398 24692 9404 24744
rect 9456 24732 9462 24744
rect 9585 24735 9643 24741
rect 9585 24732 9597 24735
rect 9456 24704 9597 24732
rect 9456 24692 9462 24704
rect 9585 24701 9597 24704
rect 9631 24701 9643 24735
rect 9585 24695 9643 24701
rect 12176 24664 12204 24840
rect 12360 24809 12388 24840
rect 13170 24828 13176 24880
rect 13228 24868 13234 24880
rect 16022 24868 16028 24880
rect 13228 24840 16028 24868
rect 13228 24828 13234 24840
rect 16022 24828 16028 24840
rect 16080 24828 16086 24880
rect 16206 24828 16212 24880
rect 16264 24868 16270 24880
rect 18049 24871 18107 24877
rect 18049 24868 18061 24871
rect 16264 24840 18061 24868
rect 16264 24828 16270 24840
rect 18049 24837 18061 24840
rect 18095 24868 18107 24871
rect 18598 24868 18604 24880
rect 18095 24840 18604 24868
rect 18095 24837 18107 24840
rect 18049 24831 18107 24837
rect 18598 24828 18604 24840
rect 18656 24828 18662 24880
rect 26326 24868 26332 24880
rect 19628 24840 20024 24868
rect 12253 24803 12311 24809
rect 12253 24769 12265 24803
rect 12299 24769 12311 24803
rect 12253 24763 12311 24769
rect 12345 24803 12403 24809
rect 12345 24769 12357 24803
rect 12391 24769 12403 24803
rect 12345 24763 12403 24769
rect 12437 24803 12495 24809
rect 12437 24769 12449 24803
rect 12483 24800 12495 24803
rect 13633 24803 13691 24809
rect 13633 24800 13645 24803
rect 12483 24772 13645 24800
rect 12483 24769 12495 24772
rect 12437 24763 12495 24769
rect 13633 24769 13645 24772
rect 13679 24800 13691 24803
rect 13722 24800 13728 24812
rect 13679 24772 13728 24800
rect 13679 24769 13691 24772
rect 13633 24763 13691 24769
rect 12268 24732 12296 24763
rect 13722 24760 13728 24772
rect 13780 24760 13786 24812
rect 14366 24800 14372 24812
rect 13832 24772 14372 24800
rect 13832 24732 13860 24772
rect 14366 24760 14372 24772
rect 14424 24760 14430 24812
rect 15470 24760 15476 24812
rect 15528 24800 15534 24812
rect 15850 24803 15908 24809
rect 15850 24800 15862 24803
rect 15528 24772 15862 24800
rect 15528 24760 15534 24772
rect 15850 24769 15862 24772
rect 15896 24769 15908 24803
rect 15850 24763 15908 24769
rect 16117 24803 16175 24809
rect 16117 24769 16129 24803
rect 16163 24800 16175 24803
rect 19628 24800 19656 24840
rect 16163 24772 19656 24800
rect 16163 24769 16175 24772
rect 16117 24763 16175 24769
rect 19702 24760 19708 24812
rect 19760 24809 19766 24812
rect 19996 24809 20024 24840
rect 25976 24840 26332 24868
rect 19760 24800 19772 24809
rect 19981 24803 20039 24809
rect 19760 24772 19805 24800
rect 19760 24763 19772 24772
rect 19981 24769 19993 24803
rect 20027 24800 20039 24803
rect 20622 24800 20628 24812
rect 20027 24772 20628 24800
rect 20027 24769 20039 24772
rect 19981 24763 20039 24769
rect 19760 24760 19766 24763
rect 20622 24760 20628 24772
rect 20680 24760 20686 24812
rect 22278 24760 22284 24812
rect 22336 24800 22342 24812
rect 23750 24800 23756 24812
rect 22336 24772 23756 24800
rect 22336 24760 22342 24772
rect 23750 24760 23756 24772
rect 23808 24760 23814 24812
rect 23842 24803 23900 24809
rect 23842 24769 23854 24803
rect 23888 24769 23900 24803
rect 23842 24763 23900 24769
rect 12268 24704 13860 24732
rect 13909 24735 13967 24741
rect 13909 24701 13921 24735
rect 13955 24732 13967 24735
rect 14274 24732 14280 24744
rect 13955 24704 14280 24732
rect 13955 24701 13967 24704
rect 13909 24695 13967 24701
rect 14274 24692 14280 24704
rect 14332 24692 14338 24744
rect 23658 24692 23664 24744
rect 23716 24732 23722 24744
rect 23857 24732 23885 24763
rect 23934 24760 23940 24812
rect 23992 24809 23998 24812
rect 23992 24800 24000 24809
rect 24121 24803 24179 24809
rect 23992 24772 24037 24800
rect 23992 24763 24000 24772
rect 24121 24769 24133 24803
rect 24167 24800 24179 24803
rect 24210 24800 24216 24812
rect 24167 24772 24216 24800
rect 24167 24769 24179 24772
rect 24121 24763 24179 24769
rect 23992 24760 23998 24763
rect 24210 24760 24216 24772
rect 24268 24800 24274 24812
rect 24578 24800 24584 24812
rect 24268 24772 24584 24800
rect 24268 24760 24274 24772
rect 24578 24760 24584 24772
rect 24636 24760 24642 24812
rect 24854 24760 24860 24812
rect 24912 24800 24918 24812
rect 25041 24803 25099 24809
rect 25041 24800 25053 24803
rect 24912 24772 25053 24800
rect 24912 24760 24918 24772
rect 25041 24769 25053 24772
rect 25087 24769 25099 24803
rect 25041 24763 25099 24769
rect 25406 24760 25412 24812
rect 25464 24800 25470 24812
rect 25593 24803 25651 24809
rect 25593 24800 25605 24803
rect 25464 24772 25605 24800
rect 25464 24760 25470 24772
rect 25593 24769 25605 24772
rect 25639 24769 25651 24803
rect 25593 24763 25651 24769
rect 25682 24760 25688 24812
rect 25740 24800 25746 24812
rect 25976 24809 26004 24840
rect 26326 24828 26332 24840
rect 26384 24828 26390 24880
rect 29822 24868 29828 24880
rect 29196 24840 29828 24868
rect 25777 24803 25835 24809
rect 25777 24800 25789 24803
rect 25740 24772 25789 24800
rect 25740 24760 25746 24772
rect 25777 24769 25789 24772
rect 25823 24769 25835 24803
rect 25777 24763 25835 24769
rect 25872 24803 25930 24809
rect 25872 24769 25884 24803
rect 25918 24769 25930 24803
rect 25872 24763 25930 24769
rect 25961 24803 26019 24809
rect 25961 24769 25973 24803
rect 26007 24769 26019 24803
rect 28086 24803 28144 24809
rect 28086 24800 28098 24803
rect 25961 24763 26019 24769
rect 26252 24772 28098 24800
rect 23716 24704 23885 24732
rect 23716 24692 23722 24704
rect 25884 24664 25912 24763
rect 26252 24741 26280 24772
rect 28086 24769 28098 24772
rect 28132 24769 28144 24803
rect 28086 24763 28144 24769
rect 28994 24760 29000 24812
rect 29052 24800 29058 24812
rect 29196 24809 29224 24840
rect 29822 24828 29828 24840
rect 29880 24828 29886 24880
rect 30745 24871 30803 24877
rect 30745 24837 30757 24871
rect 30791 24868 30803 24871
rect 31018 24868 31024 24880
rect 30791 24840 31024 24868
rect 30791 24837 30803 24840
rect 30745 24831 30803 24837
rect 29089 24803 29147 24809
rect 29089 24800 29101 24803
rect 29052 24772 29101 24800
rect 29052 24760 29058 24772
rect 29089 24769 29101 24772
rect 29135 24769 29147 24803
rect 29089 24763 29147 24769
rect 29181 24803 29239 24809
rect 29181 24769 29193 24803
rect 29227 24769 29239 24803
rect 29181 24763 29239 24769
rect 29273 24803 29331 24809
rect 29273 24769 29285 24803
rect 29319 24769 29331 24803
rect 29454 24800 29460 24812
rect 29415 24772 29460 24800
rect 29273 24763 29331 24769
rect 26237 24735 26295 24741
rect 26237 24701 26249 24735
rect 26283 24701 26295 24735
rect 26237 24695 26295 24701
rect 28353 24735 28411 24741
rect 28353 24701 28365 24735
rect 28399 24701 28411 24735
rect 29288 24732 29316 24763
rect 29454 24760 29460 24772
rect 29512 24760 29518 24812
rect 30006 24760 30012 24812
rect 30064 24800 30070 24812
rect 30101 24803 30159 24809
rect 30101 24800 30113 24803
rect 30064 24772 30113 24800
rect 30064 24760 30070 24772
rect 30101 24769 30113 24772
rect 30147 24769 30159 24803
rect 30101 24763 30159 24769
rect 30285 24803 30343 24809
rect 30285 24769 30297 24803
rect 30331 24800 30343 24803
rect 30760 24800 30788 24831
rect 31018 24828 31024 24840
rect 31076 24828 31082 24880
rect 30331 24772 30788 24800
rect 30929 24803 30987 24809
rect 30331 24769 30343 24772
rect 30285 24763 30343 24769
rect 30929 24769 30941 24803
rect 30975 24800 30987 24803
rect 31662 24800 31668 24812
rect 30975 24772 31668 24800
rect 30975 24769 30987 24772
rect 30929 24763 30987 24769
rect 31662 24760 31668 24772
rect 31720 24760 31726 24812
rect 29917 24735 29975 24741
rect 29917 24732 29929 24735
rect 29288 24704 29929 24732
rect 28353 24695 28411 24701
rect 29917 24701 29929 24704
rect 29963 24701 29975 24735
rect 29917 24695 29975 24701
rect 26050 24664 26056 24676
rect 10520 24636 12204 24664
rect 12544 24636 14872 24664
rect 25884 24636 26056 24664
rect 5169 24599 5227 24605
rect 5169 24596 5181 24599
rect 2792 24568 5181 24596
rect 5169 24565 5181 24568
rect 5215 24596 5227 24599
rect 10520 24596 10548 24636
rect 10962 24596 10968 24608
rect 5215 24568 10548 24596
rect 10923 24568 10968 24596
rect 5215 24565 5227 24568
rect 5169 24559 5227 24565
rect 10962 24556 10968 24568
rect 11020 24596 11026 24608
rect 12544 24596 12572 24636
rect 14734 24596 14740 24608
rect 11020 24568 12572 24596
rect 14695 24568 14740 24596
rect 11020 24556 11026 24568
rect 14734 24556 14740 24568
rect 14792 24556 14798 24608
rect 14844 24596 14872 24636
rect 26050 24624 26056 24636
rect 26108 24624 26114 24676
rect 17034 24596 17040 24608
rect 14844 24568 17040 24596
rect 17034 24556 17040 24568
rect 17092 24556 17098 24608
rect 18230 24556 18236 24608
rect 18288 24596 18294 24608
rect 18601 24599 18659 24605
rect 18601 24596 18613 24599
rect 18288 24568 18613 24596
rect 18288 24556 18294 24568
rect 18601 24565 18613 24568
rect 18647 24565 18659 24599
rect 20530 24596 20536 24608
rect 20491 24568 20536 24596
rect 18601 24559 18659 24565
rect 20530 24556 20536 24568
rect 20588 24556 20594 24608
rect 21818 24596 21824 24608
rect 21779 24568 21824 24596
rect 21818 24556 21824 24568
rect 21876 24556 21882 24608
rect 26142 24556 26148 24608
rect 26200 24596 26206 24608
rect 26602 24596 26608 24608
rect 26200 24568 26608 24596
rect 26200 24556 26206 24568
rect 26602 24556 26608 24568
rect 26660 24596 26666 24608
rect 26973 24599 27031 24605
rect 26973 24596 26985 24599
rect 26660 24568 26985 24596
rect 26660 24556 26666 24568
rect 26973 24565 26985 24568
rect 27019 24565 27031 24599
rect 26973 24559 27031 24565
rect 27062 24556 27068 24608
rect 27120 24596 27126 24608
rect 28368 24596 28396 24695
rect 28810 24596 28816 24608
rect 27120 24568 28396 24596
rect 28771 24568 28816 24596
rect 27120 24556 27126 24568
rect 28810 24556 28816 24568
rect 28868 24556 28874 24608
rect 1104 24506 68816 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 65654 24506
rect 65706 24454 65718 24506
rect 65770 24454 65782 24506
rect 65834 24454 65846 24506
rect 65898 24454 65910 24506
rect 65962 24454 68816 24506
rect 1104 24432 68816 24454
rect 3694 24352 3700 24404
rect 3752 24392 3758 24404
rect 3789 24395 3847 24401
rect 3789 24392 3801 24395
rect 3752 24364 3801 24392
rect 3752 24352 3758 24364
rect 3789 24361 3801 24364
rect 3835 24361 3847 24395
rect 7006 24392 7012 24404
rect 6967 24364 7012 24392
rect 3789 24355 3847 24361
rect 7006 24352 7012 24364
rect 7064 24352 7070 24404
rect 7098 24352 7104 24404
rect 7156 24392 7162 24404
rect 8110 24392 8116 24404
rect 7156 24364 8116 24392
rect 7156 24352 7162 24364
rect 8110 24352 8116 24364
rect 8168 24352 8174 24404
rect 8297 24395 8355 24401
rect 8297 24361 8309 24395
rect 8343 24392 8355 24395
rect 8846 24392 8852 24404
rect 8343 24364 8852 24392
rect 8343 24361 8355 24364
rect 8297 24355 8355 24361
rect 8846 24352 8852 24364
rect 8904 24352 8910 24404
rect 9030 24352 9036 24404
rect 9088 24392 9094 24404
rect 10962 24392 10968 24404
rect 9088 24364 10968 24392
rect 9088 24352 9094 24364
rect 10962 24352 10968 24364
rect 11020 24352 11026 24404
rect 12713 24395 12771 24401
rect 12713 24361 12725 24395
rect 12759 24392 12771 24395
rect 13354 24392 13360 24404
rect 12759 24364 13360 24392
rect 12759 24361 12771 24364
rect 12713 24355 12771 24361
rect 13354 24352 13360 24364
rect 13412 24352 13418 24404
rect 13541 24395 13599 24401
rect 13541 24361 13553 24395
rect 13587 24392 13599 24395
rect 19245 24395 19303 24401
rect 13587 24364 15792 24392
rect 13587 24361 13599 24364
rect 13541 24355 13599 24361
rect 2498 24284 2504 24336
rect 2556 24324 2562 24336
rect 3326 24324 3332 24336
rect 2556 24296 3332 24324
rect 2556 24284 2562 24296
rect 2976 24265 3004 24296
rect 3326 24284 3332 24296
rect 3384 24284 3390 24336
rect 7374 24284 7380 24336
rect 7432 24284 7438 24336
rect 10781 24327 10839 24333
rect 10781 24293 10793 24327
rect 10827 24324 10839 24327
rect 15562 24324 15568 24336
rect 10827 24296 15568 24324
rect 10827 24293 10839 24296
rect 10781 24287 10839 24293
rect 2961 24259 3019 24265
rect 2961 24225 2973 24259
rect 3007 24225 3019 24259
rect 2961 24219 3019 24225
rect 3237 24259 3295 24265
rect 3237 24225 3249 24259
rect 3283 24256 3295 24259
rect 3602 24256 3608 24268
rect 3283 24228 3608 24256
rect 3283 24225 3295 24228
rect 3237 24219 3295 24225
rect 3602 24216 3608 24228
rect 3660 24256 3666 24268
rect 3970 24256 3976 24268
rect 3660 24228 3976 24256
rect 3660 24216 3666 24228
rect 3970 24216 3976 24228
rect 4028 24216 4034 24268
rect 5166 24188 5172 24200
rect 3252 24160 5172 24188
rect 1581 24123 1639 24129
rect 1581 24089 1593 24123
rect 1627 24120 1639 24123
rect 1670 24120 1676 24132
rect 1627 24092 1676 24120
rect 1627 24089 1639 24092
rect 1581 24083 1639 24089
rect 1670 24080 1676 24092
rect 1728 24080 1734 24132
rect 1765 24123 1823 24129
rect 1765 24089 1777 24123
rect 1811 24120 1823 24123
rect 3252 24120 3280 24160
rect 5166 24148 5172 24160
rect 5224 24148 5230 24200
rect 7405 24197 7433 24284
rect 8220 24228 9536 24256
rect 7265 24191 7323 24197
rect 7265 24157 7277 24191
rect 7311 24188 7323 24191
rect 7377 24191 7435 24197
rect 7311 24157 7328 24188
rect 7265 24151 7328 24157
rect 7377 24157 7389 24191
rect 7423 24157 7435 24191
rect 7377 24151 7435 24157
rect 3878 24120 3884 24132
rect 1811 24092 3280 24120
rect 3344 24092 3884 24120
rect 1811 24089 1823 24092
rect 1765 24083 1823 24089
rect 1946 24052 1952 24064
rect 1907 24024 1952 24052
rect 1946 24012 1952 24024
rect 2004 24012 2010 24064
rect 2774 24012 2780 24064
rect 2832 24052 2838 24064
rect 3344 24052 3372 24092
rect 3878 24080 3884 24092
rect 3936 24120 3942 24132
rect 4341 24123 4399 24129
rect 4341 24120 4353 24123
rect 3936 24092 4353 24120
rect 3936 24080 3942 24092
rect 4341 24089 4353 24092
rect 4387 24089 4399 24123
rect 6270 24120 6276 24132
rect 6231 24092 6276 24120
rect 4341 24083 4399 24089
rect 6270 24080 6276 24092
rect 6328 24080 6334 24132
rect 7006 24080 7012 24132
rect 7064 24120 7070 24132
rect 7300 24120 7328 24151
rect 7466 24148 7472 24200
rect 7524 24197 7530 24200
rect 7524 24188 7532 24197
rect 7653 24191 7711 24197
rect 7524 24160 7569 24188
rect 7524 24151 7532 24160
rect 7653 24157 7665 24191
rect 7699 24188 7711 24191
rect 7742 24188 7748 24200
rect 7699 24160 7748 24188
rect 7699 24157 7711 24160
rect 7653 24151 7711 24157
rect 7524 24148 7530 24151
rect 7742 24148 7748 24160
rect 7800 24148 7806 24200
rect 8110 24188 8116 24200
rect 8071 24160 8116 24188
rect 8110 24148 8116 24160
rect 8168 24148 8174 24200
rect 8220 24120 8248 24228
rect 9398 24188 9404 24200
rect 9359 24160 9404 24188
rect 9398 24148 9404 24160
rect 9456 24148 9462 24200
rect 9508 24188 9536 24228
rect 10686 24188 10692 24200
rect 9508 24160 10692 24188
rect 10686 24148 10692 24160
rect 10744 24148 10750 24200
rect 7064 24092 8248 24120
rect 7064 24080 7070 24092
rect 8846 24080 8852 24132
rect 8904 24120 8910 24132
rect 9646 24123 9704 24129
rect 9646 24120 9658 24123
rect 8904 24092 9658 24120
rect 8904 24080 8910 24092
rect 9646 24089 9658 24092
rect 9692 24089 9704 24123
rect 9646 24083 9704 24089
rect 5718 24052 5724 24064
rect 2832 24024 3372 24052
rect 5679 24024 5724 24052
rect 2832 24012 2838 24024
rect 5718 24012 5724 24024
rect 5776 24012 5782 24064
rect 6365 24055 6423 24061
rect 6365 24021 6377 24055
rect 6411 24052 6423 24055
rect 7190 24052 7196 24064
rect 6411 24024 7196 24052
rect 6411 24021 6423 24024
rect 6365 24015 6423 24021
rect 7190 24012 7196 24024
rect 7248 24052 7254 24064
rect 7650 24052 7656 24064
rect 7248 24024 7656 24052
rect 7248 24012 7254 24024
rect 7650 24012 7656 24024
rect 7708 24012 7714 24064
rect 9306 24012 9312 24064
rect 9364 24052 9370 24064
rect 10796 24052 10824 24287
rect 15562 24284 15568 24296
rect 15620 24284 15626 24336
rect 15764 24324 15792 24364
rect 19245 24361 19257 24395
rect 19291 24392 19303 24395
rect 19702 24392 19708 24404
rect 19291 24364 19708 24392
rect 19291 24361 19303 24364
rect 19245 24355 19303 24361
rect 19702 24352 19708 24364
rect 19760 24352 19766 24404
rect 23753 24395 23811 24401
rect 23753 24361 23765 24395
rect 23799 24392 23811 24395
rect 23934 24392 23940 24404
rect 23799 24364 23940 24392
rect 23799 24361 23811 24364
rect 23753 24355 23811 24361
rect 23934 24352 23940 24364
rect 23992 24352 23998 24404
rect 26234 24352 26240 24404
rect 26292 24392 26298 24404
rect 26789 24395 26847 24401
rect 26789 24392 26801 24395
rect 26292 24364 26801 24392
rect 26292 24352 26298 24364
rect 26789 24361 26801 24364
rect 26835 24392 26847 24395
rect 26970 24392 26976 24404
rect 26835 24364 26976 24392
rect 26835 24361 26847 24364
rect 26789 24355 26847 24361
rect 26970 24352 26976 24364
rect 27028 24352 27034 24404
rect 27338 24352 27344 24404
rect 27396 24392 27402 24404
rect 30561 24395 30619 24401
rect 30561 24392 30573 24395
rect 27396 24364 30573 24392
rect 27396 24352 27402 24364
rect 30561 24361 30573 24364
rect 30607 24392 30619 24395
rect 30607 24364 31570 24392
rect 30607 24361 30619 24364
rect 30561 24355 30619 24361
rect 17218 24324 17224 24336
rect 15764 24296 17224 24324
rect 12618 24216 12624 24268
rect 12676 24256 12682 24268
rect 12676 24228 15608 24256
rect 12676 24216 12682 24228
rect 12066 24148 12072 24200
rect 12124 24188 12130 24200
rect 12529 24191 12587 24197
rect 12529 24188 12541 24191
rect 12124 24160 12541 24188
rect 12124 24148 12130 24160
rect 12529 24157 12541 24160
rect 12575 24157 12587 24191
rect 14274 24188 14280 24200
rect 14235 24160 14280 24188
rect 12529 24151 12587 24157
rect 14274 24148 14280 24160
rect 14332 24148 14338 24200
rect 15102 24148 15108 24200
rect 15160 24188 15166 24200
rect 15473 24191 15531 24197
rect 15473 24188 15485 24191
rect 15160 24160 15485 24188
rect 15160 24148 15166 24160
rect 15473 24157 15485 24160
rect 15519 24157 15531 24191
rect 15473 24151 15531 24157
rect 12345 24123 12403 24129
rect 12345 24089 12357 24123
rect 12391 24120 12403 24123
rect 13814 24120 13820 24132
rect 12391 24092 13820 24120
rect 12391 24089 12403 24092
rect 12345 24083 12403 24089
rect 12544 24064 12572 24092
rect 13814 24080 13820 24092
rect 13872 24080 13878 24132
rect 15580 24120 15608 24228
rect 15764 24197 15792 24296
rect 17218 24284 17224 24296
rect 17276 24284 17282 24336
rect 21269 24327 21327 24333
rect 21269 24293 21281 24327
rect 21315 24324 21327 24327
rect 22278 24324 22284 24336
rect 21315 24296 22284 24324
rect 21315 24293 21327 24296
rect 21269 24287 21327 24293
rect 22278 24284 22284 24296
rect 22336 24284 22342 24336
rect 26142 24284 26148 24336
rect 26200 24324 26206 24336
rect 27430 24324 27436 24336
rect 26200 24296 27436 24324
rect 26200 24284 26206 24296
rect 27430 24284 27436 24296
rect 27488 24324 27494 24336
rect 27488 24296 28028 24324
rect 27488 24284 27494 24296
rect 18322 24256 18328 24268
rect 16868 24228 18328 24256
rect 16868 24197 16896 24228
rect 18322 24216 18328 24228
rect 18380 24216 18386 24268
rect 18417 24259 18475 24265
rect 18417 24225 18429 24259
rect 18463 24256 18475 24259
rect 22189 24259 22247 24265
rect 22189 24256 22201 24259
rect 18463 24228 19748 24256
rect 18463 24225 18475 24228
rect 18417 24219 18475 24225
rect 15749 24191 15807 24197
rect 15749 24157 15761 24191
rect 15795 24157 15807 24191
rect 15749 24151 15807 24157
rect 16669 24191 16727 24197
rect 16669 24157 16681 24191
rect 16715 24157 16727 24191
rect 16669 24151 16727 24157
rect 16817 24191 16896 24197
rect 16817 24157 16829 24191
rect 16863 24160 16896 24191
rect 17034 24188 17040 24200
rect 16995 24160 17040 24188
rect 16863 24157 16875 24160
rect 16817 24151 16875 24157
rect 16684 24120 16712 24151
rect 17034 24148 17040 24160
rect 17092 24148 17098 24200
rect 17126 24148 17132 24200
rect 17184 24197 17190 24200
rect 17184 24188 17192 24197
rect 17586 24188 17592 24200
rect 17184 24160 17592 24188
rect 17184 24151 17192 24160
rect 17184 24148 17190 24151
rect 17586 24148 17592 24160
rect 17644 24148 17650 24200
rect 18230 24188 18236 24200
rect 18191 24160 18236 24188
rect 18230 24148 18236 24160
rect 18288 24148 18294 24200
rect 19334 24148 19340 24200
rect 19392 24188 19398 24200
rect 19720 24197 19748 24228
rect 22066 24228 22201 24256
rect 19521 24191 19579 24197
rect 19521 24188 19533 24191
rect 19392 24160 19533 24188
rect 19392 24148 19398 24160
rect 19521 24157 19533 24160
rect 19567 24157 19579 24191
rect 19521 24151 19579 24157
rect 19613 24191 19671 24197
rect 19613 24157 19625 24191
rect 19659 24157 19671 24191
rect 19613 24151 19671 24157
rect 19705 24191 19763 24197
rect 19705 24157 19717 24191
rect 19751 24157 19763 24191
rect 19705 24151 19763 24157
rect 19889 24191 19947 24197
rect 19889 24157 19901 24191
rect 19935 24188 19947 24191
rect 19978 24188 19984 24200
rect 19935 24160 19984 24188
rect 19935 24157 19947 24160
rect 19889 24151 19947 24157
rect 15580 24092 16712 24120
rect 16945 24123 17003 24129
rect 16945 24089 16957 24123
rect 16991 24120 17003 24123
rect 17402 24120 17408 24132
rect 16991 24092 17408 24120
rect 16991 24089 17003 24092
rect 16945 24083 17003 24089
rect 17402 24080 17408 24092
rect 17460 24080 17466 24132
rect 17494 24080 17500 24132
rect 17552 24120 17558 24132
rect 18049 24123 18107 24129
rect 17552 24092 17908 24120
rect 17552 24080 17558 24092
rect 9364 24024 10824 24052
rect 9364 24012 9370 24024
rect 12526 24012 12532 24064
rect 12584 24012 12590 24064
rect 13354 24012 13360 24064
rect 13412 24052 13418 24064
rect 14369 24055 14427 24061
rect 14369 24052 14381 24055
rect 13412 24024 14381 24052
rect 13412 24012 13418 24024
rect 14369 24021 14381 24024
rect 14415 24052 14427 24055
rect 16574 24052 16580 24064
rect 14415 24024 16580 24052
rect 14415 24021 14427 24024
rect 14369 24015 14427 24021
rect 16574 24012 16580 24024
rect 16632 24012 16638 24064
rect 17313 24055 17371 24061
rect 17313 24021 17325 24055
rect 17359 24052 17371 24055
rect 17770 24052 17776 24064
rect 17359 24024 17776 24052
rect 17359 24021 17371 24024
rect 17313 24015 17371 24021
rect 17770 24012 17776 24024
rect 17828 24012 17834 24064
rect 17880 24052 17908 24092
rect 18049 24089 18061 24123
rect 18095 24120 18107 24123
rect 18138 24120 18144 24132
rect 18095 24092 18144 24120
rect 18095 24089 18107 24092
rect 18049 24083 18107 24089
rect 18138 24080 18144 24092
rect 18196 24080 18202 24132
rect 19628 24120 19656 24151
rect 19978 24148 19984 24160
rect 20036 24148 20042 24200
rect 22066 24188 22094 24228
rect 22189 24225 22201 24228
rect 22235 24256 22247 24259
rect 22235 24228 27752 24256
rect 22235 24225 22247 24228
rect 22189 24219 22247 24225
rect 20456 24160 22094 24188
rect 20346 24120 20352 24132
rect 19628 24092 20352 24120
rect 20346 24080 20352 24092
rect 20404 24080 20410 24132
rect 20456 24052 20484 24160
rect 22370 24148 22376 24200
rect 22428 24188 22434 24200
rect 22649 24191 22707 24197
rect 22649 24188 22661 24191
rect 22428 24160 22661 24188
rect 22428 24148 22434 24160
rect 22649 24157 22661 24160
rect 22695 24157 22707 24191
rect 22649 24151 22707 24157
rect 23290 24148 23296 24200
rect 23348 24188 23354 24200
rect 27724 24197 27752 24228
rect 23569 24191 23627 24197
rect 23569 24188 23581 24191
rect 23348 24160 23581 24188
rect 23348 24148 23354 24160
rect 23569 24157 23581 24160
rect 23615 24157 23627 24191
rect 23569 24151 23627 24157
rect 27709 24191 27767 24197
rect 27709 24157 27721 24191
rect 27755 24157 27767 24191
rect 27709 24151 27767 24157
rect 27798 24148 27804 24200
rect 27856 24188 27862 24200
rect 28000 24197 28028 24296
rect 27893 24191 27951 24197
rect 27893 24188 27905 24191
rect 27856 24160 27905 24188
rect 27856 24148 27862 24160
rect 27893 24157 27905 24160
rect 27939 24157 27951 24191
rect 27893 24151 27951 24157
rect 27985 24191 28043 24197
rect 27985 24157 27997 24191
rect 28031 24157 28043 24191
rect 27985 24151 28043 24157
rect 28077 24191 28135 24197
rect 28077 24157 28089 24191
rect 28123 24188 28135 24191
rect 28994 24188 29000 24200
rect 28123 24160 29000 24188
rect 28123 24157 28135 24160
rect 28077 24151 28135 24157
rect 20533 24123 20591 24129
rect 20533 24089 20545 24123
rect 20579 24120 20591 24123
rect 21085 24123 21143 24129
rect 21085 24120 21097 24123
rect 20579 24092 21097 24120
rect 20579 24089 20591 24092
rect 20533 24083 20591 24089
rect 21085 24089 21097 24092
rect 21131 24120 21143 24123
rect 21910 24120 21916 24132
rect 21131 24092 21916 24120
rect 21131 24089 21143 24092
rect 21085 24083 21143 24089
rect 21910 24080 21916 24092
rect 21968 24080 21974 24132
rect 22005 24123 22063 24129
rect 22005 24089 22017 24123
rect 22051 24089 22063 24123
rect 22005 24083 22063 24089
rect 17880 24024 20484 24052
rect 21818 24012 21824 24064
rect 21876 24052 21882 24064
rect 22020 24052 22048 24083
rect 23198 24080 23204 24132
rect 23256 24120 23262 24132
rect 23385 24123 23443 24129
rect 23385 24120 23397 24123
rect 23256 24092 23397 24120
rect 23256 24080 23262 24092
rect 23385 24089 23397 24092
rect 23431 24089 23443 24123
rect 23385 24083 23443 24089
rect 23750 24080 23756 24132
rect 23808 24120 23814 24132
rect 25501 24123 25559 24129
rect 23808 24092 25452 24120
rect 23808 24080 23814 24092
rect 21876 24024 22048 24052
rect 22833 24055 22891 24061
rect 21876 24012 21882 24024
rect 22833 24021 22845 24055
rect 22879 24052 22891 24055
rect 23216 24052 23244 24080
rect 22879 24024 23244 24052
rect 24765 24055 24823 24061
rect 22879 24021 22891 24024
rect 22833 24015 22891 24021
rect 24765 24021 24777 24055
rect 24811 24052 24823 24055
rect 24854 24052 24860 24064
rect 24811 24024 24860 24052
rect 24811 24021 24823 24024
rect 24765 24015 24823 24021
rect 24854 24012 24860 24024
rect 24912 24012 24918 24064
rect 25424 24052 25452 24092
rect 25501 24089 25513 24123
rect 25547 24120 25559 24123
rect 27246 24120 27252 24132
rect 25547 24092 27252 24120
rect 25547 24089 25559 24092
rect 25501 24083 25559 24089
rect 27246 24080 27252 24092
rect 27304 24080 27310 24132
rect 28092 24052 28120 24151
rect 28994 24148 29000 24160
rect 29052 24148 29058 24200
rect 29454 24148 29460 24200
rect 29512 24188 29518 24200
rect 31113 24191 31171 24197
rect 31113 24188 31125 24191
rect 29512 24160 31125 24188
rect 29512 24148 29518 24160
rect 31113 24157 31125 24160
rect 31159 24157 31171 24191
rect 31276 24191 31334 24197
rect 31276 24188 31288 24191
rect 31113 24151 31171 24157
rect 31220 24160 31288 24188
rect 31220 24064 31248 24160
rect 31276 24157 31288 24160
rect 31322 24157 31334 24191
rect 31276 24151 31334 24157
rect 31386 24148 31392 24200
rect 31444 24188 31450 24200
rect 31542 24197 31570 24364
rect 31527 24191 31585 24197
rect 31444 24160 31489 24188
rect 31444 24148 31450 24160
rect 31527 24157 31539 24191
rect 31573 24157 31585 24191
rect 33962 24188 33968 24200
rect 33923 24160 33968 24188
rect 31527 24151 31585 24157
rect 33962 24148 33968 24160
rect 34020 24148 34026 24200
rect 68094 24188 68100 24200
rect 68055 24160 68100 24188
rect 68094 24148 68100 24160
rect 68152 24148 68158 24200
rect 31757 24123 31815 24129
rect 31757 24089 31769 24123
rect 31803 24120 31815 24123
rect 33698 24123 33756 24129
rect 33698 24120 33710 24123
rect 31803 24092 33710 24120
rect 31803 24089 31815 24092
rect 31757 24083 31815 24089
rect 33698 24089 33710 24092
rect 33744 24089 33756 24123
rect 33698 24083 33756 24089
rect 28350 24052 28356 24064
rect 25424 24024 28120 24052
rect 28311 24024 28356 24052
rect 28350 24012 28356 24024
rect 28408 24012 28414 24064
rect 31202 24012 31208 24064
rect 31260 24012 31266 24064
rect 32582 24052 32588 24064
rect 32543 24024 32588 24052
rect 32582 24012 32588 24024
rect 32640 24012 32646 24064
rect 1104 23962 68816 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 68816 23962
rect 1104 23888 68816 23910
rect 3697 23851 3755 23857
rect 3697 23817 3709 23851
rect 3743 23848 3755 23851
rect 4062 23848 4068 23860
rect 3743 23820 4068 23848
rect 3743 23817 3755 23820
rect 3697 23811 3755 23817
rect 4062 23808 4068 23820
rect 4120 23808 4126 23860
rect 5350 23808 5356 23860
rect 5408 23848 5414 23860
rect 5445 23851 5503 23857
rect 5445 23848 5457 23851
rect 5408 23820 5457 23848
rect 5408 23808 5414 23820
rect 5445 23817 5457 23820
rect 5491 23817 5503 23851
rect 8570 23848 8576 23860
rect 5445 23811 5503 23817
rect 8496 23820 8576 23848
rect 4249 23783 4307 23789
rect 4249 23749 4261 23783
rect 4295 23780 4307 23783
rect 5534 23780 5540 23792
rect 4295 23752 5540 23780
rect 4295 23749 4307 23752
rect 4249 23743 4307 23749
rect 3053 23715 3111 23721
rect 3053 23712 3065 23715
rect 2332 23684 3065 23712
rect 2332 23656 2360 23684
rect 3053 23681 3065 23684
rect 3099 23681 3111 23715
rect 3234 23712 3240 23724
rect 3195 23684 3240 23712
rect 3053 23675 3111 23681
rect 3234 23672 3240 23684
rect 3292 23672 3298 23724
rect 3326 23672 3332 23724
rect 3384 23712 3390 23724
rect 3467 23715 3525 23721
rect 3384 23684 3429 23712
rect 3384 23672 3390 23684
rect 3467 23681 3479 23715
rect 3513 23712 3525 23715
rect 4264 23712 4292 23743
rect 5534 23740 5540 23752
rect 5592 23740 5598 23792
rect 6822 23780 6828 23792
rect 6196 23752 6828 23780
rect 3513 23684 4292 23712
rect 5629 23715 5687 23721
rect 3513 23681 3525 23684
rect 3467 23675 3525 23681
rect 5629 23681 5641 23715
rect 5675 23712 5687 23715
rect 5718 23712 5724 23724
rect 5675 23684 5724 23712
rect 5675 23681 5687 23684
rect 5629 23675 5687 23681
rect 5718 23672 5724 23684
rect 5776 23712 5782 23724
rect 6196 23712 6224 23752
rect 6822 23740 6828 23752
rect 6880 23780 6886 23792
rect 7926 23780 7932 23792
rect 6880 23752 7932 23780
rect 6880 23740 6886 23752
rect 7926 23740 7932 23752
rect 7984 23740 7990 23792
rect 8496 23780 8524 23820
rect 8570 23808 8576 23820
rect 8628 23808 8634 23860
rect 8846 23848 8852 23860
rect 8807 23820 8852 23848
rect 8846 23808 8852 23820
rect 8904 23808 8910 23860
rect 9309 23851 9367 23857
rect 9309 23848 9321 23851
rect 8956 23820 9321 23848
rect 8956 23780 8984 23820
rect 9309 23817 9321 23820
rect 9355 23817 9367 23851
rect 9309 23811 9367 23817
rect 9858 23808 9864 23860
rect 9916 23848 9922 23860
rect 12894 23848 12900 23860
rect 9916 23820 12900 23848
rect 9916 23808 9922 23820
rect 12894 23808 12900 23820
rect 12952 23808 12958 23860
rect 15010 23808 15016 23860
rect 15068 23808 15074 23860
rect 15470 23848 15476 23860
rect 15431 23820 15476 23848
rect 15470 23808 15476 23820
rect 15528 23808 15534 23860
rect 15562 23808 15568 23860
rect 15620 23848 15626 23860
rect 15620 23820 17540 23848
rect 15620 23808 15626 23820
rect 13354 23780 13360 23792
rect 8023 23752 8524 23780
rect 6914 23712 6920 23724
rect 5776 23684 6224 23712
rect 6827 23684 6920 23712
rect 5776 23672 5782 23684
rect 6914 23672 6920 23684
rect 6972 23712 6978 23724
rect 7282 23712 7288 23724
rect 6972 23684 7288 23712
rect 6972 23672 6978 23684
rect 7282 23672 7288 23684
rect 7340 23672 7346 23724
rect 7374 23672 7380 23724
rect 7432 23712 7438 23724
rect 8023 23712 8051 23752
rect 7432 23684 8051 23712
rect 8205 23715 8263 23721
rect 7432 23672 7438 23684
rect 8205 23681 8217 23715
rect 8251 23681 8263 23715
rect 8205 23675 8263 23681
rect 2314 23644 2320 23656
rect 2275 23616 2320 23644
rect 2314 23604 2320 23616
rect 2372 23604 2378 23656
rect 2593 23647 2651 23653
rect 2593 23613 2605 23647
rect 2639 23644 2651 23647
rect 2774 23644 2780 23656
rect 2639 23616 2780 23644
rect 2639 23613 2651 23616
rect 2593 23607 2651 23613
rect 2774 23604 2780 23616
rect 2832 23604 2838 23656
rect 4985 23647 5043 23653
rect 4985 23613 4997 23647
rect 5031 23644 5043 23647
rect 5813 23647 5871 23653
rect 5813 23644 5825 23647
rect 5031 23616 5825 23644
rect 5031 23613 5043 23616
rect 4985 23607 5043 23613
rect 5813 23613 5825 23616
rect 5859 23644 5871 23647
rect 6454 23644 6460 23656
rect 5859 23616 6460 23644
rect 5859 23613 5871 23616
rect 5813 23607 5871 23613
rect 6454 23604 6460 23616
rect 6512 23604 6518 23656
rect 7193 23647 7251 23653
rect 7193 23613 7205 23647
rect 7239 23644 7251 23647
rect 7392 23644 7420 23672
rect 7239 23616 7420 23644
rect 7239 23613 7251 23616
rect 7193 23607 7251 23613
rect 8018 23604 8024 23656
rect 8076 23644 8082 23656
rect 8220 23644 8248 23675
rect 8294 23672 8300 23724
rect 8352 23712 8358 23724
rect 8496 23721 8524 23752
rect 8588 23752 8984 23780
rect 9048 23752 13360 23780
rect 8588 23721 8616 23752
rect 8389 23715 8447 23721
rect 8389 23712 8401 23715
rect 8352 23684 8401 23712
rect 8352 23672 8358 23684
rect 8389 23681 8401 23684
rect 8435 23681 8447 23715
rect 8389 23675 8447 23681
rect 8481 23715 8539 23721
rect 8481 23681 8493 23715
rect 8527 23681 8539 23715
rect 8481 23675 8539 23681
rect 8573 23715 8631 23721
rect 8573 23681 8585 23715
rect 8619 23710 8631 23715
rect 8619 23682 8708 23710
rect 8619 23681 8631 23682
rect 8573 23675 8631 23681
rect 8076 23616 8248 23644
rect 8076 23604 8082 23616
rect 3694 23536 3700 23588
rect 3752 23576 3758 23588
rect 6365 23579 6423 23585
rect 6365 23576 6377 23579
rect 3752 23548 6377 23576
rect 3752 23536 3758 23548
rect 6365 23545 6377 23548
rect 6411 23576 6423 23579
rect 7006 23576 7012 23588
rect 6411 23548 7012 23576
rect 6411 23545 6423 23548
rect 6365 23539 6423 23545
rect 7006 23536 7012 23548
rect 7064 23536 7070 23588
rect 8680 23576 8708 23682
rect 7852 23548 8708 23576
rect 3878 23468 3884 23520
rect 3936 23508 3942 23520
rect 7852 23508 7880 23548
rect 3936 23480 7880 23508
rect 3936 23468 3942 23480
rect 7926 23468 7932 23520
rect 7984 23508 7990 23520
rect 9048 23508 9076 23752
rect 13354 23740 13360 23752
rect 13412 23740 13418 23792
rect 15028 23780 15056 23808
rect 17512 23789 17540 23820
rect 18598 23808 18604 23860
rect 18656 23848 18662 23860
rect 20438 23848 20444 23860
rect 18656 23820 20444 23848
rect 18656 23808 18662 23820
rect 20438 23808 20444 23820
rect 20496 23808 20502 23860
rect 27341 23851 27399 23857
rect 27341 23817 27353 23851
rect 27387 23848 27399 23851
rect 27798 23848 27804 23860
rect 27387 23820 27804 23848
rect 27387 23817 27399 23820
rect 27341 23811 27399 23817
rect 27798 23808 27804 23820
rect 27856 23808 27862 23860
rect 27893 23851 27951 23857
rect 27893 23817 27905 23851
rect 27939 23848 27951 23851
rect 29086 23848 29092 23860
rect 27939 23820 29092 23848
rect 27939 23817 27951 23820
rect 27893 23811 27951 23817
rect 17497 23783 17555 23789
rect 13648 23752 15148 23780
rect 12437 23715 12495 23721
rect 12437 23681 12449 23715
rect 12483 23712 12495 23715
rect 12526 23712 12532 23724
rect 12483 23684 12532 23712
rect 12483 23681 12495 23684
rect 12437 23675 12495 23681
rect 12526 23672 12532 23684
rect 12584 23672 12590 23724
rect 12621 23715 12679 23721
rect 12621 23681 12633 23715
rect 12667 23712 12679 23715
rect 12986 23712 12992 23724
rect 12667 23684 12992 23712
rect 12667 23681 12679 23684
rect 12621 23675 12679 23681
rect 12986 23672 12992 23684
rect 13044 23672 13050 23724
rect 13538 23712 13544 23724
rect 13499 23684 13544 23712
rect 13538 23672 13544 23684
rect 13596 23672 13602 23724
rect 13648 23721 13676 23752
rect 13633 23715 13691 23721
rect 13633 23681 13645 23715
rect 13679 23681 13691 23715
rect 13633 23675 13691 23681
rect 13725 23715 13783 23721
rect 13725 23681 13737 23715
rect 13771 23681 13783 23715
rect 13725 23675 13783 23681
rect 12805 23647 12863 23653
rect 12805 23613 12817 23647
rect 12851 23644 12863 23647
rect 13740 23644 13768 23675
rect 13906 23672 13912 23724
rect 13964 23712 13970 23724
rect 14829 23715 14887 23721
rect 14829 23712 14841 23715
rect 13964 23684 14841 23712
rect 13964 23672 13970 23684
rect 14829 23681 14841 23684
rect 14875 23681 14887 23715
rect 15010 23712 15016 23724
rect 14971 23684 15016 23712
rect 14829 23675 14887 23681
rect 12851 23616 13768 23644
rect 12851 23613 12863 23616
rect 12805 23607 12863 23613
rect 14844 23576 14872 23675
rect 15010 23672 15016 23684
rect 15068 23672 15074 23724
rect 15120 23721 15148 23752
rect 17497 23749 17509 23783
rect 17543 23749 17555 23783
rect 17497 23743 17555 23749
rect 18322 23740 18328 23792
rect 18380 23780 18386 23792
rect 19429 23783 19487 23789
rect 19429 23780 19441 23783
rect 18380 23752 19441 23780
rect 18380 23740 18386 23752
rect 19429 23749 19441 23752
rect 19475 23780 19487 23783
rect 21910 23780 21916 23792
rect 19475 23752 21916 23780
rect 19475 23749 19487 23752
rect 19429 23743 19487 23749
rect 21910 23740 21916 23752
rect 21968 23740 21974 23792
rect 25590 23740 25596 23792
rect 25648 23780 25654 23792
rect 27157 23783 27215 23789
rect 27157 23780 27169 23783
rect 25648 23752 27169 23780
rect 25648 23740 25654 23752
rect 27157 23749 27169 23752
rect 27203 23749 27215 23783
rect 27157 23743 27215 23749
rect 27246 23740 27252 23792
rect 27304 23780 27310 23792
rect 27908 23780 27936 23811
rect 29086 23808 29092 23820
rect 29144 23848 29150 23860
rect 29270 23848 29276 23860
rect 29144 23820 29276 23848
rect 29144 23808 29150 23820
rect 29270 23808 29276 23820
rect 29328 23808 29334 23860
rect 31202 23808 31208 23860
rect 31260 23848 31266 23860
rect 31297 23851 31355 23857
rect 31297 23848 31309 23851
rect 31260 23820 31309 23848
rect 31260 23808 31266 23820
rect 31297 23817 31309 23820
rect 31343 23817 31355 23851
rect 31297 23811 31355 23817
rect 28810 23789 28816 23792
rect 28804 23780 28816 23789
rect 27304 23752 27936 23780
rect 28771 23752 28816 23780
rect 27304 23740 27310 23752
rect 28804 23743 28816 23752
rect 28810 23740 28816 23743
rect 28868 23740 28874 23792
rect 15105 23715 15163 23721
rect 15105 23681 15117 23715
rect 15151 23681 15163 23715
rect 15105 23675 15163 23681
rect 15197 23715 15255 23721
rect 15197 23681 15209 23715
rect 15243 23681 15255 23715
rect 15197 23675 15255 23681
rect 15212 23644 15240 23675
rect 15654 23672 15660 23724
rect 15712 23712 15718 23724
rect 17310 23721 17316 23724
rect 17129 23715 17187 23721
rect 17129 23712 17141 23715
rect 15712 23684 17141 23712
rect 15712 23672 15718 23684
rect 17129 23681 17141 23684
rect 17175 23681 17187 23715
rect 17129 23675 17187 23681
rect 17277 23715 17316 23721
rect 17277 23681 17289 23715
rect 17277 23675 17316 23681
rect 17310 23672 17316 23675
rect 17368 23672 17374 23724
rect 17402 23672 17408 23724
rect 17460 23712 17466 23724
rect 17460 23684 17505 23712
rect 17460 23672 17466 23684
rect 17586 23672 17592 23724
rect 17644 23721 17650 23724
rect 17644 23712 17652 23721
rect 17644 23684 17689 23712
rect 17644 23675 17652 23684
rect 17644 23672 17650 23675
rect 18138 23672 18144 23724
rect 18196 23712 18202 23724
rect 19245 23715 19303 23721
rect 19245 23712 19257 23715
rect 18196 23684 19257 23712
rect 18196 23672 18202 23684
rect 19245 23681 19257 23684
rect 19291 23681 19303 23715
rect 21818 23712 21824 23724
rect 19245 23675 19303 23681
rect 21192 23684 21824 23712
rect 16025 23647 16083 23653
rect 16025 23644 16037 23647
rect 15212 23616 16037 23644
rect 16025 23613 16037 23616
rect 16071 23644 16083 23647
rect 16206 23644 16212 23656
rect 16071 23616 16212 23644
rect 16071 23613 16083 23616
rect 16025 23607 16083 23613
rect 16206 23604 16212 23616
rect 16264 23644 16270 23656
rect 18785 23647 18843 23653
rect 18785 23644 18797 23647
rect 16264 23616 18797 23644
rect 16264 23604 16270 23616
rect 18785 23613 18797 23616
rect 18831 23644 18843 23647
rect 19334 23644 19340 23656
rect 18831 23616 19340 23644
rect 18831 23613 18843 23616
rect 18785 23607 18843 23613
rect 19334 23604 19340 23616
rect 19392 23604 19398 23656
rect 19610 23644 19616 23656
rect 19571 23616 19616 23644
rect 19610 23604 19616 23616
rect 19668 23604 19674 23656
rect 17494 23576 17500 23588
rect 14844 23548 17500 23576
rect 17494 23536 17500 23548
rect 17552 23536 17558 23588
rect 17773 23579 17831 23585
rect 17773 23545 17785 23579
rect 17819 23576 17831 23579
rect 19242 23576 19248 23588
rect 17819 23548 19248 23576
rect 17819 23545 17831 23548
rect 17773 23539 17831 23545
rect 19242 23536 19248 23548
rect 19300 23536 19306 23588
rect 21192 23585 21220 23684
rect 21818 23672 21824 23684
rect 21876 23712 21882 23724
rect 22097 23715 22155 23721
rect 22097 23712 22109 23715
rect 21876 23684 22109 23712
rect 21876 23672 21882 23684
rect 22097 23681 22109 23684
rect 22143 23681 22155 23715
rect 22097 23675 22155 23681
rect 23106 23672 23112 23724
rect 23164 23712 23170 23724
rect 23569 23715 23627 23721
rect 23569 23712 23581 23715
rect 23164 23684 23581 23712
rect 23164 23672 23170 23684
rect 23569 23681 23581 23684
rect 23615 23681 23627 23715
rect 24578 23712 24584 23724
rect 24539 23684 24584 23712
rect 23569 23675 23627 23681
rect 24578 23672 24584 23684
rect 24636 23672 24642 23724
rect 26878 23672 26884 23724
rect 26936 23712 26942 23724
rect 26973 23715 27031 23721
rect 26973 23712 26985 23715
rect 26936 23684 26985 23712
rect 26936 23672 26942 23684
rect 26973 23681 26985 23684
rect 27019 23681 27031 23715
rect 26973 23675 27031 23681
rect 30929 23715 30987 23721
rect 30929 23681 30941 23715
rect 30975 23712 30987 23715
rect 31018 23712 31024 23724
rect 30975 23684 31024 23712
rect 30975 23681 30987 23684
rect 30929 23675 30987 23681
rect 31018 23672 31024 23684
rect 31076 23672 31082 23724
rect 31113 23715 31171 23721
rect 31113 23681 31125 23715
rect 31159 23712 31171 23715
rect 31294 23712 31300 23724
rect 31159 23684 31300 23712
rect 31159 23681 31171 23684
rect 31113 23675 31171 23681
rect 31294 23672 31300 23684
rect 31352 23712 31358 23724
rect 32582 23712 32588 23724
rect 31352 23684 32588 23712
rect 31352 23672 31358 23684
rect 32582 23672 32588 23684
rect 32640 23672 32646 23724
rect 23293 23647 23351 23653
rect 23293 23613 23305 23647
rect 23339 23644 23351 23647
rect 23658 23644 23664 23656
rect 23339 23616 23664 23644
rect 23339 23613 23351 23616
rect 23293 23607 23351 23613
rect 23658 23604 23664 23616
rect 23716 23604 23722 23656
rect 24857 23647 24915 23653
rect 24857 23613 24869 23647
rect 24903 23644 24915 23647
rect 24946 23644 24952 23656
rect 24903 23616 24952 23644
rect 24903 23613 24915 23616
rect 24857 23607 24915 23613
rect 24946 23604 24952 23616
rect 25004 23604 25010 23656
rect 25317 23647 25375 23653
rect 25317 23613 25329 23647
rect 25363 23613 25375 23647
rect 25317 23607 25375 23613
rect 25593 23647 25651 23653
rect 25593 23613 25605 23647
rect 25639 23644 25651 23647
rect 26142 23644 26148 23656
rect 25639 23616 26148 23644
rect 25639 23613 25651 23616
rect 25593 23607 25651 23613
rect 21177 23579 21235 23585
rect 21177 23576 21189 23579
rect 19536 23548 21189 23576
rect 13262 23508 13268 23520
rect 7984 23480 9076 23508
rect 13223 23480 13268 23508
rect 7984 23468 7990 23480
rect 13262 23468 13268 23480
rect 13320 23468 13326 23520
rect 17218 23468 17224 23520
rect 17276 23508 17282 23520
rect 19536 23508 19564 23548
rect 21177 23545 21189 23548
rect 21223 23545 21235 23579
rect 21177 23539 21235 23545
rect 22738 23536 22744 23588
rect 22796 23576 22802 23588
rect 25332 23576 25360 23607
rect 26142 23604 26148 23616
rect 26200 23604 26206 23656
rect 28537 23647 28595 23653
rect 28537 23644 28549 23647
rect 26988 23616 28549 23644
rect 26988 23588 27016 23616
rect 28537 23613 28549 23616
rect 28583 23613 28595 23647
rect 28537 23607 28595 23613
rect 22796 23548 25360 23576
rect 22796 23536 22802 23548
rect 26970 23536 26976 23588
rect 27028 23536 27034 23588
rect 29472 23548 30512 23576
rect 17276 23480 19564 23508
rect 17276 23468 17282 23480
rect 22094 23468 22100 23520
rect 22152 23508 22158 23520
rect 22189 23511 22247 23517
rect 22189 23508 22201 23511
rect 22152 23480 22201 23508
rect 22152 23468 22158 23480
rect 22189 23477 22201 23480
rect 22235 23508 22247 23511
rect 25406 23508 25412 23520
rect 22235 23480 25412 23508
rect 22235 23477 22247 23480
rect 22189 23471 22247 23477
rect 25406 23468 25412 23480
rect 25464 23468 25470 23520
rect 26326 23468 26332 23520
rect 26384 23508 26390 23520
rect 29472 23508 29500 23548
rect 26384 23480 29500 23508
rect 29917 23511 29975 23517
rect 26384 23468 26390 23480
rect 29917 23477 29929 23511
rect 29963 23508 29975 23511
rect 30006 23508 30012 23520
rect 29963 23480 30012 23508
rect 29963 23477 29975 23480
rect 29917 23471 29975 23477
rect 30006 23468 30012 23480
rect 30064 23468 30070 23520
rect 30484 23517 30512 23548
rect 30469 23511 30527 23517
rect 30469 23477 30481 23511
rect 30515 23508 30527 23511
rect 30650 23508 30656 23520
rect 30515 23480 30656 23508
rect 30515 23477 30527 23480
rect 30469 23471 30527 23477
rect 30650 23468 30656 23480
rect 30708 23468 30714 23520
rect 1104 23418 68816 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 65654 23418
rect 65706 23366 65718 23418
rect 65770 23366 65782 23418
rect 65834 23366 65846 23418
rect 65898 23366 65910 23418
rect 65962 23366 68816 23418
rect 1104 23344 68816 23366
rect 1673 23307 1731 23313
rect 1673 23273 1685 23307
rect 1719 23304 1731 23307
rect 2406 23304 2412 23316
rect 1719 23276 2412 23304
rect 1719 23273 1731 23276
rect 1673 23267 1731 23273
rect 2406 23264 2412 23276
rect 2464 23304 2470 23316
rect 2590 23304 2596 23316
rect 2464 23276 2596 23304
rect 2464 23264 2470 23276
rect 2590 23264 2596 23276
rect 2648 23264 2654 23316
rect 6641 23307 6699 23313
rect 6641 23273 6653 23307
rect 6687 23304 6699 23307
rect 6914 23304 6920 23316
rect 6687 23276 6920 23304
rect 6687 23273 6699 23276
rect 6641 23267 6699 23273
rect 6914 23264 6920 23276
rect 6972 23264 6978 23316
rect 7193 23307 7251 23313
rect 7193 23273 7205 23307
rect 7239 23304 7251 23307
rect 8294 23304 8300 23316
rect 7239 23276 8300 23304
rect 7239 23273 7251 23276
rect 7193 23267 7251 23273
rect 8294 23264 8300 23276
rect 8352 23264 8358 23316
rect 8389 23307 8447 23313
rect 8389 23273 8401 23307
rect 8435 23304 8447 23307
rect 8662 23304 8668 23316
rect 8435 23276 8668 23304
rect 8435 23273 8447 23276
rect 8389 23267 8447 23273
rect 8662 23264 8668 23276
rect 8720 23264 8726 23316
rect 12986 23304 12992 23316
rect 12947 23276 12992 23304
rect 12986 23264 12992 23276
rect 13044 23264 13050 23316
rect 14645 23307 14703 23313
rect 14645 23273 14657 23307
rect 14691 23304 14703 23307
rect 15010 23304 15016 23316
rect 14691 23276 15016 23304
rect 14691 23273 14703 23276
rect 14645 23267 14703 23273
rect 15010 23264 15016 23276
rect 15068 23264 15074 23316
rect 15654 23304 15660 23316
rect 15615 23276 15660 23304
rect 15654 23264 15660 23276
rect 15712 23264 15718 23316
rect 15746 23264 15752 23316
rect 15804 23304 15810 23316
rect 21910 23304 21916 23316
rect 15804 23276 21496 23304
rect 21871 23276 21916 23304
rect 15804 23264 15810 23276
rect 5626 23236 5632 23248
rect 5587 23208 5632 23236
rect 5626 23196 5632 23208
rect 5684 23196 5690 23248
rect 13538 23236 13544 23248
rect 13451 23208 13544 23236
rect 13538 23196 13544 23208
rect 13596 23236 13602 23248
rect 17494 23236 17500 23248
rect 13596 23208 17500 23236
rect 13596 23196 13602 23208
rect 17494 23196 17500 23208
rect 17552 23196 17558 23248
rect 17586 23196 17592 23248
rect 17644 23196 17650 23248
rect 21468 23236 21496 23276
rect 21910 23264 21916 23276
rect 21968 23264 21974 23316
rect 25590 23304 25596 23316
rect 25551 23276 25596 23304
rect 25590 23264 25596 23276
rect 25648 23264 25654 23316
rect 23750 23236 23756 23248
rect 21468 23208 23756 23236
rect 1946 23128 1952 23180
rect 2004 23168 2010 23180
rect 3326 23168 3332 23180
rect 2004 23140 2452 23168
rect 2004 23128 2010 23140
rect 1854 23100 1860 23112
rect 1815 23072 1860 23100
rect 1854 23060 1860 23072
rect 1912 23060 1918 23112
rect 2314 23100 2320 23112
rect 2275 23072 2320 23100
rect 2314 23060 2320 23072
rect 2372 23060 2378 23112
rect 2424 23100 2452 23140
rect 2608 23140 3332 23168
rect 2608 23109 2636 23140
rect 3326 23128 3332 23140
rect 3384 23128 3390 23180
rect 9306 23168 9312 23180
rect 7392 23140 9312 23168
rect 2480 23103 2538 23109
rect 2480 23100 2492 23103
rect 2424 23072 2492 23100
rect 2480 23069 2492 23072
rect 2526 23069 2538 23103
rect 2480 23063 2538 23069
rect 2593 23103 2651 23109
rect 2593 23069 2605 23103
rect 2639 23069 2651 23103
rect 2593 23063 2651 23069
rect 2685 23103 2743 23109
rect 2685 23069 2697 23103
rect 2731 23069 2743 23103
rect 2685 23063 2743 23069
rect 2038 22992 2044 23044
rect 2096 23032 2102 23044
rect 2608 23032 2636 23063
rect 2096 23004 2636 23032
rect 2700 23032 2728 23063
rect 2866 23060 2872 23112
rect 2924 23100 2930 23112
rect 3789 23103 3847 23109
rect 3789 23100 3801 23103
rect 2924 23072 3801 23100
rect 2924 23060 2930 23072
rect 3789 23069 3801 23072
rect 3835 23069 3847 23103
rect 3789 23063 3847 23069
rect 6362 23060 6368 23112
rect 6420 23100 6426 23112
rect 6549 23103 6607 23109
rect 6549 23100 6561 23103
rect 6420 23072 6561 23100
rect 6420 23060 6426 23072
rect 6549 23069 6561 23072
rect 6595 23069 6607 23103
rect 6549 23063 6607 23069
rect 6733 23103 6791 23109
rect 6733 23069 6745 23103
rect 6779 23100 6791 23103
rect 7282 23100 7288 23112
rect 6779 23072 7288 23100
rect 6779 23069 6791 23072
rect 6733 23063 6791 23069
rect 7282 23060 7288 23072
rect 7340 23060 7346 23112
rect 7392 23109 7420 23140
rect 9306 23128 9312 23140
rect 9364 23128 9370 23180
rect 9398 23128 9404 23180
rect 9456 23168 9462 23180
rect 9769 23171 9827 23177
rect 9769 23168 9781 23171
rect 9456 23140 9781 23168
rect 9456 23128 9462 23140
rect 9769 23137 9781 23140
rect 9815 23137 9827 23171
rect 9769 23131 9827 23137
rect 14274 23128 14280 23180
rect 14332 23168 14338 23180
rect 17313 23171 17371 23177
rect 14332 23140 15516 23168
rect 14332 23128 14338 23140
rect 7377 23103 7435 23109
rect 7377 23069 7389 23103
rect 7423 23069 7435 23103
rect 7377 23063 7435 23069
rect 7561 23103 7619 23109
rect 7561 23069 7573 23103
rect 7607 23100 7619 23103
rect 8021 23103 8079 23109
rect 8021 23100 8033 23103
rect 7607 23072 8033 23100
rect 7607 23069 7619 23072
rect 7561 23063 7619 23069
rect 8021 23069 8033 23072
rect 8067 23100 8079 23103
rect 8938 23100 8944 23112
rect 8067 23072 8944 23100
rect 8067 23069 8079 23072
rect 8021 23063 8079 23069
rect 8938 23060 8944 23072
rect 8996 23060 9002 23112
rect 9030 23060 9036 23112
rect 9088 23060 9094 23112
rect 11609 23103 11667 23109
rect 11609 23069 11621 23103
rect 11655 23100 11667 23103
rect 12434 23100 12440 23112
rect 11655 23072 12440 23100
rect 11655 23069 11667 23072
rect 11609 23063 11667 23069
rect 12434 23060 12440 23072
rect 12492 23060 12498 23112
rect 13814 23060 13820 23112
rect 13872 23100 13878 23112
rect 14461 23103 14519 23109
rect 13872 23072 14412 23100
rect 13872 23060 13878 23072
rect 2961 23035 3019 23041
rect 2700 23004 2912 23032
rect 2096 22992 2102 23004
rect 2884 22964 2912 23004
rect 2961 23001 2973 23035
rect 3007 23032 3019 23035
rect 4034 23035 4092 23041
rect 4034 23032 4046 23035
rect 3007 23004 4046 23032
rect 3007 23001 3019 23004
rect 2961 22995 3019 23001
rect 4034 23001 4046 23004
rect 4080 23001 4092 23035
rect 4034 22995 4092 23001
rect 5813 23035 5871 23041
rect 5813 23001 5825 23035
rect 5859 23032 5871 23035
rect 6086 23032 6092 23044
rect 5859 23004 6092 23032
rect 5859 23001 5871 23004
rect 5813 22995 5871 23001
rect 6086 22992 6092 23004
rect 6144 22992 6150 23044
rect 8205 23035 8263 23041
rect 8205 23001 8217 23035
rect 8251 23032 8263 23035
rect 9048 23032 9076 23060
rect 8251 23004 9076 23032
rect 9125 23035 9183 23041
rect 8251 23001 8263 23004
rect 8205 22995 8263 23001
rect 9125 23001 9137 23035
rect 9171 23032 9183 23035
rect 9171 23004 9444 23032
rect 9171 23001 9183 23004
rect 9125 22995 9183 23001
rect 3050 22964 3056 22976
rect 2884 22936 3056 22964
rect 3050 22924 3056 22936
rect 3108 22964 3114 22976
rect 3878 22964 3884 22976
rect 3108 22936 3884 22964
rect 3108 22924 3114 22936
rect 3878 22924 3884 22936
rect 3936 22924 3942 22976
rect 5166 22964 5172 22976
rect 5127 22936 5172 22964
rect 5166 22924 5172 22936
rect 5224 22924 5230 22976
rect 9030 22924 9036 22976
rect 9088 22964 9094 22976
rect 9309 22967 9367 22973
rect 9309 22964 9321 22967
rect 9088 22936 9321 22964
rect 9088 22924 9094 22936
rect 9309 22933 9321 22936
rect 9355 22933 9367 22967
rect 9416 22964 9444 23004
rect 9490 22992 9496 23044
rect 9548 23032 9554 23044
rect 10014 23035 10072 23041
rect 10014 23032 10026 23035
rect 9548 23004 10026 23032
rect 9548 22992 9554 23004
rect 10014 23001 10026 23004
rect 10060 23001 10072 23035
rect 10014 22995 10072 23001
rect 11876 23035 11934 23041
rect 11876 23001 11888 23035
rect 11922 23032 11934 23035
rect 13262 23032 13268 23044
rect 11922 23004 13268 23032
rect 11922 23001 11934 23004
rect 11876 22995 11934 23001
rect 13262 22992 13268 23004
rect 13320 22992 13326 23044
rect 13372 23004 13584 23032
rect 11149 22967 11207 22973
rect 11149 22964 11161 22967
rect 9416 22936 11161 22964
rect 9309 22927 9367 22933
rect 11149 22933 11161 22936
rect 11195 22964 11207 22967
rect 13372 22964 13400 23004
rect 11195 22936 13400 22964
rect 13556 22964 13584 23004
rect 13906 22992 13912 23044
rect 13964 23032 13970 23044
rect 14277 23035 14335 23041
rect 14277 23032 14289 23035
rect 13964 23004 14289 23032
rect 13964 22992 13970 23004
rect 14277 23001 14289 23004
rect 14323 23001 14335 23035
rect 14384 23032 14412 23072
rect 14461 23069 14473 23103
rect 14507 23100 14519 23103
rect 14734 23100 14740 23112
rect 14507 23072 14740 23100
rect 14507 23069 14519 23072
rect 14461 23063 14519 23069
rect 14734 23060 14740 23072
rect 14792 23100 14798 23112
rect 15488 23109 15516 23140
rect 17313 23137 17325 23171
rect 17359 23168 17371 23171
rect 17604 23168 17632 23196
rect 17359 23140 17632 23168
rect 17359 23137 17371 23140
rect 17313 23131 17371 23137
rect 19334 23128 19340 23180
rect 19392 23168 19398 23180
rect 20346 23168 20352 23180
rect 19392 23140 20352 23168
rect 19392 23128 19398 23140
rect 15105 23103 15163 23109
rect 15105 23100 15117 23103
rect 14792 23072 15117 23100
rect 14792 23060 14798 23072
rect 15105 23069 15117 23072
rect 15151 23069 15163 23103
rect 15105 23063 15163 23069
rect 15473 23103 15531 23109
rect 15473 23069 15485 23103
rect 15519 23069 15531 23103
rect 17586 23100 17592 23112
rect 17547 23072 17592 23100
rect 15473 23063 15531 23069
rect 17586 23060 17592 23072
rect 17644 23060 17650 23112
rect 19426 23100 19432 23112
rect 19387 23072 19432 23100
rect 19426 23060 19432 23072
rect 19484 23060 19490 23112
rect 19610 23100 19616 23112
rect 19571 23072 19616 23100
rect 19610 23060 19616 23072
rect 19668 23060 19674 23112
rect 19720 23109 19748 23140
rect 20346 23128 20352 23140
rect 20404 23128 20410 23180
rect 19705 23103 19763 23109
rect 19705 23069 19717 23103
rect 19751 23069 19763 23103
rect 19705 23063 19763 23069
rect 19797 23103 19855 23109
rect 19797 23069 19809 23103
rect 19843 23069 19855 23103
rect 19797 23063 19855 23069
rect 14918 23032 14924 23044
rect 14384 23004 14924 23032
rect 14277 22995 14335 23001
rect 14918 22992 14924 23004
rect 14976 23032 14982 23044
rect 15289 23035 15347 23041
rect 15289 23032 15301 23035
rect 14976 23004 15301 23032
rect 14976 22992 14982 23004
rect 15120 22976 15148 23004
rect 15289 23001 15301 23004
rect 15335 23001 15347 23035
rect 15289 22995 15347 23001
rect 15378 22992 15384 23044
rect 15436 23032 15442 23044
rect 15436 23004 15481 23032
rect 15436 22992 15442 23004
rect 16022 22992 16028 23044
rect 16080 23032 16086 23044
rect 17034 23032 17040 23044
rect 16080 23004 17040 23032
rect 16080 22992 16086 23004
rect 17034 22992 17040 23004
rect 17092 23032 17098 23044
rect 18601 23035 18659 23041
rect 18601 23032 18613 23035
rect 17092 23004 18613 23032
rect 17092 22992 17098 23004
rect 18601 23001 18613 23004
rect 18647 23032 18659 23035
rect 19812 23032 19840 23063
rect 20070 23060 20076 23112
rect 20128 23100 20134 23112
rect 20533 23103 20591 23109
rect 20533 23100 20545 23103
rect 20128 23072 20545 23100
rect 20128 23060 20134 23072
rect 20533 23069 20545 23072
rect 20579 23100 20591 23103
rect 20622 23100 20628 23112
rect 20579 23072 20628 23100
rect 20579 23069 20591 23072
rect 20533 23063 20591 23069
rect 20622 23060 20628 23072
rect 20680 23060 20686 23112
rect 22646 23100 22652 23112
rect 22607 23072 22652 23100
rect 22646 23060 22652 23072
rect 22704 23060 22710 23112
rect 22830 23100 22836 23112
rect 22791 23072 22836 23100
rect 22830 23060 22836 23072
rect 22888 23060 22894 23112
rect 23032 23109 23060 23208
rect 23750 23196 23756 23208
rect 23808 23196 23814 23248
rect 26970 23168 26976 23180
rect 26931 23140 26976 23168
rect 26970 23128 26976 23140
rect 27028 23168 27034 23180
rect 27617 23171 27675 23177
rect 27617 23168 27629 23171
rect 27028 23140 27629 23168
rect 27028 23128 27034 23140
rect 27617 23137 27629 23140
rect 27663 23137 27675 23171
rect 29822 23168 29828 23180
rect 29735 23140 29828 23168
rect 27617 23131 27675 23137
rect 29822 23128 29828 23140
rect 29880 23168 29886 23180
rect 30466 23168 30472 23180
rect 29880 23140 30472 23168
rect 29880 23128 29886 23140
rect 30466 23128 30472 23140
rect 30524 23168 30530 23180
rect 31386 23168 31392 23180
rect 30524 23140 31392 23168
rect 30524 23128 30530 23140
rect 31386 23128 31392 23140
rect 31444 23128 31450 23180
rect 22925 23103 22983 23109
rect 22925 23069 22937 23103
rect 22971 23069 22983 23103
rect 22925 23063 22983 23069
rect 23017 23103 23075 23109
rect 23017 23069 23029 23103
rect 23063 23069 23075 23103
rect 23017 23063 23075 23069
rect 26717 23103 26775 23109
rect 26717 23069 26729 23103
rect 26763 23100 26775 23103
rect 28350 23100 28356 23112
rect 26763 23072 28356 23100
rect 26763 23069 26775 23072
rect 26717 23063 26775 23069
rect 20778 23035 20836 23041
rect 20778 23032 20790 23035
rect 18647 23004 19840 23032
rect 20088 23004 20790 23032
rect 18647 23001 18659 23004
rect 18601 22995 18659 23001
rect 15010 22964 15016 22976
rect 13556 22936 15016 22964
rect 11195 22933 11207 22936
rect 11149 22927 11207 22933
rect 15010 22924 15016 22936
rect 15068 22924 15074 22976
rect 15102 22924 15108 22976
rect 15160 22924 15166 22976
rect 15838 22924 15844 22976
rect 15896 22964 15902 22976
rect 20088 22973 20116 23004
rect 20778 23001 20790 23004
rect 20824 23001 20836 23035
rect 22940 23032 22968 23063
rect 28350 23060 28356 23072
rect 28408 23060 28414 23112
rect 28902 23060 28908 23112
rect 28960 23100 28966 23112
rect 29549 23103 29607 23109
rect 29549 23100 29561 23103
rect 28960 23072 29561 23100
rect 28960 23060 28966 23072
rect 29549 23069 29561 23072
rect 29595 23069 29607 23103
rect 29549 23063 29607 23069
rect 29914 23060 29920 23112
rect 29972 23100 29978 23112
rect 30837 23103 30895 23109
rect 30837 23100 30849 23103
rect 29972 23072 30849 23100
rect 29972 23060 29978 23072
rect 30837 23069 30849 23072
rect 30883 23069 30895 23103
rect 30837 23063 30895 23069
rect 30926 23060 30932 23112
rect 30984 23100 30990 23112
rect 31573 23103 31631 23109
rect 31573 23100 31585 23103
rect 30984 23072 31585 23100
rect 30984 23060 30990 23072
rect 31573 23069 31585 23072
rect 31619 23069 31631 23103
rect 31573 23063 31631 23069
rect 23106 23032 23112 23044
rect 22940 23004 23112 23032
rect 20778 22995 20836 23001
rect 23106 22992 23112 23004
rect 23164 22992 23170 23044
rect 27884 23035 27942 23041
rect 27884 23001 27896 23035
rect 27930 23032 27942 23035
rect 28074 23032 28080 23044
rect 27930 23004 28080 23032
rect 27930 23001 27942 23004
rect 27884 22995 27942 23001
rect 28074 22992 28080 23004
rect 28132 22992 28138 23044
rect 31110 22992 31116 23044
rect 31168 23032 31174 23044
rect 31818 23035 31876 23041
rect 31818 23032 31830 23035
rect 31168 23004 31830 23032
rect 31168 22992 31174 23004
rect 31818 23001 31830 23004
rect 31864 23001 31876 23035
rect 31818 22995 31876 23001
rect 16209 22967 16267 22973
rect 16209 22964 16221 22967
rect 15896 22936 16221 22964
rect 15896 22924 15902 22936
rect 16209 22933 16221 22936
rect 16255 22933 16267 22967
rect 16209 22927 16267 22933
rect 20073 22967 20131 22973
rect 20073 22933 20085 22967
rect 20119 22933 20131 22967
rect 23290 22964 23296 22976
rect 23251 22936 23296 22964
rect 20073 22927 20131 22933
rect 23290 22924 23296 22936
rect 23348 22924 23354 22976
rect 23750 22964 23756 22976
rect 23711 22936 23756 22964
rect 23750 22924 23756 22936
rect 23808 22924 23814 22976
rect 28994 22964 29000 22976
rect 28955 22936 29000 22964
rect 28994 22924 29000 22936
rect 29052 22924 29058 22976
rect 31018 22964 31024 22976
rect 30979 22936 31024 22964
rect 31018 22924 31024 22936
rect 31076 22924 31082 22976
rect 32950 22964 32956 22976
rect 32911 22936 32956 22964
rect 32950 22924 32956 22936
rect 33008 22924 33014 22976
rect 1104 22874 68816 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 68816 22874
rect 1104 22800 68816 22822
rect 2498 22720 2504 22772
rect 2556 22760 2562 22772
rect 9490 22760 9496 22772
rect 2556 22732 9240 22760
rect 9451 22732 9496 22760
rect 2556 22720 2562 22732
rect 2314 22692 2320 22704
rect 1780 22664 2320 22692
rect 1780 22633 1808 22664
rect 2314 22652 2320 22664
rect 2372 22652 2378 22704
rect 2409 22695 2467 22701
rect 2409 22661 2421 22695
rect 2455 22692 2467 22695
rect 3114 22695 3172 22701
rect 3114 22692 3126 22695
rect 2455 22664 3126 22692
rect 2455 22661 2467 22664
rect 2409 22655 2467 22661
rect 3114 22661 3126 22664
rect 3160 22661 3172 22695
rect 3114 22655 3172 22661
rect 3970 22652 3976 22704
rect 4028 22692 4034 22704
rect 4028 22664 5120 22692
rect 4028 22652 4034 22664
rect 1765 22627 1823 22633
rect 1765 22593 1777 22627
rect 1811 22593 1823 22627
rect 1946 22624 1952 22636
rect 1907 22596 1952 22624
rect 1765 22587 1823 22593
rect 1946 22584 1952 22596
rect 2004 22584 2010 22636
rect 2038 22584 2044 22636
rect 2096 22624 2102 22636
rect 2179 22627 2237 22633
rect 2096 22596 2141 22624
rect 2096 22584 2102 22596
rect 2179 22593 2191 22627
rect 2225 22624 2237 22627
rect 2498 22624 2504 22636
rect 2225 22596 2504 22624
rect 2225 22593 2237 22596
rect 2179 22587 2237 22593
rect 2498 22584 2504 22596
rect 2556 22584 2562 22636
rect 2866 22624 2872 22636
rect 2827 22596 2872 22624
rect 2866 22584 2872 22596
rect 2924 22584 2930 22636
rect 5092 22633 5120 22664
rect 6914 22652 6920 22704
rect 6972 22692 6978 22704
rect 8018 22692 8024 22704
rect 6972 22664 7236 22692
rect 6972 22652 6978 22664
rect 4985 22627 5043 22633
rect 4985 22593 4997 22627
rect 5031 22593 5043 22627
rect 4985 22587 5043 22593
rect 5077 22627 5135 22633
rect 5077 22593 5089 22627
rect 5123 22593 5135 22627
rect 5077 22587 5135 22593
rect 5000 22556 5028 22587
rect 5166 22584 5172 22636
rect 5224 22624 5230 22636
rect 5350 22624 5356 22636
rect 5224 22596 5269 22624
rect 5311 22596 5356 22624
rect 5224 22584 5230 22596
rect 5350 22584 5356 22596
rect 5408 22584 5414 22636
rect 7208 22633 7236 22664
rect 7484 22664 8024 22692
rect 7484 22633 7512 22664
rect 8018 22652 8024 22664
rect 8076 22692 8082 22704
rect 8478 22692 8484 22704
rect 8076 22664 8484 22692
rect 8076 22652 8082 22664
rect 8478 22652 8484 22664
rect 8536 22692 8542 22704
rect 8536 22664 8892 22692
rect 8536 22652 8542 22664
rect 8864 22636 8892 22664
rect 7101 22627 7159 22633
rect 7101 22593 7113 22627
rect 7147 22593 7159 22627
rect 7101 22587 7159 22593
rect 7193 22627 7251 22633
rect 7193 22593 7205 22627
rect 7239 22593 7251 22627
rect 7193 22587 7251 22593
rect 7285 22627 7343 22633
rect 7285 22593 7297 22627
rect 7331 22593 7343 22627
rect 7285 22587 7343 22593
rect 7469 22627 7527 22633
rect 7469 22593 7481 22627
rect 7515 22593 7527 22627
rect 8110 22624 8116 22636
rect 8071 22596 8116 22624
rect 7469 22587 7527 22593
rect 7116 22556 7144 22587
rect 5000 22528 7144 22556
rect 7300 22556 7328 22587
rect 8110 22584 8116 22596
rect 8168 22584 8174 22636
rect 8202 22584 8208 22636
rect 8260 22624 8266 22636
rect 8297 22627 8355 22633
rect 8297 22624 8309 22627
rect 8260 22596 8309 22624
rect 8260 22584 8266 22596
rect 8297 22593 8309 22596
rect 8343 22593 8355 22627
rect 8846 22624 8852 22636
rect 8807 22596 8852 22624
rect 8297 22587 8355 22593
rect 8846 22584 8852 22596
rect 8904 22584 8910 22636
rect 9030 22624 9036 22636
rect 8991 22596 9036 22624
rect 9030 22584 9036 22596
rect 9088 22584 9094 22636
rect 9212 22633 9240 22732
rect 9490 22720 9496 22732
rect 9548 22720 9554 22772
rect 14185 22763 14243 22769
rect 14185 22729 14197 22763
rect 14231 22729 14243 22763
rect 14185 22723 14243 22729
rect 13814 22692 13820 22704
rect 13775 22664 13820 22692
rect 13814 22652 13820 22664
rect 13872 22652 13878 22704
rect 13906 22652 13912 22704
rect 13964 22692 13970 22704
rect 13964 22664 14009 22692
rect 13964 22652 13970 22664
rect 9125 22627 9183 22633
rect 9125 22593 9137 22627
rect 9171 22593 9183 22627
rect 9212 22627 9275 22633
rect 9212 22596 9229 22627
rect 9125 22587 9183 22593
rect 9217 22593 9229 22596
rect 9263 22624 9275 22627
rect 9953 22627 10011 22633
rect 9953 22624 9965 22627
rect 9263 22596 9965 22624
rect 9263 22593 9275 22596
rect 9217 22587 9275 22593
rect 9953 22593 9965 22596
rect 9999 22593 10011 22627
rect 9953 22587 10011 22593
rect 7929 22559 7987 22565
rect 7929 22556 7941 22559
rect 7300 22528 7941 22556
rect 4249 22491 4307 22497
rect 4249 22457 4261 22491
rect 4295 22488 4307 22491
rect 4614 22488 4620 22500
rect 4295 22460 4620 22488
rect 4295 22457 4307 22460
rect 4249 22451 4307 22457
rect 4614 22448 4620 22460
rect 4672 22448 4678 22500
rect 7116 22488 7144 22528
rect 7929 22525 7941 22528
rect 7975 22525 7987 22559
rect 7929 22519 7987 22525
rect 7374 22488 7380 22500
rect 7116 22460 7380 22488
rect 7374 22448 7380 22460
rect 7432 22448 7438 22500
rect 7466 22448 7472 22500
rect 7524 22488 7530 22500
rect 8220 22488 8248 22584
rect 8570 22516 8576 22568
rect 8628 22556 8634 22568
rect 9140 22556 9168 22587
rect 12986 22584 12992 22636
rect 13044 22624 13050 22636
rect 13633 22627 13691 22633
rect 13633 22624 13645 22627
rect 13044 22596 13645 22624
rect 13044 22584 13050 22596
rect 13633 22593 13645 22596
rect 13679 22593 13691 22627
rect 13633 22587 13691 22593
rect 14001 22627 14059 22633
rect 14001 22593 14013 22627
rect 14047 22593 14059 22627
rect 14200 22624 14228 22723
rect 22646 22720 22652 22772
rect 22704 22760 22710 22772
rect 26145 22763 26203 22769
rect 26145 22760 26157 22763
rect 22704 22732 26157 22760
rect 22704 22720 22710 22732
rect 26145 22729 26157 22732
rect 26191 22729 26203 22763
rect 28074 22760 28080 22772
rect 28035 22732 28080 22760
rect 26145 22723 26203 22729
rect 15010 22692 15016 22704
rect 14971 22664 15016 22692
rect 15010 22652 15016 22664
rect 15068 22652 15074 22704
rect 17804 22695 17862 22701
rect 17804 22661 17816 22695
rect 17850 22692 17862 22695
rect 18601 22695 18659 22701
rect 18601 22692 18613 22695
rect 17850 22664 18613 22692
rect 17850 22661 17862 22664
rect 17804 22655 17862 22661
rect 18601 22661 18613 22664
rect 18647 22661 18659 22695
rect 19334 22692 19340 22704
rect 18601 22655 18659 22661
rect 18984 22664 19340 22692
rect 14645 22627 14703 22633
rect 14645 22624 14657 22627
rect 14200 22596 14657 22624
rect 14001 22587 14059 22593
rect 14645 22593 14657 22596
rect 14691 22593 14703 22627
rect 14645 22587 14703 22593
rect 14738 22627 14796 22633
rect 14738 22593 14750 22627
rect 14784 22593 14796 22627
rect 14918 22624 14924 22636
rect 14879 22596 14924 22624
rect 14738 22587 14796 22593
rect 8628 22528 9168 22556
rect 14016 22556 14044 22587
rect 14274 22556 14280 22568
rect 14016 22528 14280 22556
rect 8628 22516 8634 22528
rect 14274 22516 14280 22528
rect 14332 22516 14338 22568
rect 14752 22556 14780 22587
rect 14918 22584 14924 22596
rect 14976 22584 14982 22636
rect 15151 22627 15209 22633
rect 15151 22593 15163 22627
rect 15197 22624 15209 22627
rect 15838 22624 15844 22636
rect 15197 22596 15844 22624
rect 15197 22593 15209 22596
rect 15151 22587 15209 22593
rect 15838 22584 15844 22596
rect 15896 22584 15902 22636
rect 17494 22584 17500 22636
rect 17552 22624 17558 22636
rect 18874 22624 18880 22636
rect 17552 22596 18880 22624
rect 17552 22584 17558 22596
rect 18874 22584 18880 22596
rect 18932 22584 18938 22636
rect 18984 22633 19012 22664
rect 19334 22652 19340 22664
rect 19392 22652 19398 22704
rect 23290 22652 23296 22704
rect 23348 22692 23354 22704
rect 24314 22695 24372 22701
rect 24314 22692 24326 22695
rect 23348 22664 24326 22692
rect 23348 22652 23354 22664
rect 24314 22661 24326 22664
rect 24360 22661 24372 22695
rect 24314 22655 24372 22661
rect 25222 22652 25228 22704
rect 25280 22692 25286 22704
rect 25317 22695 25375 22701
rect 25317 22692 25329 22695
rect 25280 22664 25329 22692
rect 25280 22652 25286 22664
rect 25317 22661 25329 22664
rect 25363 22661 25375 22695
rect 26160 22692 26188 22723
rect 28074 22720 28080 22732
rect 28132 22720 28138 22772
rect 30837 22763 30895 22769
rect 30837 22729 30849 22763
rect 30883 22760 30895 22763
rect 31110 22760 31116 22772
rect 30883 22732 31116 22760
rect 30883 22729 30895 22732
rect 30837 22723 30895 22729
rect 31110 22720 31116 22732
rect 31168 22720 31174 22772
rect 28902 22692 28908 22704
rect 26160 22664 27568 22692
rect 25317 22655 25375 22661
rect 18969 22627 19027 22633
rect 18969 22593 18981 22627
rect 19015 22593 19027 22627
rect 18969 22587 19027 22593
rect 19058 22584 19064 22636
rect 19116 22624 19122 22636
rect 19245 22627 19303 22633
rect 19116 22596 19161 22624
rect 19116 22584 19122 22596
rect 19245 22593 19257 22627
rect 19291 22593 19303 22627
rect 19245 22587 19303 22593
rect 18049 22559 18107 22565
rect 14752 22528 16712 22556
rect 7524 22460 8248 22488
rect 7524 22448 7530 22460
rect 4706 22420 4712 22432
rect 4667 22392 4712 22420
rect 4706 22380 4712 22392
rect 4764 22380 4770 22432
rect 6825 22423 6883 22429
rect 6825 22389 6837 22423
rect 6871 22420 6883 22423
rect 6914 22420 6920 22432
rect 6871 22392 6920 22420
rect 6871 22389 6883 22392
rect 6825 22383 6883 22389
rect 6914 22380 6920 22392
rect 6972 22380 6978 22432
rect 15286 22420 15292 22432
rect 15247 22392 15292 22420
rect 15286 22380 15292 22392
rect 15344 22380 15350 22432
rect 15930 22420 15936 22432
rect 15891 22392 15936 22420
rect 15930 22380 15936 22392
rect 15988 22420 15994 22432
rect 16390 22420 16396 22432
rect 15988 22392 16396 22420
rect 15988 22380 15994 22392
rect 16390 22380 16396 22392
rect 16448 22380 16454 22432
rect 16684 22429 16712 22528
rect 18049 22525 18061 22559
rect 18095 22556 18107 22559
rect 18095 22528 19196 22556
rect 18095 22525 18107 22528
rect 18049 22519 18107 22525
rect 16669 22423 16727 22429
rect 16669 22389 16681 22423
rect 16715 22420 16727 22423
rect 18506 22420 18512 22432
rect 16715 22392 18512 22420
rect 16715 22389 16727 22392
rect 16669 22383 16727 22389
rect 18506 22380 18512 22392
rect 18564 22380 18570 22432
rect 19168 22420 19196 22528
rect 19260 22488 19288 22587
rect 19426 22584 19432 22636
rect 19484 22624 19490 22636
rect 20717 22627 20775 22633
rect 20717 22624 20729 22627
rect 19484 22596 20729 22624
rect 19484 22584 19490 22596
rect 20717 22593 20729 22596
rect 20763 22593 20775 22627
rect 25501 22627 25559 22633
rect 25501 22624 25513 22627
rect 20717 22587 20775 22593
rect 21836 22596 25513 22624
rect 20993 22559 21051 22565
rect 20993 22525 21005 22559
rect 21039 22556 21051 22559
rect 21634 22556 21640 22568
rect 21039 22528 21640 22556
rect 21039 22525 21051 22528
rect 20993 22519 21051 22525
rect 21634 22516 21640 22528
rect 21692 22556 21698 22568
rect 21836 22565 21864 22596
rect 25501 22593 25513 22596
rect 25547 22624 25559 22627
rect 26234 22624 26240 22636
rect 25547 22596 26240 22624
rect 25547 22593 25559 22596
rect 25501 22587 25559 22593
rect 26234 22584 26240 22596
rect 26292 22584 26298 22636
rect 27430 22624 27436 22636
rect 27080 22596 27436 22624
rect 21821 22559 21879 22565
rect 21821 22556 21833 22559
rect 21692 22528 21833 22556
rect 21692 22516 21698 22528
rect 21821 22525 21833 22528
rect 21867 22525 21879 22559
rect 21821 22519 21879 22525
rect 22097 22559 22155 22565
rect 22097 22525 22109 22559
rect 22143 22525 22155 22559
rect 22097 22519 22155 22525
rect 19978 22488 19984 22500
rect 19260 22460 19984 22488
rect 19978 22448 19984 22460
rect 20036 22488 20042 22500
rect 22112 22488 22140 22519
rect 24578 22516 24584 22568
rect 24636 22556 24642 22568
rect 26786 22556 26792 22568
rect 24636 22528 26792 22556
rect 24636 22516 24642 22528
rect 26786 22516 26792 22528
rect 26844 22556 26850 22568
rect 26970 22556 26976 22568
rect 26844 22528 26976 22556
rect 26844 22516 26850 22528
rect 26970 22516 26976 22528
rect 27028 22516 27034 22568
rect 20036 22460 22140 22488
rect 20036 22448 20042 22460
rect 25222 22448 25228 22500
rect 25280 22488 25286 22500
rect 27080 22488 27108 22596
rect 27430 22584 27436 22596
rect 27488 22584 27494 22636
rect 25280 22460 27108 22488
rect 27540 22488 27568 22664
rect 27724 22664 28908 22692
rect 27724 22633 27752 22664
rect 28902 22652 28908 22664
rect 28960 22652 28966 22704
rect 28994 22652 29000 22704
rect 29052 22692 29058 22704
rect 29181 22695 29239 22701
rect 29181 22692 29193 22695
rect 29052 22664 29193 22692
rect 29052 22652 29058 22664
rect 29181 22661 29193 22664
rect 29227 22692 29239 22695
rect 29546 22692 29552 22704
rect 29227 22664 29552 22692
rect 29227 22661 29239 22664
rect 29181 22655 29239 22661
rect 29546 22652 29552 22664
rect 29604 22652 29610 22704
rect 27617 22627 27675 22633
rect 27617 22593 27629 22627
rect 27663 22593 27675 22627
rect 27617 22587 27675 22593
rect 27709 22627 27767 22633
rect 27709 22593 27721 22627
rect 27755 22593 27767 22627
rect 27709 22587 27767 22593
rect 27632 22556 27660 22587
rect 27798 22584 27804 22636
rect 27856 22624 27862 22636
rect 27856 22596 27901 22624
rect 27856 22584 27862 22596
rect 29086 22584 29092 22636
rect 29144 22624 29150 22636
rect 29365 22627 29423 22633
rect 29365 22624 29377 22627
rect 29144 22596 29377 22624
rect 29144 22584 29150 22596
rect 29365 22593 29377 22596
rect 29411 22624 29423 22627
rect 29914 22624 29920 22636
rect 29411 22596 29920 22624
rect 29411 22593 29423 22596
rect 29365 22587 29423 22593
rect 29914 22584 29920 22596
rect 29972 22584 29978 22636
rect 30190 22624 30196 22636
rect 30151 22596 30196 22624
rect 30190 22584 30196 22596
rect 30248 22584 30254 22636
rect 30374 22624 30380 22636
rect 30335 22596 30380 22624
rect 30374 22584 30380 22596
rect 30432 22584 30438 22636
rect 30466 22584 30472 22636
rect 30524 22624 30530 22636
rect 30650 22633 30656 22636
rect 30607 22627 30656 22633
rect 30524 22596 30569 22624
rect 30524 22584 30530 22596
rect 30607 22593 30619 22627
rect 30653 22593 30656 22627
rect 30607 22587 30656 22593
rect 30650 22584 30656 22587
rect 30708 22584 30714 22636
rect 31478 22624 31484 22636
rect 31391 22596 31484 22624
rect 31478 22584 31484 22596
rect 31536 22624 31542 22636
rect 32125 22627 32183 22633
rect 32125 22624 32137 22627
rect 31536 22596 32137 22624
rect 31536 22584 31542 22596
rect 32125 22593 32137 22596
rect 32171 22593 32183 22627
rect 32125 22587 32183 22593
rect 28997 22559 29055 22565
rect 28997 22556 29009 22559
rect 27632 22528 29009 22556
rect 28997 22525 29009 22528
rect 29043 22525 29055 22559
rect 28997 22519 29055 22525
rect 29454 22488 29460 22500
rect 27540 22460 29460 22488
rect 25280 22448 25286 22460
rect 29454 22448 29460 22460
rect 29512 22448 29518 22500
rect 31110 22448 31116 22500
rect 31168 22488 31174 22500
rect 31297 22491 31355 22497
rect 31297 22488 31309 22491
rect 31168 22460 31309 22488
rect 31168 22448 31174 22460
rect 31297 22457 31309 22460
rect 31343 22457 31355 22491
rect 67634 22488 67640 22500
rect 67595 22460 67640 22488
rect 31297 22451 31355 22457
rect 67634 22448 67640 22460
rect 67692 22448 67698 22500
rect 20070 22420 20076 22432
rect 19168 22392 20076 22420
rect 20070 22380 20076 22392
rect 20128 22380 20134 22432
rect 22922 22380 22928 22432
rect 22980 22420 22986 22432
rect 23201 22423 23259 22429
rect 23201 22420 23213 22423
rect 22980 22392 23213 22420
rect 22980 22380 22986 22392
rect 23201 22389 23213 22392
rect 23247 22389 23259 22423
rect 23201 22383 23259 22389
rect 28994 22380 29000 22432
rect 29052 22420 29058 22432
rect 29178 22420 29184 22432
rect 29052 22392 29184 22420
rect 29052 22380 29058 22392
rect 29178 22380 29184 22392
rect 29236 22380 29242 22432
rect 1104 22330 68816 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 65654 22330
rect 65706 22278 65718 22330
rect 65770 22278 65782 22330
rect 65834 22278 65846 22330
rect 65898 22278 65910 22330
rect 65962 22278 68816 22330
rect 1104 22256 68816 22278
rect 1946 22176 1952 22228
rect 2004 22216 2010 22228
rect 2041 22219 2099 22225
rect 2041 22216 2053 22219
rect 2004 22188 2053 22216
rect 2004 22176 2010 22188
rect 2041 22185 2053 22188
rect 2087 22185 2099 22219
rect 2041 22179 2099 22185
rect 5077 22219 5135 22225
rect 5077 22185 5089 22219
rect 5123 22216 5135 22219
rect 5166 22216 5172 22228
rect 5123 22188 5172 22216
rect 5123 22185 5135 22188
rect 5077 22179 5135 22185
rect 5166 22176 5172 22188
rect 5224 22176 5230 22228
rect 7282 22176 7288 22228
rect 7340 22216 7346 22228
rect 15930 22216 15936 22228
rect 7340 22188 15936 22216
rect 7340 22176 7346 22188
rect 15930 22176 15936 22188
rect 15988 22176 15994 22228
rect 18693 22219 18751 22225
rect 18693 22185 18705 22219
rect 18739 22216 18751 22219
rect 19058 22216 19064 22228
rect 18739 22188 19064 22216
rect 18739 22185 18751 22188
rect 18693 22179 18751 22185
rect 19058 22176 19064 22188
rect 19116 22176 19122 22228
rect 22741 22219 22799 22225
rect 22741 22185 22753 22219
rect 22787 22216 22799 22219
rect 22830 22216 22836 22228
rect 22787 22188 22836 22216
rect 22787 22185 22799 22188
rect 22741 22179 22799 22185
rect 22830 22176 22836 22188
rect 22888 22176 22894 22228
rect 23106 22176 23112 22228
rect 23164 22216 23170 22228
rect 23293 22219 23351 22225
rect 23293 22216 23305 22219
rect 23164 22188 23305 22216
rect 23164 22176 23170 22188
rect 23293 22185 23305 22188
rect 23339 22185 23351 22219
rect 23293 22179 23351 22185
rect 23750 22176 23756 22228
rect 23808 22216 23814 22228
rect 27617 22219 27675 22225
rect 27617 22216 27629 22219
rect 23808 22188 27629 22216
rect 23808 22176 23814 22188
rect 27617 22185 27629 22188
rect 27663 22216 27675 22219
rect 27798 22216 27804 22228
rect 27663 22188 27804 22216
rect 27663 22185 27675 22188
rect 27617 22179 27675 22185
rect 27798 22176 27804 22188
rect 27856 22176 27862 22228
rect 30374 22216 30380 22228
rect 30335 22188 30380 22216
rect 30374 22176 30380 22188
rect 30432 22176 30438 22228
rect 14274 22108 14280 22160
rect 14332 22148 14338 22160
rect 14332 22120 15332 22148
rect 14332 22108 14338 22120
rect 3050 22080 3056 22092
rect 3011 22052 3056 22080
rect 3050 22040 3056 22052
rect 3108 22040 3114 22092
rect 5258 22040 5264 22092
rect 5316 22080 5322 22092
rect 5316 22052 5488 22080
rect 5316 22040 5322 22052
rect 1670 22012 1676 22024
rect 1631 21984 1676 22012
rect 1670 21972 1676 21984
rect 1728 21972 1734 22024
rect 1857 22015 1915 22021
rect 1857 21981 1869 22015
rect 1903 22012 1915 22015
rect 4614 22012 4620 22024
rect 1903 21984 4620 22012
rect 1903 21981 1915 21984
rect 1857 21975 1915 21981
rect 4614 21972 4620 21984
rect 4672 21972 4678 22024
rect 5460 22021 5488 22052
rect 6270 22040 6276 22092
rect 6328 22080 6334 22092
rect 7098 22080 7104 22092
rect 6328 22052 7104 22080
rect 6328 22040 6334 22052
rect 7098 22040 7104 22052
rect 7156 22080 7162 22092
rect 7285 22083 7343 22089
rect 7285 22080 7297 22083
rect 7156 22052 7297 22080
rect 7156 22040 7162 22052
rect 7285 22049 7297 22052
rect 7331 22049 7343 22083
rect 7285 22043 7343 22049
rect 8110 22040 8116 22092
rect 8168 22080 8174 22092
rect 8168 22052 11100 22080
rect 8168 22040 8174 22052
rect 5445 22015 5503 22021
rect 5445 21981 5457 22015
rect 5491 21981 5503 22015
rect 5445 21975 5503 21981
rect 7009 22015 7067 22021
rect 7009 21981 7021 22015
rect 7055 22012 7067 22015
rect 8846 22012 8852 22024
rect 7055 21984 8852 22012
rect 7055 21981 7067 21984
rect 7009 21975 7067 21981
rect 8846 21972 8852 21984
rect 8904 21972 8910 22024
rect 5261 21947 5319 21953
rect 5261 21913 5273 21947
rect 5307 21944 5319 21947
rect 5810 21944 5816 21956
rect 5307 21916 5816 21944
rect 5307 21913 5319 21916
rect 5261 21907 5319 21913
rect 5810 21904 5816 21916
rect 5868 21904 5874 21956
rect 9030 21904 9036 21956
rect 9088 21944 9094 21956
rect 9125 21947 9183 21953
rect 9125 21944 9137 21947
rect 9088 21916 9137 21944
rect 9088 21904 9094 21916
rect 9125 21913 9137 21916
rect 9171 21913 9183 21947
rect 9306 21944 9312 21956
rect 9267 21916 9312 21944
rect 9125 21907 9183 21913
rect 9306 21904 9312 21916
rect 9364 21944 9370 21956
rect 9861 21947 9919 21953
rect 9861 21944 9873 21947
rect 9364 21916 9873 21944
rect 9364 21904 9370 21916
rect 9861 21913 9873 21916
rect 9907 21913 9919 21947
rect 9861 21907 9919 21913
rect 10045 21947 10103 21953
rect 10045 21913 10057 21947
rect 10091 21944 10103 21947
rect 10962 21944 10968 21956
rect 10091 21916 10968 21944
rect 10091 21913 10103 21916
rect 10045 21907 10103 21913
rect 10962 21904 10968 21916
rect 11020 21904 11026 21956
rect 11072 21944 11100 22052
rect 11146 22040 11152 22092
rect 11204 22080 11210 22092
rect 11204 22052 15240 22080
rect 11204 22040 11210 22052
rect 14826 21972 14832 22024
rect 14884 22012 14890 22024
rect 15212 22021 15240 22052
rect 15304 22021 15332 22120
rect 15838 22108 15844 22160
rect 15896 22148 15902 22160
rect 28534 22148 28540 22160
rect 15896 22120 16804 22148
rect 15896 22108 15902 22120
rect 15396 22052 16712 22080
rect 14921 22015 14979 22021
rect 14921 22012 14933 22015
rect 14884 21984 14933 22012
rect 14884 21972 14890 21984
rect 14921 21981 14933 21984
rect 14967 21981 14979 22015
rect 14921 21975 14979 21981
rect 15197 22015 15255 22021
rect 15197 21981 15209 22015
rect 15243 21981 15255 22015
rect 15197 21975 15255 21981
rect 15289 22015 15347 22021
rect 15289 21981 15301 22015
rect 15335 21981 15347 22015
rect 15289 21975 15347 21981
rect 11072 21916 14596 21944
rect 2498 21876 2504 21888
rect 2459 21848 2504 21876
rect 2498 21836 2504 21848
rect 2556 21836 2562 21888
rect 3878 21836 3884 21888
rect 3936 21876 3942 21888
rect 3973 21879 4031 21885
rect 3973 21876 3985 21879
rect 3936 21848 3985 21876
rect 3936 21836 3942 21848
rect 3973 21845 3985 21848
rect 4019 21845 4031 21879
rect 3973 21839 4031 21845
rect 5997 21879 6055 21885
rect 5997 21845 6009 21879
rect 6043 21876 6055 21879
rect 6086 21876 6092 21888
rect 6043 21848 6092 21876
rect 6043 21845 6055 21848
rect 5997 21839 6055 21845
rect 6086 21836 6092 21848
rect 6144 21836 6150 21888
rect 6546 21836 6552 21888
rect 6604 21876 6610 21888
rect 6822 21876 6828 21888
rect 6604 21848 6828 21876
rect 6604 21836 6610 21848
rect 6822 21836 6828 21848
rect 6880 21876 6886 21888
rect 7745 21879 7803 21885
rect 7745 21876 7757 21879
rect 6880 21848 7757 21876
rect 6880 21836 6886 21848
rect 7745 21845 7757 21848
rect 7791 21845 7803 21879
rect 7745 21839 7803 21845
rect 8294 21836 8300 21888
rect 8352 21876 8358 21888
rect 8941 21879 8999 21885
rect 8941 21876 8953 21879
rect 8352 21848 8953 21876
rect 8352 21836 8358 21848
rect 8941 21845 8953 21848
rect 8987 21845 8999 21879
rect 8941 21839 8999 21845
rect 10134 21836 10140 21888
rect 10192 21876 10198 21888
rect 10229 21879 10287 21885
rect 10229 21876 10241 21879
rect 10192 21848 10241 21876
rect 10192 21836 10198 21848
rect 10229 21845 10241 21848
rect 10275 21845 10287 21879
rect 10229 21839 10287 21845
rect 12802 21836 12808 21888
rect 12860 21876 12866 21888
rect 14366 21876 14372 21888
rect 12860 21848 14372 21876
rect 12860 21836 12866 21848
rect 14366 21836 14372 21848
rect 14424 21836 14430 21888
rect 14568 21876 14596 21916
rect 14734 21904 14740 21956
rect 14792 21944 14798 21956
rect 15102 21944 15108 21956
rect 14792 21916 15108 21944
rect 14792 21904 14798 21916
rect 15102 21904 15108 21916
rect 15160 21904 15166 21956
rect 15396 21876 15424 22052
rect 16684 22021 16712 22052
rect 16776 22021 16804 22120
rect 19306 22120 22692 22148
rect 18046 22040 18052 22092
rect 18104 22080 18110 22092
rect 19306 22080 19334 22120
rect 22664 22092 22692 22120
rect 23308 22120 28540 22148
rect 21634 22080 21640 22092
rect 18104 22052 19334 22080
rect 21595 22052 21640 22080
rect 18104 22040 18110 22052
rect 21634 22040 21640 22052
rect 21692 22040 21698 22092
rect 22646 22040 22652 22092
rect 22704 22080 22710 22092
rect 23308 22080 23336 22120
rect 28534 22108 28540 22120
rect 28592 22108 28598 22160
rect 26234 22080 26240 22092
rect 22704 22052 23336 22080
rect 26195 22052 26240 22080
rect 22704 22040 22710 22052
rect 16301 22015 16359 22021
rect 16301 21981 16313 22015
rect 16347 21981 16359 22015
rect 16301 21975 16359 21981
rect 16449 22015 16507 22021
rect 16449 21981 16461 22015
rect 16495 22012 16507 22015
rect 16669 22015 16727 22021
rect 16495 21981 16528 22012
rect 16449 21975 16528 21981
rect 16669 21981 16681 22015
rect 16715 21981 16727 22015
rect 16669 21975 16727 21981
rect 16766 22015 16824 22021
rect 16766 21981 16778 22015
rect 16812 22012 16824 22015
rect 17405 22015 17463 22021
rect 17405 22012 17417 22015
rect 16812 21984 17417 22012
rect 16812 21981 16824 21984
rect 16766 21975 16824 21981
rect 17405 21981 17417 21984
rect 17451 22012 17463 22015
rect 17586 22012 17592 22024
rect 17451 21984 17592 22012
rect 17451 21981 17463 21984
rect 17405 21975 17463 21981
rect 14568 21848 15424 21876
rect 15473 21879 15531 21885
rect 15473 21845 15485 21879
rect 15519 21876 15531 21879
rect 16316 21876 16344 21975
rect 15519 21848 16344 21876
rect 16500 21876 16528 21975
rect 17586 21972 17592 21984
rect 17644 21972 17650 22024
rect 18322 22012 18328 22024
rect 18283 21984 18328 22012
rect 18322 21972 18328 21984
rect 18380 21972 18386 22024
rect 18506 22012 18512 22024
rect 18467 21984 18512 22012
rect 18506 21972 18512 21984
rect 18564 21972 18570 22024
rect 20254 21972 20260 22024
rect 20312 22012 20318 22024
rect 20625 22015 20683 22021
rect 20625 22012 20637 22015
rect 20312 21984 20637 22012
rect 20312 21972 20318 21984
rect 20625 21981 20637 21984
rect 20671 22012 20683 22015
rect 21910 22012 21916 22024
rect 20671 21984 21916 22012
rect 20671 21981 20683 21984
rect 20625 21975 20683 21981
rect 21910 21972 21916 21984
rect 21968 21972 21974 22024
rect 22370 22012 22376 22024
rect 22331 21984 22376 22012
rect 22370 21972 22376 21984
rect 22428 21972 22434 22024
rect 23201 22015 23259 22021
rect 23201 21981 23213 22015
rect 23247 22012 23259 22015
rect 23308 22012 23336 22052
rect 26234 22040 26240 22052
rect 26292 22040 26298 22092
rect 30926 22080 30932 22092
rect 30887 22052 30932 22080
rect 30926 22040 30932 22052
rect 30984 22040 30990 22092
rect 23247 21984 23336 22012
rect 23385 22015 23443 22021
rect 23247 21981 23259 21984
rect 23201 21975 23259 21981
rect 23385 21981 23397 22015
rect 23431 22012 23443 22015
rect 23566 22012 23572 22024
rect 23431 21984 23572 22012
rect 23431 21981 23443 21984
rect 23385 21975 23443 21981
rect 23566 21972 23572 21984
rect 23624 21972 23630 22024
rect 25866 22012 25872 22024
rect 25536 21984 25872 22012
rect 16574 21904 16580 21956
rect 16632 21944 16638 21956
rect 17954 21944 17960 21956
rect 16632 21916 16677 21944
rect 16868 21916 17960 21944
rect 16632 21904 16638 21916
rect 16868 21876 16896 21916
rect 17954 21904 17960 21916
rect 18012 21904 18018 21956
rect 22557 21947 22615 21953
rect 22557 21913 22569 21947
rect 22603 21944 22615 21947
rect 22830 21944 22836 21956
rect 22603 21916 22836 21944
rect 22603 21913 22615 21916
rect 22557 21907 22615 21913
rect 22830 21904 22836 21916
rect 22888 21904 22894 21956
rect 25536 21944 25564 21984
rect 25866 21972 25872 21984
rect 25924 21972 25930 22024
rect 26510 22012 26516 22024
rect 26471 21984 26516 22012
rect 26510 21972 26516 21984
rect 26568 21972 26574 22024
rect 30009 22015 30067 22021
rect 30009 21981 30021 22015
rect 30055 22012 30067 22015
rect 31018 22012 31024 22024
rect 30055 21984 31024 22012
rect 30055 21981 30067 21984
rect 30009 21975 30067 21981
rect 31018 21972 31024 21984
rect 31076 21972 31082 22024
rect 32950 22012 32956 22024
rect 31128 21984 32956 22012
rect 24826 21916 25564 21944
rect 25593 21947 25651 21953
rect 16500 21848 16896 21876
rect 16945 21879 17003 21885
rect 15519 21845 15531 21848
rect 15473 21839 15531 21845
rect 16945 21845 16957 21879
rect 16991 21876 17003 21879
rect 17218 21876 17224 21888
rect 16991 21848 17224 21876
rect 16991 21845 17003 21848
rect 16945 21839 17003 21845
rect 17218 21836 17224 21848
rect 17276 21836 17282 21888
rect 18874 21836 18880 21888
rect 18932 21876 18938 21888
rect 19337 21879 19395 21885
rect 19337 21876 19349 21879
rect 18932 21848 19349 21876
rect 18932 21836 18938 21848
rect 19337 21845 19349 21848
rect 19383 21876 19395 21879
rect 24826 21876 24854 21916
rect 25593 21913 25605 21947
rect 25639 21913 25651 21947
rect 25593 21907 25651 21913
rect 25777 21947 25835 21953
rect 25777 21913 25789 21947
rect 25823 21944 25835 21947
rect 27338 21944 27344 21956
rect 25823 21916 27344 21944
rect 25823 21913 25835 21916
rect 25777 21907 25835 21913
rect 19383 21848 24854 21876
rect 25041 21879 25099 21885
rect 19383 21845 19395 21848
rect 19337 21839 19395 21845
rect 25041 21845 25053 21879
rect 25087 21876 25099 21879
rect 25314 21876 25320 21888
rect 25087 21848 25320 21876
rect 25087 21845 25099 21848
rect 25041 21839 25099 21845
rect 25314 21836 25320 21848
rect 25372 21876 25378 21888
rect 25608 21876 25636 21907
rect 27338 21904 27344 21916
rect 27396 21904 27402 21956
rect 29822 21904 29828 21956
rect 29880 21944 29886 21956
rect 30193 21947 30251 21953
rect 30193 21944 30205 21947
rect 29880 21916 30205 21944
rect 29880 21904 29886 21916
rect 30193 21913 30205 21916
rect 30239 21944 30251 21947
rect 31128 21944 31156 21984
rect 32950 21972 32956 21984
rect 33008 21972 33014 22024
rect 34146 22012 34152 22024
rect 34107 21984 34152 22012
rect 34146 21972 34152 21984
rect 34204 21972 34210 22024
rect 31202 21953 31208 21956
rect 30239 21916 31156 21944
rect 30239 21913 30251 21916
rect 30193 21907 30251 21913
rect 31196 21907 31208 21953
rect 31260 21944 31266 21956
rect 31260 21916 31296 21944
rect 31202 21904 31208 21907
rect 31260 21904 31266 21916
rect 33594 21904 33600 21956
rect 33652 21944 33658 21956
rect 33882 21947 33940 21953
rect 33882 21944 33894 21947
rect 33652 21916 33894 21944
rect 33652 21904 33658 21916
rect 33882 21913 33894 21916
rect 33928 21913 33940 21947
rect 36357 21947 36415 21953
rect 36357 21944 36369 21947
rect 33882 21907 33940 21913
rect 35912 21916 36369 21944
rect 35912 21888 35940 21916
rect 36357 21913 36369 21916
rect 36403 21913 36415 21947
rect 36357 21907 36415 21913
rect 25372 21848 25636 21876
rect 25372 21836 25378 21848
rect 28074 21836 28080 21888
rect 28132 21876 28138 21888
rect 32122 21876 32128 21888
rect 28132 21848 32128 21876
rect 28132 21836 28138 21848
rect 32122 21836 32128 21848
rect 32180 21836 32186 21888
rect 32306 21876 32312 21888
rect 32267 21848 32312 21876
rect 32306 21836 32312 21848
rect 32364 21836 32370 21888
rect 32766 21876 32772 21888
rect 32727 21848 32772 21876
rect 32766 21836 32772 21848
rect 32824 21836 32830 21888
rect 35894 21876 35900 21888
rect 35855 21848 35900 21876
rect 35894 21836 35900 21848
rect 35952 21836 35958 21888
rect 37642 21876 37648 21888
rect 37603 21848 37648 21876
rect 37642 21836 37648 21848
rect 37700 21836 37706 21888
rect 1104 21786 68816 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 68816 21786
rect 1104 21712 68816 21734
rect 2961 21675 3019 21681
rect 2961 21641 2973 21675
rect 3007 21672 3019 21675
rect 3142 21672 3148 21684
rect 3007 21644 3148 21672
rect 3007 21641 3019 21644
rect 2961 21635 3019 21641
rect 3142 21632 3148 21644
rect 3200 21632 3206 21684
rect 3970 21632 3976 21684
rect 4028 21672 4034 21684
rect 6365 21675 6423 21681
rect 6365 21672 6377 21675
rect 4028 21644 6377 21672
rect 4028 21632 4034 21644
rect 6365 21641 6377 21644
rect 6411 21641 6423 21675
rect 6365 21635 6423 21641
rect 7101 21675 7159 21681
rect 7101 21641 7113 21675
rect 7147 21672 7159 21675
rect 7282 21672 7288 21684
rect 7147 21644 7288 21672
rect 7147 21641 7159 21644
rect 7101 21635 7159 21641
rect 7282 21632 7288 21644
rect 7340 21632 7346 21684
rect 8018 21632 8024 21684
rect 8076 21672 8082 21684
rect 9306 21672 9312 21684
rect 8076 21644 9312 21672
rect 8076 21632 8082 21644
rect 9306 21632 9312 21644
rect 9364 21672 9370 21684
rect 13817 21675 13875 21681
rect 9364 21644 11652 21672
rect 9364 21632 9370 21644
rect 11624 21616 11652 21644
rect 13817 21641 13829 21675
rect 13863 21641 13875 21675
rect 13817 21635 13875 21641
rect 2866 21564 2872 21616
rect 2924 21604 2930 21616
rect 4706 21613 4712 21616
rect 4700 21604 4712 21613
rect 2924 21576 4108 21604
rect 4667 21576 4712 21604
rect 2924 21564 2930 21576
rect 4080 21548 4108 21576
rect 4700 21567 4712 21576
rect 4706 21564 4712 21567
rect 4764 21564 4770 21616
rect 11146 21604 11152 21616
rect 8680 21576 11152 21604
rect 3145 21539 3203 21545
rect 3145 21505 3157 21539
rect 3191 21536 3203 21539
rect 3326 21536 3332 21548
rect 3191 21508 3332 21536
rect 3191 21505 3203 21508
rect 3145 21499 3203 21505
rect 3326 21496 3332 21508
rect 3384 21496 3390 21548
rect 3697 21539 3755 21545
rect 3697 21505 3709 21539
rect 3743 21536 3755 21539
rect 3878 21536 3884 21548
rect 3743 21508 3884 21536
rect 3743 21505 3755 21508
rect 3697 21499 3755 21505
rect 3878 21496 3884 21508
rect 3936 21496 3942 21548
rect 4062 21496 4068 21548
rect 4120 21536 4126 21548
rect 4433 21539 4491 21545
rect 4433 21536 4445 21539
rect 4120 21508 4445 21536
rect 4120 21496 4126 21508
rect 4433 21505 4445 21508
rect 4479 21505 4491 21539
rect 6362 21536 6368 21548
rect 6323 21508 6368 21536
rect 4433 21499 4491 21505
rect 6362 21496 6368 21508
rect 6420 21496 6426 21548
rect 6546 21536 6552 21548
rect 6507 21508 6552 21536
rect 6546 21496 6552 21508
rect 6604 21496 6610 21548
rect 7742 21496 7748 21548
rect 7800 21536 7806 21548
rect 7909 21539 7967 21545
rect 7909 21536 7921 21539
rect 7800 21508 7921 21536
rect 7800 21496 7806 21508
rect 7909 21505 7921 21508
rect 7955 21505 7967 21539
rect 7909 21499 7967 21505
rect 6638 21428 6644 21480
rect 6696 21468 6702 21480
rect 7653 21471 7711 21477
rect 7653 21468 7665 21471
rect 6696 21440 7665 21468
rect 6696 21428 6702 21440
rect 7653 21437 7665 21440
rect 7699 21437 7711 21471
rect 7653 21431 7711 21437
rect 5810 21400 5816 21412
rect 5723 21372 5816 21400
rect 5810 21360 5816 21372
rect 5868 21360 5874 21412
rect 1854 21292 1860 21344
rect 1912 21332 1918 21344
rect 2041 21335 2099 21341
rect 2041 21332 2053 21335
rect 1912 21304 2053 21332
rect 1912 21292 1918 21304
rect 2041 21301 2053 21304
rect 2087 21332 2099 21335
rect 2590 21332 2596 21344
rect 2087 21304 2596 21332
rect 2087 21301 2099 21304
rect 2041 21295 2099 21301
rect 2590 21292 2596 21304
rect 2648 21292 2654 21344
rect 3234 21292 3240 21344
rect 3292 21332 3298 21344
rect 3789 21335 3847 21341
rect 3789 21332 3801 21335
rect 3292 21304 3801 21332
rect 3292 21292 3298 21304
rect 3789 21301 3801 21304
rect 3835 21332 3847 21335
rect 5718 21332 5724 21344
rect 3835 21304 5724 21332
rect 3835 21301 3847 21304
rect 3789 21295 3847 21301
rect 5718 21292 5724 21304
rect 5776 21292 5782 21344
rect 5828 21332 5856 21360
rect 8680 21332 8708 21576
rect 11146 21564 11152 21576
rect 11204 21564 11210 21616
rect 11606 21604 11612 21616
rect 11519 21576 11612 21604
rect 11606 21564 11612 21576
rect 11664 21564 11670 21616
rect 11793 21607 11851 21613
rect 11793 21573 11805 21607
rect 11839 21604 11851 21607
rect 13832 21604 13860 21635
rect 15010 21632 15016 21684
rect 15068 21672 15074 21684
rect 16574 21672 16580 21684
rect 15068 21644 16580 21672
rect 15068 21632 15074 21644
rect 16574 21632 16580 21644
rect 16632 21632 16638 21684
rect 16761 21675 16819 21681
rect 16761 21641 16773 21675
rect 16807 21672 16819 21675
rect 17678 21672 17684 21684
rect 16807 21644 17684 21672
rect 16807 21641 16819 21644
rect 16761 21635 16819 21641
rect 17678 21632 17684 21644
rect 17736 21632 17742 21684
rect 17957 21675 18015 21681
rect 17957 21641 17969 21675
rect 18003 21672 18015 21675
rect 18046 21672 18052 21684
rect 18003 21644 18052 21672
rect 18003 21641 18015 21644
rect 17957 21635 18015 21641
rect 18046 21632 18052 21644
rect 18104 21632 18110 21684
rect 21269 21675 21327 21681
rect 21269 21641 21281 21675
rect 21315 21672 21327 21675
rect 22370 21672 22376 21684
rect 21315 21644 22376 21672
rect 21315 21641 21327 21644
rect 21269 21635 21327 21641
rect 22370 21632 22376 21644
rect 22428 21632 22434 21684
rect 26694 21672 26700 21684
rect 25332 21644 26700 21672
rect 23569 21607 23627 21613
rect 23569 21604 23581 21607
rect 11839 21576 23581 21604
rect 11839 21573 11851 21576
rect 11793 21567 11851 21573
rect 23569 21573 23581 21576
rect 23615 21573 23627 21607
rect 24305 21607 24363 21613
rect 24305 21604 24317 21607
rect 23569 21567 23627 21573
rect 23676 21576 24317 21604
rect 23676 21548 23704 21576
rect 24305 21573 24317 21576
rect 24351 21573 24363 21607
rect 24305 21567 24363 21573
rect 9674 21496 9680 21548
rect 9732 21536 9738 21548
rect 9841 21539 9899 21545
rect 9841 21536 9853 21539
rect 9732 21508 9853 21536
rect 9732 21496 9738 21508
rect 9841 21505 9853 21508
rect 9887 21505 9899 21539
rect 12434 21536 12440 21548
rect 12395 21508 12440 21536
rect 9841 21499 9899 21505
rect 12434 21496 12440 21508
rect 12492 21496 12498 21548
rect 12710 21545 12716 21548
rect 12704 21499 12716 21545
rect 12768 21536 12774 21548
rect 12768 21508 12804 21536
rect 12710 21496 12716 21499
rect 12768 21496 12774 21508
rect 14366 21496 14372 21548
rect 14424 21536 14430 21548
rect 15565 21539 15623 21545
rect 15565 21536 15577 21539
rect 14424 21508 15577 21536
rect 14424 21496 14430 21508
rect 15565 21505 15577 21508
rect 15611 21536 15623 21539
rect 15838 21536 15844 21548
rect 15611 21508 15844 21536
rect 15611 21505 15623 21508
rect 15565 21499 15623 21505
rect 15838 21496 15844 21508
rect 15896 21496 15902 21548
rect 16942 21536 16948 21548
rect 16903 21508 16948 21536
rect 16942 21496 16948 21508
rect 17000 21496 17006 21548
rect 17586 21496 17592 21548
rect 17644 21536 17650 21548
rect 17865 21539 17923 21545
rect 17865 21536 17877 21539
rect 17644 21508 17877 21536
rect 17644 21496 17650 21508
rect 17865 21505 17877 21508
rect 17911 21505 17923 21539
rect 19794 21536 19800 21548
rect 19852 21545 19858 21548
rect 19764 21508 19800 21536
rect 17865 21499 17923 21505
rect 19794 21496 19800 21508
rect 19852 21499 19864 21545
rect 20070 21536 20076 21548
rect 20031 21508 20076 21536
rect 19852 21496 19858 21499
rect 20070 21496 20076 21508
rect 20128 21496 20134 21548
rect 21082 21536 21088 21548
rect 21043 21508 21088 21536
rect 21082 21496 21088 21508
rect 21140 21496 21146 21548
rect 22649 21539 22707 21545
rect 22649 21505 22661 21539
rect 22695 21536 22707 21539
rect 23106 21536 23112 21548
rect 22695 21508 23112 21536
rect 22695 21505 22707 21508
rect 22649 21499 22707 21505
rect 23106 21496 23112 21508
rect 23164 21496 23170 21548
rect 23293 21539 23351 21545
rect 23293 21505 23305 21539
rect 23339 21505 23351 21539
rect 23293 21499 23351 21505
rect 23477 21539 23535 21545
rect 23477 21505 23489 21539
rect 23523 21505 23535 21539
rect 23658 21536 23664 21548
rect 23619 21508 23664 21536
rect 23477 21499 23535 21505
rect 9214 21428 9220 21480
rect 9272 21468 9278 21480
rect 9585 21471 9643 21477
rect 9585 21468 9597 21471
rect 9272 21440 9597 21468
rect 9272 21428 9278 21440
rect 9585 21437 9597 21440
rect 9631 21437 9643 21471
rect 9585 21431 9643 21437
rect 20714 21428 20720 21480
rect 20772 21468 20778 21480
rect 20901 21471 20959 21477
rect 20901 21468 20913 21471
rect 20772 21440 20913 21468
rect 20772 21428 20778 21440
rect 20901 21437 20913 21440
rect 20947 21437 20959 21471
rect 20901 21431 20959 21437
rect 22373 21471 22431 21477
rect 22373 21437 22385 21471
rect 22419 21437 22431 21471
rect 22373 21431 22431 21437
rect 10962 21400 10968 21412
rect 10923 21372 10968 21400
rect 10962 21360 10968 21372
rect 11020 21360 11026 21412
rect 20070 21360 20076 21412
rect 20128 21400 20134 21412
rect 22388 21400 22416 21431
rect 20128 21372 22416 21400
rect 20128 21360 20134 21372
rect 9030 21332 9036 21344
rect 5828 21304 8708 21332
rect 8991 21304 9036 21332
rect 9030 21292 9036 21304
rect 9088 21292 9094 21344
rect 11790 21292 11796 21344
rect 11848 21332 11854 21344
rect 11977 21335 12035 21341
rect 11977 21332 11989 21335
rect 11848 21304 11989 21332
rect 11848 21292 11854 21304
rect 11977 21301 11989 21304
rect 12023 21301 12035 21335
rect 11977 21295 12035 21301
rect 18693 21335 18751 21341
rect 18693 21301 18705 21335
rect 18739 21332 18751 21335
rect 18874 21332 18880 21344
rect 18739 21304 18880 21332
rect 18739 21301 18751 21304
rect 18693 21295 18751 21301
rect 18874 21292 18880 21304
rect 18932 21292 18938 21344
rect 23308 21332 23336 21499
rect 23492 21468 23520 21499
rect 23658 21496 23664 21508
rect 23716 21496 23722 21548
rect 25332 21545 25360 21644
rect 26694 21632 26700 21644
rect 26752 21632 26758 21684
rect 28629 21675 28687 21681
rect 28629 21641 28641 21675
rect 28675 21672 28687 21675
rect 28902 21672 28908 21684
rect 28675 21644 28908 21672
rect 28675 21641 28687 21644
rect 28629 21635 28687 21641
rect 28902 21632 28908 21644
rect 28960 21632 28966 21684
rect 31113 21675 31171 21681
rect 31113 21641 31125 21675
rect 31159 21672 31171 21675
rect 31202 21672 31208 21684
rect 31159 21644 31208 21672
rect 31159 21641 31171 21644
rect 31113 21635 31171 21641
rect 31202 21632 31208 21644
rect 31260 21632 31266 21684
rect 25501 21607 25559 21613
rect 25501 21573 25513 21607
rect 25547 21604 25559 21607
rect 25547 21576 28856 21604
rect 25547 21573 25559 21576
rect 25501 21567 25559 21573
rect 25133 21539 25191 21545
rect 25133 21536 25145 21539
rect 23860 21508 25145 21536
rect 23566 21468 23572 21480
rect 23492 21440 23572 21468
rect 23566 21428 23572 21440
rect 23624 21428 23630 21480
rect 23860 21409 23888 21508
rect 25133 21505 25145 21508
rect 25179 21505 25191 21539
rect 25133 21499 25191 21505
rect 25281 21539 25360 21545
rect 25281 21505 25293 21539
rect 25327 21508 25360 21539
rect 25327 21505 25339 21508
rect 25281 21499 25339 21505
rect 25406 21496 25412 21548
rect 25464 21536 25470 21548
rect 25598 21539 25656 21545
rect 25464 21508 25509 21536
rect 25464 21496 25470 21508
rect 25598 21505 25610 21539
rect 25644 21505 25656 21539
rect 25598 21499 25656 21505
rect 25498 21428 25504 21480
rect 25556 21468 25562 21480
rect 25613 21468 25641 21499
rect 25866 21496 25872 21548
rect 25924 21536 25930 21548
rect 26421 21539 26479 21545
rect 26421 21536 26433 21539
rect 25924 21508 26433 21536
rect 25924 21496 25930 21508
rect 26421 21505 26433 21508
rect 26467 21536 26479 21539
rect 27249 21539 27307 21545
rect 27249 21536 27261 21539
rect 26467 21508 27261 21536
rect 26467 21505 26479 21508
rect 26421 21499 26479 21505
rect 27249 21505 27261 21508
rect 27295 21505 27307 21539
rect 27249 21499 27307 21505
rect 27341 21539 27399 21545
rect 27341 21505 27353 21539
rect 27387 21505 27399 21539
rect 27341 21499 27399 21505
rect 27433 21539 27491 21545
rect 27433 21505 27445 21539
rect 27479 21505 27491 21539
rect 27433 21499 27491 21505
rect 25556 21440 25641 21468
rect 25556 21428 25562 21440
rect 23845 21403 23903 21409
rect 23845 21369 23857 21403
rect 23891 21369 23903 21403
rect 26418 21400 26424 21412
rect 23845 21363 23903 21369
rect 23952 21372 26424 21400
rect 23952 21332 23980 21372
rect 26418 21360 26424 21372
rect 26476 21360 26482 21412
rect 27356 21400 27384 21499
rect 27448 21468 27476 21499
rect 27522 21496 27528 21548
rect 27580 21536 27586 21548
rect 27617 21539 27675 21545
rect 27617 21536 27629 21539
rect 27580 21508 27629 21536
rect 27580 21496 27586 21508
rect 27617 21505 27629 21508
rect 27663 21505 27675 21539
rect 28534 21536 28540 21548
rect 28495 21508 28540 21536
rect 27617 21499 27675 21505
rect 28534 21496 28540 21508
rect 28592 21496 28598 21548
rect 28718 21536 28724 21548
rect 28679 21508 28724 21536
rect 28718 21496 28724 21508
rect 28776 21496 28782 21548
rect 27706 21468 27712 21480
rect 27448 21440 27712 21468
rect 27706 21428 27712 21440
rect 27764 21428 27770 21480
rect 28828 21468 28856 21576
rect 28920 21536 28948 21632
rect 32766 21604 32772 21616
rect 29288 21576 32772 21604
rect 29181 21539 29239 21545
rect 29181 21536 29193 21539
rect 28920 21508 29193 21536
rect 29181 21505 29193 21508
rect 29227 21505 29239 21539
rect 29181 21499 29239 21505
rect 29288 21468 29316 21576
rect 32766 21564 32772 21576
rect 32824 21604 32830 21616
rect 33137 21607 33195 21613
rect 33137 21604 33149 21607
rect 32824 21576 33149 21604
rect 32824 21564 32830 21576
rect 33137 21573 33149 21576
rect 33183 21573 33195 21607
rect 33137 21567 33195 21573
rect 33962 21564 33968 21616
rect 34020 21604 34026 21616
rect 37642 21604 37648 21616
rect 34020 21576 37648 21604
rect 34020 21564 34026 21576
rect 30190 21496 30196 21548
rect 30248 21536 30254 21548
rect 30469 21539 30527 21545
rect 30469 21536 30481 21539
rect 30248 21508 30481 21536
rect 30248 21496 30254 21508
rect 30469 21505 30481 21508
rect 30515 21505 30527 21539
rect 30650 21536 30656 21548
rect 30611 21508 30656 21536
rect 30469 21499 30527 21505
rect 30650 21496 30656 21508
rect 30708 21496 30714 21548
rect 30745 21539 30803 21545
rect 30745 21505 30757 21539
rect 30791 21505 30803 21539
rect 30745 21499 30803 21505
rect 28828 21440 29316 21468
rect 29457 21471 29515 21477
rect 29457 21437 29469 21471
rect 29503 21468 29515 21471
rect 30760 21468 30788 21499
rect 30834 21496 30840 21548
rect 30892 21536 30898 21548
rect 32953 21539 33011 21545
rect 30892 21508 30937 21536
rect 30892 21496 30898 21508
rect 32953 21505 32965 21539
rect 32999 21536 33011 21539
rect 33410 21536 33416 21548
rect 32999 21508 33416 21536
rect 32999 21505 33011 21508
rect 32953 21499 33011 21505
rect 33410 21496 33416 21508
rect 33468 21536 33474 21548
rect 34517 21539 34575 21545
rect 34517 21536 34529 21539
rect 33468 21508 34529 21536
rect 33468 21496 33474 21508
rect 34517 21505 34529 21508
rect 34563 21505 34575 21539
rect 34517 21499 34575 21505
rect 34701 21539 34759 21545
rect 34701 21505 34713 21539
rect 34747 21505 34759 21539
rect 34701 21499 34759 21505
rect 31386 21468 31392 21480
rect 29503 21440 31392 21468
rect 29503 21437 29515 21440
rect 29457 21431 29515 21437
rect 27430 21400 27436 21412
rect 27343 21372 27436 21400
rect 27430 21360 27436 21372
rect 27488 21400 27494 21412
rect 29472 21400 29500 21431
rect 31386 21428 31392 21440
rect 31444 21428 31450 21480
rect 32122 21428 32128 21480
rect 32180 21468 32186 21480
rect 34716 21468 34744 21499
rect 35618 21496 35624 21548
rect 35676 21536 35682 21548
rect 36740 21545 36768 21576
rect 37642 21564 37648 21576
rect 37700 21564 37706 21616
rect 36458 21539 36516 21545
rect 36458 21536 36470 21539
rect 35676 21508 36470 21536
rect 35676 21496 35682 21508
rect 36458 21505 36470 21508
rect 36504 21505 36516 21539
rect 36458 21499 36516 21505
rect 36725 21539 36783 21545
rect 36725 21505 36737 21539
rect 36771 21505 36783 21539
rect 36725 21499 36783 21505
rect 32180 21440 35388 21468
rect 32180 21428 32186 21440
rect 35360 21409 35388 21440
rect 27488 21372 29500 21400
rect 35345 21403 35403 21409
rect 27488 21360 27494 21372
rect 35345 21369 35357 21403
rect 35391 21369 35403 21403
rect 35345 21363 35403 21369
rect 23308 21304 23980 21332
rect 25777 21335 25835 21341
rect 25777 21301 25789 21335
rect 25823 21332 25835 21335
rect 26050 21332 26056 21344
rect 25823 21304 26056 21332
rect 25823 21301 25835 21304
rect 25777 21295 25835 21301
rect 26050 21292 26056 21304
rect 26108 21292 26114 21344
rect 26973 21335 27031 21341
rect 26973 21301 26985 21335
rect 27019 21332 27031 21335
rect 27062 21332 27068 21344
rect 27019 21304 27068 21332
rect 27019 21301 27031 21304
rect 26973 21295 27031 21301
rect 27062 21292 27068 21304
rect 27120 21292 27126 21344
rect 33134 21292 33140 21344
rect 33192 21332 33198 21344
rect 33321 21335 33379 21341
rect 33321 21332 33333 21335
rect 33192 21304 33333 21332
rect 33192 21292 33198 21304
rect 33321 21301 33333 21304
rect 33367 21301 33379 21335
rect 33321 21295 33379 21301
rect 34790 21292 34796 21344
rect 34848 21332 34854 21344
rect 34885 21335 34943 21341
rect 34885 21332 34897 21335
rect 34848 21304 34897 21332
rect 34848 21292 34854 21304
rect 34885 21301 34897 21304
rect 34931 21301 34943 21335
rect 67634 21332 67640 21344
rect 67595 21304 67640 21332
rect 34885 21295 34943 21301
rect 67634 21292 67640 21304
rect 67692 21292 67698 21344
rect 1104 21242 68816 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 65654 21242
rect 65706 21190 65718 21242
rect 65770 21190 65782 21242
rect 65834 21190 65846 21242
rect 65898 21190 65910 21242
rect 65962 21190 68816 21242
rect 1104 21168 68816 21190
rect 5718 21088 5724 21140
rect 5776 21128 5782 21140
rect 8021 21131 8079 21137
rect 5776 21100 7972 21128
rect 5776 21088 5782 21100
rect 7944 21060 7972 21100
rect 8021 21097 8033 21131
rect 8067 21128 8079 21131
rect 8110 21128 8116 21140
rect 8067 21100 8116 21128
rect 8067 21097 8079 21100
rect 8021 21091 8079 21097
rect 8110 21088 8116 21100
rect 8168 21088 8174 21140
rect 9585 21131 9643 21137
rect 9585 21097 9597 21131
rect 9631 21128 9643 21131
rect 9674 21128 9680 21140
rect 9631 21100 9680 21128
rect 9631 21097 9643 21100
rect 9585 21091 9643 21097
rect 9674 21088 9680 21100
rect 9732 21088 9738 21140
rect 12345 21131 12403 21137
rect 12345 21097 12357 21131
rect 12391 21128 12403 21131
rect 12710 21128 12716 21140
rect 12391 21100 12716 21128
rect 12391 21097 12403 21100
rect 12345 21091 12403 21097
rect 12710 21088 12716 21100
rect 12768 21088 12774 21140
rect 16577 21131 16635 21137
rect 16577 21097 16589 21131
rect 16623 21128 16635 21131
rect 16942 21128 16948 21140
rect 16623 21100 16948 21128
rect 16623 21097 16635 21100
rect 16577 21091 16635 21097
rect 16942 21088 16948 21100
rect 17000 21128 17006 21140
rect 17678 21128 17684 21140
rect 17000 21100 17684 21128
rect 17000 21088 17006 21100
rect 17678 21088 17684 21100
rect 17736 21088 17742 21140
rect 19794 21088 19800 21140
rect 19852 21128 19858 21140
rect 19889 21131 19947 21137
rect 19889 21128 19901 21131
rect 19852 21100 19901 21128
rect 19852 21088 19858 21100
rect 19889 21097 19901 21100
rect 19935 21097 19947 21131
rect 21637 21131 21695 21137
rect 19889 21091 19947 21097
rect 20456 21100 21496 21128
rect 20456 21072 20484 21100
rect 9033 21063 9091 21069
rect 9033 21060 9045 21063
rect 7944 21032 9045 21060
rect 9033 21029 9045 21032
rect 9079 21029 9091 21063
rect 10594 21060 10600 21072
rect 9033 21023 9091 21029
rect 9968 21032 10600 21060
rect 4062 20952 4068 21004
rect 4120 20992 4126 21004
rect 6181 20995 6239 21001
rect 6181 20992 6193 20995
rect 4120 20964 6193 20992
rect 4120 20952 4126 20964
rect 6181 20961 6193 20964
rect 6227 20992 6239 20995
rect 6638 20992 6644 21004
rect 6227 20964 6644 20992
rect 6227 20961 6239 20964
rect 6181 20955 6239 20961
rect 6638 20952 6644 20964
rect 6696 20952 6702 21004
rect 2314 20924 2320 20936
rect 2275 20896 2320 20924
rect 2314 20884 2320 20896
rect 2372 20884 2378 20936
rect 2593 20927 2651 20933
rect 2593 20893 2605 20927
rect 2639 20924 2651 20927
rect 2774 20924 2780 20936
rect 2639 20896 2780 20924
rect 2639 20893 2651 20896
rect 2593 20887 2651 20893
rect 2774 20884 2780 20896
rect 2832 20884 2838 20936
rect 8386 20924 8392 20936
rect 6748 20896 8392 20924
rect 3973 20859 4031 20865
rect 3973 20825 3985 20859
rect 4019 20856 4031 20859
rect 4433 20859 4491 20865
rect 4433 20856 4445 20859
rect 4019 20828 4445 20856
rect 4019 20825 4031 20828
rect 3973 20819 4031 20825
rect 4433 20825 4445 20828
rect 4479 20856 4491 20859
rect 6748 20856 6776 20896
rect 8386 20884 8392 20896
rect 8444 20884 8450 20936
rect 9048 20924 9076 21023
rect 9968 20933 9996 21032
rect 10594 21020 10600 21032
rect 10652 21060 10658 21072
rect 17034 21060 17040 21072
rect 10652 21032 12020 21060
rect 16995 21032 17040 21060
rect 10652 21020 10658 21032
rect 10134 20992 10140 21004
rect 10060 20964 10140 20992
rect 10060 20933 10088 20964
rect 10134 20952 10140 20964
rect 10192 20952 10198 21004
rect 9815 20927 9873 20933
rect 9815 20924 9827 20927
rect 9048 20896 9827 20924
rect 9815 20893 9827 20896
rect 9861 20893 9873 20927
rect 9815 20887 9873 20893
rect 9953 20927 10011 20933
rect 9953 20893 9965 20927
rect 9999 20893 10011 20927
rect 9953 20887 10011 20893
rect 10045 20927 10103 20933
rect 10045 20893 10057 20927
rect 10091 20893 10103 20927
rect 10045 20887 10103 20893
rect 10229 20927 10287 20933
rect 10229 20893 10241 20927
rect 10275 20924 10287 20927
rect 10318 20924 10324 20936
rect 10275 20896 10324 20924
rect 10275 20893 10287 20896
rect 10229 20887 10287 20893
rect 10318 20884 10324 20896
rect 10376 20924 10382 20936
rect 11992 20933 12020 21032
rect 17034 21020 17040 21032
rect 17092 21060 17098 21072
rect 18230 21060 18236 21072
rect 17092 21032 18236 21060
rect 17092 21020 17098 21032
rect 18230 21020 18236 21032
rect 18288 21020 18294 21072
rect 19978 21020 19984 21072
rect 20036 21060 20042 21072
rect 20438 21060 20444 21072
rect 20036 21032 20444 21060
rect 20036 21020 20042 21032
rect 20438 21020 20444 21032
rect 20496 21020 20502 21072
rect 21082 21020 21088 21072
rect 21140 21020 21146 21072
rect 21468 21060 21496 21100
rect 21637 21097 21649 21131
rect 21683 21128 21695 21131
rect 21726 21128 21732 21140
rect 21683 21100 21732 21128
rect 21683 21097 21695 21100
rect 21637 21091 21695 21097
rect 21726 21088 21732 21100
rect 21784 21088 21790 21140
rect 22462 21088 22468 21140
rect 22520 21128 22526 21140
rect 22649 21131 22707 21137
rect 22649 21128 22661 21131
rect 22520 21100 22661 21128
rect 22520 21088 22526 21100
rect 22649 21097 22661 21100
rect 22695 21128 22707 21131
rect 22738 21128 22744 21140
rect 22695 21100 22744 21128
rect 22695 21097 22707 21100
rect 22649 21091 22707 21097
rect 22738 21088 22744 21100
rect 22796 21088 22802 21140
rect 28997 21131 29055 21137
rect 23676 21100 28672 21128
rect 23676 21060 23704 21100
rect 21468 21032 23704 21060
rect 23753 21063 23811 21069
rect 23753 21029 23765 21063
rect 23799 21029 23811 21063
rect 23753 21023 23811 21029
rect 18693 20995 18751 21001
rect 18693 20961 18705 20995
rect 18739 20992 18751 20995
rect 20070 20992 20076 21004
rect 18739 20964 19472 20992
rect 18739 20961 18751 20964
rect 18693 20955 18751 20961
rect 11701 20927 11759 20933
rect 11701 20924 11713 20927
rect 10376 20896 11713 20924
rect 10376 20884 10382 20896
rect 11701 20893 11713 20896
rect 11747 20893 11759 20927
rect 11701 20887 11759 20893
rect 11885 20927 11943 20933
rect 11885 20893 11897 20927
rect 11931 20893 11943 20927
rect 11885 20887 11943 20893
rect 11980 20927 12038 20933
rect 11980 20893 11992 20927
rect 12026 20893 12038 20927
rect 11980 20887 12038 20893
rect 12069 20927 12127 20933
rect 12069 20893 12081 20927
rect 12115 20918 12127 20927
rect 12158 20918 12164 20936
rect 12115 20893 12164 20918
rect 12069 20890 12164 20893
rect 12069 20887 12127 20890
rect 6914 20865 6920 20868
rect 4479 20828 6776 20856
rect 4479 20825 4491 20828
rect 4433 20819 4491 20825
rect 6908 20819 6920 20865
rect 6972 20856 6978 20868
rect 6972 20828 7008 20856
rect 6914 20816 6920 20819
rect 6972 20816 6978 20828
rect 7558 20816 7564 20868
rect 7616 20856 7622 20868
rect 8110 20856 8116 20868
rect 7616 20828 8116 20856
rect 7616 20816 7622 20828
rect 8110 20816 8116 20828
rect 8168 20816 8174 20868
rect 9582 20816 9588 20868
rect 9640 20856 9646 20868
rect 11149 20859 11207 20865
rect 11149 20856 11161 20859
rect 9640 20828 11161 20856
rect 9640 20816 9646 20828
rect 11149 20825 11161 20828
rect 11195 20825 11207 20859
rect 11149 20819 11207 20825
rect 3237 20791 3295 20797
rect 3237 20757 3249 20791
rect 3283 20788 3295 20791
rect 3326 20788 3332 20800
rect 3283 20760 3332 20788
rect 3283 20757 3295 20760
rect 3237 20751 3295 20757
rect 3326 20748 3332 20760
rect 3384 20748 3390 20800
rect 6362 20748 6368 20800
rect 6420 20788 6426 20800
rect 7834 20788 7840 20800
rect 6420 20760 7840 20788
rect 6420 20748 6426 20760
rect 7834 20748 7840 20760
rect 7892 20748 7898 20800
rect 11164 20788 11192 20819
rect 11790 20816 11796 20868
rect 11848 20856 11854 20868
rect 11891 20856 11919 20887
rect 12158 20884 12164 20890
rect 12216 20884 12222 20936
rect 15470 20924 15476 20936
rect 15431 20896 15476 20924
rect 15470 20884 15476 20896
rect 15528 20884 15534 20936
rect 18340 20896 19012 20924
rect 18340 20868 18368 20896
rect 11848 20828 11919 20856
rect 11848 20816 11854 20828
rect 14366 20816 14372 20868
rect 14424 20856 14430 20868
rect 15228 20859 15286 20865
rect 14424 20828 15148 20856
rect 14424 20816 14430 20828
rect 12158 20788 12164 20800
rect 11164 20760 12164 20788
rect 12158 20748 12164 20760
rect 12216 20748 12222 20800
rect 14093 20791 14151 20797
rect 14093 20757 14105 20791
rect 14139 20788 14151 20791
rect 15010 20788 15016 20800
rect 14139 20760 15016 20788
rect 14139 20757 14151 20760
rect 14093 20751 14151 20757
rect 15010 20748 15016 20760
rect 15068 20748 15074 20800
rect 15120 20788 15148 20828
rect 15228 20825 15240 20859
rect 15274 20856 15286 20859
rect 15378 20856 15384 20868
rect 15274 20828 15384 20856
rect 15274 20825 15286 20828
rect 15228 20819 15286 20825
rect 15378 20816 15384 20828
rect 15436 20816 15442 20868
rect 16298 20816 16304 20868
rect 16356 20856 16362 20868
rect 17586 20856 17592 20868
rect 16356 20828 17592 20856
rect 16356 20816 16362 20828
rect 17586 20816 17592 20828
rect 17644 20816 17650 20868
rect 18322 20856 18328 20868
rect 18283 20828 18328 20856
rect 18322 20816 18328 20828
rect 18380 20816 18386 20868
rect 18509 20859 18567 20865
rect 18509 20825 18521 20859
rect 18555 20856 18567 20859
rect 18874 20856 18880 20868
rect 18555 20828 18880 20856
rect 18555 20825 18567 20828
rect 18509 20819 18567 20825
rect 18874 20816 18880 20828
rect 18932 20816 18938 20868
rect 18984 20856 19012 20896
rect 19150 20884 19156 20936
rect 19208 20924 19214 20936
rect 19444 20933 19472 20964
rect 19536 20964 20076 20992
rect 19536 20933 19564 20964
rect 20070 20952 20076 20964
rect 20128 20952 20134 21004
rect 20622 20952 20628 21004
rect 20680 20952 20686 21004
rect 21100 20992 21128 21020
rect 23382 20992 23388 21004
rect 21100 20964 23152 20992
rect 19245 20927 19303 20933
rect 19245 20924 19257 20927
rect 19208 20896 19257 20924
rect 19208 20884 19214 20896
rect 19245 20893 19257 20896
rect 19291 20893 19303 20927
rect 19245 20887 19303 20893
rect 19429 20927 19487 20933
rect 19429 20893 19441 20927
rect 19475 20893 19487 20927
rect 19429 20887 19487 20893
rect 19521 20927 19579 20933
rect 19521 20893 19533 20927
rect 19567 20893 19579 20927
rect 19521 20887 19579 20893
rect 19610 20884 19616 20936
rect 19668 20924 19674 20936
rect 20640 20924 20668 20952
rect 19668 20896 20668 20924
rect 21085 20927 21143 20933
rect 19668 20884 19674 20896
rect 21085 20893 21097 20927
rect 21131 20924 21143 20927
rect 22370 20924 22376 20936
rect 21131 20896 22376 20924
rect 21131 20893 21143 20896
rect 21085 20887 21143 20893
rect 22370 20884 22376 20896
rect 22428 20884 22434 20936
rect 22557 20927 22615 20933
rect 22557 20893 22569 20927
rect 22603 20924 22615 20927
rect 22646 20924 22652 20936
rect 22603 20896 22652 20924
rect 22603 20893 22615 20896
rect 22557 20887 22615 20893
rect 22646 20884 22652 20896
rect 22704 20884 22710 20936
rect 22738 20884 22744 20936
rect 22796 20924 22802 20936
rect 22796 20896 22841 20924
rect 22796 20884 22802 20896
rect 20622 20856 20628 20868
rect 18984 20828 20628 20856
rect 20622 20816 20628 20828
rect 20680 20856 20686 20868
rect 20680 20828 20944 20856
rect 20680 20816 20686 20828
rect 20254 20788 20260 20800
rect 15120 20760 20260 20788
rect 20254 20748 20260 20760
rect 20312 20748 20318 20800
rect 20441 20791 20499 20797
rect 20441 20757 20453 20791
rect 20487 20788 20499 20791
rect 20714 20788 20720 20800
rect 20487 20760 20720 20788
rect 20487 20757 20499 20760
rect 20441 20751 20499 20757
rect 20714 20748 20720 20760
rect 20772 20748 20778 20800
rect 20916 20797 20944 20828
rect 21542 20816 21548 20868
rect 21600 20856 21606 20868
rect 21729 20859 21787 20865
rect 21729 20856 21741 20859
rect 21600 20828 21741 20856
rect 21600 20816 21606 20828
rect 21729 20825 21741 20828
rect 21775 20825 21787 20859
rect 23124 20856 23152 20964
rect 23216 20964 23388 20992
rect 23216 20933 23244 20964
rect 23382 20952 23388 20964
rect 23440 20952 23446 21004
rect 23768 20992 23796 21023
rect 24854 21020 24860 21072
rect 24912 21060 24918 21072
rect 25866 21060 25872 21072
rect 24912 21032 25872 21060
rect 24912 21020 24918 21032
rect 25866 21020 25872 21032
rect 25924 21020 25930 21072
rect 26786 20992 26792 21004
rect 23768 20964 25636 20992
rect 26747 20964 26792 20992
rect 23201 20927 23259 20933
rect 23201 20893 23213 20927
rect 23247 20893 23259 20927
rect 23474 20924 23480 20936
rect 23435 20896 23480 20924
rect 23201 20887 23259 20893
rect 23474 20884 23480 20896
rect 23532 20884 23538 20936
rect 23569 20927 23627 20933
rect 23569 20893 23581 20927
rect 23615 20924 23627 20927
rect 23658 20924 23664 20936
rect 23615 20896 23664 20924
rect 23615 20893 23627 20896
rect 23569 20887 23627 20893
rect 23658 20884 23664 20896
rect 23716 20924 23722 20936
rect 24397 20927 24455 20933
rect 24397 20924 24409 20927
rect 23716 20896 24409 20924
rect 23716 20884 23722 20896
rect 24397 20893 24409 20896
rect 24443 20893 24455 20927
rect 24397 20887 24455 20893
rect 25128 20927 25186 20933
rect 25128 20893 25140 20927
rect 25174 20893 25186 20927
rect 25128 20887 25186 20893
rect 25317 20927 25375 20933
rect 25317 20893 25329 20927
rect 25363 20924 25375 20927
rect 25406 20924 25412 20936
rect 25363 20896 25412 20924
rect 25363 20893 25375 20896
rect 25317 20887 25375 20893
rect 23382 20856 23388 20868
rect 23124 20828 23388 20856
rect 21729 20819 21787 20825
rect 23382 20816 23388 20828
rect 23440 20816 23446 20868
rect 25143 20800 25171 20887
rect 25406 20884 25412 20896
rect 25464 20884 25470 20936
rect 25608 20933 25636 20964
rect 26786 20952 26792 20964
rect 26844 20952 26850 21004
rect 28534 20952 28540 21004
rect 28592 20992 28598 21004
rect 28644 21001 28672 21100
rect 28997 21097 29009 21131
rect 29043 21128 29055 21131
rect 29086 21128 29092 21140
rect 29043 21100 29092 21128
rect 29043 21097 29055 21100
rect 28997 21091 29055 21097
rect 29086 21088 29092 21100
rect 29144 21088 29150 21140
rect 30377 21131 30435 21137
rect 30377 21097 30389 21131
rect 30423 21128 30435 21131
rect 30650 21128 30656 21140
rect 30423 21100 30656 21128
rect 30423 21097 30435 21100
rect 30377 21091 30435 21097
rect 30650 21088 30656 21100
rect 30708 21088 30714 21140
rect 33594 21128 33600 21140
rect 33555 21100 33600 21128
rect 33594 21088 33600 21100
rect 33652 21088 33658 21140
rect 35618 21128 35624 21140
rect 35579 21100 35624 21128
rect 35618 21088 35624 21100
rect 35676 21088 35682 21140
rect 37642 21088 37648 21140
rect 37700 21128 37706 21140
rect 37700 21100 38056 21128
rect 37700 21088 37706 21100
rect 34149 21063 34207 21069
rect 34149 21029 34161 21063
rect 34195 21060 34207 21063
rect 34195 21032 35388 21060
rect 34195 21029 34207 21032
rect 34149 21023 34207 21029
rect 28629 20995 28687 21001
rect 28629 20992 28641 20995
rect 28592 20964 28641 20992
rect 28592 20952 28598 20964
rect 28629 20961 28641 20964
rect 28675 20961 28687 20995
rect 32401 20995 32459 21001
rect 32401 20992 32413 20995
rect 28629 20955 28687 20961
rect 28736 20964 32413 20992
rect 27062 20933 27068 20936
rect 25500 20927 25558 20933
rect 25500 20893 25512 20927
rect 25546 20893 25558 20927
rect 25500 20887 25558 20893
rect 25593 20927 25651 20933
rect 25593 20893 25605 20927
rect 25639 20893 25651 20927
rect 27056 20924 27068 20933
rect 27023 20896 27068 20924
rect 25593 20887 25651 20893
rect 27056 20887 27068 20896
rect 25225 20859 25283 20865
rect 25225 20825 25237 20859
rect 25271 20856 25283 20859
rect 25516 20856 25544 20887
rect 27062 20884 27068 20887
rect 27120 20884 27126 20936
rect 27338 20884 27344 20936
rect 27396 20924 27402 20936
rect 28736 20924 28764 20964
rect 32401 20961 32413 20964
rect 32447 20992 32459 20995
rect 34514 20992 34520 21004
rect 32447 20964 34520 20992
rect 32447 20961 32459 20964
rect 32401 20955 32459 20961
rect 27396 20896 28764 20924
rect 27396 20884 27402 20896
rect 28810 20884 28816 20936
rect 28868 20924 28874 20936
rect 30009 20927 30067 20933
rect 28868 20896 28913 20924
rect 28868 20884 28874 20896
rect 30009 20893 30021 20927
rect 30055 20924 30067 20927
rect 30282 20924 30288 20936
rect 30055 20896 30288 20924
rect 30055 20893 30067 20896
rect 30009 20887 30067 20893
rect 30282 20884 30288 20896
rect 30340 20884 30346 20936
rect 32953 20927 33011 20933
rect 32953 20893 32965 20927
rect 32999 20893 33011 20927
rect 33134 20924 33140 20936
rect 33095 20896 33140 20924
rect 32953 20887 33011 20893
rect 28994 20856 29000 20868
rect 25271 20828 25452 20856
rect 25516 20828 29000 20856
rect 25271 20825 25283 20828
rect 25225 20819 25283 20825
rect 20901 20791 20959 20797
rect 20901 20757 20913 20791
rect 20947 20757 20959 20791
rect 20901 20751 20959 20757
rect 24854 20748 24860 20800
rect 24912 20788 24918 20800
rect 24949 20791 25007 20797
rect 24949 20788 24961 20791
rect 24912 20760 24961 20788
rect 24912 20748 24918 20760
rect 24949 20757 24961 20760
rect 24995 20757 25007 20791
rect 24949 20751 25007 20757
rect 25130 20748 25136 20800
rect 25188 20748 25194 20800
rect 25424 20788 25452 20828
rect 28994 20816 29000 20828
rect 29052 20816 29058 20868
rect 30098 20816 30104 20868
rect 30156 20856 30162 20868
rect 30193 20859 30251 20865
rect 30193 20856 30205 20859
rect 30156 20828 30205 20856
rect 30156 20816 30162 20828
rect 30193 20825 30205 20828
rect 30239 20856 30251 20859
rect 32306 20856 32312 20868
rect 30239 20828 32312 20856
rect 30239 20825 30251 20828
rect 30193 20819 30251 20825
rect 32306 20816 32312 20828
rect 32364 20816 32370 20868
rect 28074 20788 28080 20800
rect 25424 20760 28080 20788
rect 28074 20748 28080 20760
rect 28132 20748 28138 20800
rect 28169 20791 28227 20797
rect 28169 20757 28181 20791
rect 28215 20788 28227 20791
rect 28258 20788 28264 20800
rect 28215 20760 28264 20788
rect 28215 20757 28227 20760
rect 28169 20751 28227 20757
rect 28258 20748 28264 20760
rect 28316 20748 28322 20800
rect 30834 20788 30840 20800
rect 30795 20760 30840 20788
rect 30834 20748 30840 20760
rect 30892 20748 30898 20800
rect 31941 20791 31999 20797
rect 31941 20757 31953 20791
rect 31987 20788 31999 20791
rect 32968 20788 32996 20887
rect 33134 20884 33140 20896
rect 33192 20884 33198 20936
rect 33336 20933 33364 20964
rect 34514 20952 34520 20964
rect 34572 20952 34578 21004
rect 34790 20952 34796 21004
rect 34848 20992 34854 21004
rect 34848 20964 35204 20992
rect 34848 20952 34854 20964
rect 33229 20927 33287 20933
rect 33229 20893 33241 20927
rect 33275 20893 33287 20927
rect 33229 20887 33287 20893
rect 33321 20927 33379 20933
rect 33321 20893 33333 20927
rect 33367 20893 33379 20927
rect 34974 20924 34980 20936
rect 34935 20896 34980 20924
rect 33321 20887 33379 20893
rect 33244 20856 33272 20887
rect 34974 20884 34980 20896
rect 35032 20884 35038 20936
rect 35176 20933 35204 20964
rect 35360 20933 35388 21032
rect 38028 21001 38056 21100
rect 38013 20995 38071 21001
rect 38013 20961 38025 20995
rect 38059 20992 38071 20995
rect 38194 20992 38200 21004
rect 38059 20964 38200 20992
rect 38059 20961 38071 20964
rect 38013 20955 38071 20961
rect 38194 20952 38200 20964
rect 38252 20952 38258 21004
rect 35161 20927 35219 20933
rect 35161 20893 35173 20927
rect 35207 20893 35219 20927
rect 35161 20887 35219 20893
rect 35253 20927 35311 20933
rect 35253 20893 35265 20927
rect 35299 20893 35311 20927
rect 35253 20887 35311 20893
rect 35345 20927 35403 20933
rect 35345 20893 35357 20927
rect 35391 20924 35403 20927
rect 37458 20924 37464 20936
rect 35391 20896 37464 20924
rect 35391 20893 35403 20896
rect 35345 20887 35403 20893
rect 33502 20856 33508 20868
rect 33244 20828 33508 20856
rect 33502 20816 33508 20828
rect 33560 20856 33566 20868
rect 35268 20856 35296 20887
rect 37458 20884 37464 20896
rect 37516 20884 37522 20936
rect 35434 20856 35440 20868
rect 33560 20828 35440 20856
rect 33560 20816 33566 20828
rect 35434 20816 35440 20828
rect 35492 20816 35498 20868
rect 35710 20816 35716 20868
rect 35768 20856 35774 20868
rect 37746 20859 37804 20865
rect 37746 20856 37758 20859
rect 35768 20828 37758 20856
rect 35768 20816 35774 20828
rect 37746 20825 37758 20828
rect 37792 20825 37804 20859
rect 37746 20819 37804 20825
rect 34790 20788 34796 20800
rect 31987 20760 34796 20788
rect 31987 20757 31999 20760
rect 31941 20751 31999 20757
rect 34790 20748 34796 20760
rect 34848 20788 34854 20800
rect 34974 20788 34980 20800
rect 34848 20760 34980 20788
rect 34848 20748 34854 20760
rect 34974 20748 34980 20760
rect 35032 20788 35038 20800
rect 36081 20791 36139 20797
rect 36081 20788 36093 20791
rect 35032 20760 36093 20788
rect 35032 20748 35038 20760
rect 36081 20757 36093 20760
rect 36127 20757 36139 20791
rect 36630 20788 36636 20800
rect 36591 20760 36636 20788
rect 36081 20751 36139 20757
rect 36630 20748 36636 20760
rect 36688 20748 36694 20800
rect 1104 20698 68816 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 68816 20698
rect 1104 20624 68816 20646
rect 6730 20584 6736 20596
rect 4816 20556 6736 20584
rect 2866 20476 2872 20528
rect 2924 20476 2930 20528
rect 4816 20525 4844 20556
rect 6730 20544 6736 20556
rect 6788 20544 6794 20596
rect 7285 20587 7343 20593
rect 7285 20553 7297 20587
rect 7331 20584 7343 20587
rect 7466 20584 7472 20596
rect 7331 20556 7472 20584
rect 7331 20553 7343 20556
rect 7285 20547 7343 20553
rect 7466 20544 7472 20556
rect 7524 20544 7530 20596
rect 7742 20584 7748 20596
rect 7703 20556 7748 20584
rect 7742 20544 7748 20556
rect 7800 20544 7806 20596
rect 10965 20587 11023 20593
rect 10965 20553 10977 20587
rect 11011 20584 11023 20587
rect 11011 20556 12204 20584
rect 11011 20553 11023 20556
rect 10965 20547 11023 20553
rect 4801 20519 4859 20525
rect 4801 20485 4813 20519
rect 4847 20485 4859 20519
rect 4801 20479 4859 20485
rect 5626 20476 5632 20528
rect 5684 20516 5690 20528
rect 6365 20519 6423 20525
rect 6365 20516 6377 20519
rect 5684 20488 6377 20516
rect 5684 20476 5690 20488
rect 6365 20485 6377 20488
rect 6411 20516 6423 20519
rect 11517 20519 11575 20525
rect 11517 20516 11529 20519
rect 6411 20488 8064 20516
rect 6411 20485 6423 20488
rect 6365 20479 6423 20485
rect 1946 20448 1952 20460
rect 1907 20420 1952 20448
rect 1946 20408 1952 20420
rect 2004 20408 2010 20460
rect 2130 20448 2136 20460
rect 2091 20420 2136 20448
rect 2130 20408 2136 20420
rect 2188 20408 2194 20460
rect 2784 20383 2842 20389
rect 2784 20349 2796 20383
rect 2830 20380 2842 20383
rect 2884 20380 2912 20476
rect 3050 20457 3056 20460
rect 3044 20411 3056 20457
rect 3108 20448 3114 20460
rect 4617 20451 4675 20457
rect 3108 20420 3144 20448
rect 3050 20408 3056 20411
rect 3108 20408 3114 20420
rect 4617 20417 4629 20451
rect 4663 20448 4675 20451
rect 4706 20448 4712 20460
rect 4663 20420 4712 20448
rect 4663 20417 4675 20420
rect 4617 20411 4675 20417
rect 4706 20408 4712 20420
rect 4764 20408 4770 20460
rect 8036 20457 8064 20488
rect 10499 20488 11529 20516
rect 10499 20460 10527 20488
rect 11517 20485 11529 20488
rect 11563 20485 11575 20519
rect 11517 20479 11575 20485
rect 11701 20519 11759 20525
rect 11701 20485 11713 20519
rect 11747 20516 11759 20519
rect 12176 20516 12204 20556
rect 15378 20544 15384 20596
rect 15436 20584 15442 20596
rect 15473 20587 15531 20593
rect 15473 20584 15485 20587
rect 15436 20556 15485 20584
rect 15436 20544 15442 20556
rect 15473 20553 15485 20556
rect 15519 20553 15531 20587
rect 16390 20584 16396 20596
rect 15473 20547 15531 20553
rect 16224 20556 16396 20584
rect 12682 20519 12740 20525
rect 12682 20516 12694 20519
rect 11747 20488 12112 20516
rect 12176 20488 12694 20516
rect 11747 20485 11759 20488
rect 11701 20479 11759 20485
rect 7101 20451 7159 20457
rect 7101 20417 7113 20451
rect 7147 20417 7159 20451
rect 7101 20411 7159 20417
rect 8021 20451 8079 20457
rect 8021 20417 8033 20451
rect 8067 20417 8079 20451
rect 8021 20411 8079 20417
rect 8113 20451 8171 20457
rect 8113 20417 8125 20451
rect 8159 20417 8171 20451
rect 8113 20411 8171 20417
rect 8205 20451 8263 20457
rect 8205 20417 8217 20451
rect 8251 20448 8263 20451
rect 8294 20448 8300 20460
rect 8251 20420 8300 20448
rect 8251 20417 8263 20420
rect 8205 20411 8263 20417
rect 2830 20352 2912 20380
rect 6917 20383 6975 20389
rect 2830 20349 2842 20352
rect 2784 20343 2842 20349
rect 6917 20349 6929 20383
rect 6963 20349 6975 20383
rect 7116 20380 7144 20411
rect 8128 20380 8156 20411
rect 8294 20408 8300 20420
rect 8352 20408 8358 20460
rect 8389 20451 8447 20457
rect 8389 20417 8401 20451
rect 8435 20448 8447 20451
rect 8846 20448 8852 20460
rect 8435 20420 8852 20448
rect 8435 20417 8447 20420
rect 8389 20411 8447 20417
rect 8846 20408 8852 20420
rect 8904 20408 8910 20460
rect 10318 20448 10324 20460
rect 10279 20420 10324 20448
rect 10318 20408 10324 20420
rect 10376 20408 10382 20460
rect 10484 20454 10542 20460
rect 10484 20420 10496 20454
rect 10530 20420 10542 20454
rect 10484 20414 10542 20420
rect 10594 20408 10600 20460
rect 10652 20448 10658 20460
rect 10735 20451 10793 20457
rect 10652 20420 10697 20448
rect 10652 20408 10658 20420
rect 10735 20417 10747 20451
rect 10781 20448 10793 20451
rect 11054 20448 11060 20460
rect 10781 20420 11060 20448
rect 10781 20417 10793 20420
rect 10735 20411 10793 20417
rect 11054 20408 11060 20420
rect 11112 20408 11118 20460
rect 11606 20408 11612 20460
rect 11664 20448 11670 20460
rect 11885 20451 11943 20457
rect 11885 20448 11897 20451
rect 11664 20420 11897 20448
rect 11664 20408 11670 20420
rect 11885 20417 11897 20420
rect 11931 20417 11943 20451
rect 12084 20448 12112 20488
rect 12682 20485 12694 20488
rect 12728 20485 12740 20519
rect 16022 20516 16028 20528
rect 12682 20479 12740 20485
rect 15948 20488 16028 20516
rect 15746 20448 15752 20460
rect 12084 20420 13860 20448
rect 15707 20420 15752 20448
rect 11885 20411 11943 20417
rect 8754 20380 8760 20392
rect 7116 20352 8064 20380
rect 8128 20352 8760 20380
rect 6917 20343 6975 20349
rect 4154 20272 4160 20324
rect 4212 20312 4218 20324
rect 5258 20312 5264 20324
rect 4212 20284 5264 20312
rect 4212 20272 4218 20284
rect 5258 20272 5264 20284
rect 5316 20272 5322 20324
rect 5813 20315 5871 20321
rect 5813 20281 5825 20315
rect 5859 20312 5871 20315
rect 6932 20312 6960 20343
rect 7926 20312 7932 20324
rect 5859 20284 7932 20312
rect 5859 20281 5871 20284
rect 5813 20275 5871 20281
rect 7926 20272 7932 20284
rect 7984 20272 7990 20324
rect 8036 20312 8064 20352
rect 8754 20340 8760 20352
rect 8812 20380 8818 20392
rect 10612 20380 10640 20408
rect 12434 20380 12440 20392
rect 8812 20352 10640 20380
rect 12395 20352 12440 20380
rect 8812 20340 8818 20352
rect 12434 20340 12440 20352
rect 12492 20340 12498 20392
rect 13832 20321 13860 20420
rect 15746 20408 15752 20420
rect 15804 20408 15810 20460
rect 15948 20457 15976 20488
rect 16022 20476 16028 20488
rect 16080 20476 16086 20528
rect 16224 20516 16252 20556
rect 16390 20544 16396 20556
rect 16448 20544 16454 20596
rect 20070 20584 20076 20596
rect 17052 20556 20076 20584
rect 17052 20516 17080 20556
rect 20070 20544 20076 20556
rect 20128 20544 20134 20596
rect 20714 20544 20720 20596
rect 20772 20584 20778 20596
rect 22278 20584 22284 20596
rect 20772 20556 22284 20584
rect 20772 20544 20778 20556
rect 22278 20544 22284 20556
rect 22336 20544 22342 20596
rect 22922 20544 22928 20596
rect 22980 20584 22986 20596
rect 24578 20584 24584 20596
rect 22980 20556 24584 20584
rect 22980 20544 22986 20556
rect 24578 20544 24584 20556
rect 24636 20544 24642 20596
rect 25498 20584 25504 20596
rect 25470 20544 25504 20584
rect 25556 20544 25562 20596
rect 27706 20584 27712 20596
rect 27667 20556 27712 20584
rect 27706 20544 27712 20556
rect 27764 20544 27770 20596
rect 28534 20584 28540 20596
rect 28495 20556 28540 20584
rect 28534 20544 28540 20556
rect 28592 20544 28598 20596
rect 35710 20584 35716 20596
rect 28644 20556 35388 20584
rect 35671 20556 35716 20584
rect 17773 20519 17831 20525
rect 17773 20516 17785 20519
rect 16132 20488 16252 20516
rect 16321 20488 17080 20516
rect 16132 20457 16160 20488
rect 15841 20451 15899 20457
rect 15841 20417 15853 20451
rect 15887 20417 15899 20451
rect 15841 20411 15899 20417
rect 15933 20451 15991 20457
rect 15933 20417 15945 20451
rect 15979 20417 15991 20451
rect 15933 20411 15991 20417
rect 16129 20451 16187 20457
rect 16129 20417 16141 20451
rect 16175 20417 16187 20451
rect 16129 20411 16187 20417
rect 15562 20340 15568 20392
rect 15620 20380 15626 20392
rect 15856 20380 15884 20411
rect 16321 20380 16349 20488
rect 16942 20448 16948 20460
rect 16903 20420 16948 20448
rect 16942 20408 16948 20420
rect 17000 20408 17006 20460
rect 17052 20457 17080 20488
rect 17144 20488 17785 20516
rect 17144 20457 17172 20488
rect 17773 20485 17785 20488
rect 17819 20485 17831 20519
rect 18141 20519 18199 20525
rect 18141 20516 18153 20519
rect 17773 20479 17831 20485
rect 17880 20488 18153 20516
rect 17037 20451 17095 20457
rect 17037 20417 17049 20451
rect 17083 20417 17095 20451
rect 17037 20411 17095 20417
rect 17129 20451 17187 20457
rect 17129 20417 17141 20451
rect 17175 20417 17187 20451
rect 17129 20411 17187 20417
rect 17313 20451 17371 20457
rect 17313 20417 17325 20451
rect 17359 20417 17371 20451
rect 17313 20411 17371 20417
rect 15620 20352 16349 20380
rect 15620 20340 15626 20352
rect 16390 20340 16396 20392
rect 16448 20380 16454 20392
rect 17328 20380 17356 20411
rect 17586 20408 17592 20460
rect 17644 20448 17650 20460
rect 17880 20448 17908 20488
rect 18141 20485 18153 20488
rect 18187 20516 18199 20519
rect 18322 20516 18328 20528
rect 18187 20488 18328 20516
rect 18187 20485 18199 20488
rect 18141 20479 18199 20485
rect 18322 20476 18328 20488
rect 18380 20476 18386 20528
rect 23474 20516 23480 20528
rect 23435 20488 23480 20516
rect 23474 20476 23480 20488
rect 23532 20476 23538 20528
rect 23566 20476 23572 20528
rect 23624 20516 23630 20528
rect 23624 20488 23669 20516
rect 23624 20476 23630 20488
rect 17644 20420 17908 20448
rect 17957 20451 18015 20457
rect 17644 20408 17650 20420
rect 17957 20417 17969 20451
rect 18003 20448 18015 20451
rect 18046 20448 18052 20460
rect 18003 20420 18052 20448
rect 18003 20417 18015 20420
rect 17957 20411 18015 20417
rect 18046 20408 18052 20420
rect 18104 20408 18110 20460
rect 18230 20408 18236 20460
rect 18288 20448 18294 20460
rect 20717 20451 20775 20457
rect 18288 20420 20668 20448
rect 18288 20408 18294 20420
rect 19150 20380 19156 20392
rect 16448 20352 19156 20380
rect 16448 20340 16454 20352
rect 19150 20340 19156 20352
rect 19208 20340 19214 20392
rect 19334 20340 19340 20392
rect 19392 20380 19398 20392
rect 20441 20383 20499 20389
rect 20441 20380 20453 20383
rect 19392 20352 20453 20380
rect 19392 20340 19398 20352
rect 20441 20349 20453 20352
rect 20487 20349 20499 20383
rect 20640 20380 20668 20420
rect 20717 20417 20729 20451
rect 20763 20448 20775 20451
rect 21082 20448 21088 20460
rect 20763 20420 21088 20448
rect 20763 20417 20775 20420
rect 20717 20411 20775 20417
rect 21082 20408 21088 20420
rect 21140 20408 21146 20460
rect 23198 20408 23204 20460
rect 23256 20448 23262 20460
rect 23293 20451 23351 20457
rect 23293 20448 23305 20451
rect 23256 20420 23305 20448
rect 23256 20408 23262 20420
rect 23293 20417 23305 20420
rect 23339 20417 23351 20451
rect 23293 20411 23351 20417
rect 23661 20451 23719 20457
rect 23661 20417 23673 20451
rect 23707 20448 23719 20451
rect 23707 20420 23796 20448
rect 23707 20417 23719 20420
rect 23661 20411 23719 20417
rect 21266 20380 21272 20392
rect 20640 20352 21272 20380
rect 20441 20343 20499 20349
rect 21266 20340 21272 20352
rect 21324 20340 21330 20392
rect 8849 20315 8907 20321
rect 8849 20312 8861 20315
rect 8036 20284 8861 20312
rect 8849 20281 8861 20284
rect 8895 20312 8907 20315
rect 13817 20315 13875 20321
rect 8895 20284 10456 20312
rect 8895 20281 8907 20284
rect 8849 20275 8907 20281
rect 1765 20247 1823 20253
rect 1765 20213 1777 20247
rect 1811 20244 1823 20247
rect 2038 20244 2044 20256
rect 1811 20216 2044 20244
rect 1811 20213 1823 20216
rect 1765 20207 1823 20213
rect 2038 20204 2044 20216
rect 2096 20204 2102 20256
rect 4614 20204 4620 20256
rect 4672 20244 4678 20256
rect 4985 20247 5043 20253
rect 4985 20244 4997 20247
rect 4672 20216 4997 20244
rect 4672 20204 4678 20216
rect 4985 20213 4997 20216
rect 5031 20213 5043 20247
rect 4985 20207 5043 20213
rect 7282 20204 7288 20256
rect 7340 20244 7346 20256
rect 9401 20247 9459 20253
rect 9401 20244 9413 20247
rect 7340 20216 9413 20244
rect 7340 20204 7346 20216
rect 9401 20213 9413 20216
rect 9447 20213 9459 20247
rect 10428 20244 10456 20284
rect 13817 20281 13829 20315
rect 13863 20312 13875 20315
rect 15838 20312 15844 20324
rect 13863 20284 15844 20312
rect 13863 20281 13875 20284
rect 13817 20275 13875 20281
rect 15838 20272 15844 20284
rect 15896 20272 15902 20324
rect 20714 20272 20720 20324
rect 20772 20312 20778 20324
rect 22741 20315 22799 20321
rect 22741 20312 22753 20315
rect 20772 20284 22753 20312
rect 20772 20272 20778 20284
rect 22741 20281 22753 20284
rect 22787 20312 22799 20315
rect 23658 20312 23664 20324
rect 22787 20284 23664 20312
rect 22787 20281 22799 20284
rect 22741 20275 22799 20281
rect 23658 20272 23664 20284
rect 23716 20312 23722 20324
rect 23768 20312 23796 20420
rect 25222 20408 25228 20460
rect 25280 20448 25286 20460
rect 25470 20457 25498 20544
rect 25593 20519 25651 20525
rect 25593 20485 25605 20519
rect 25639 20516 25651 20519
rect 28644 20516 28672 20556
rect 30926 20516 30932 20528
rect 25639 20488 28672 20516
rect 30887 20488 30932 20516
rect 25639 20485 25651 20488
rect 25593 20479 25651 20485
rect 30926 20476 30932 20488
rect 30984 20476 30990 20528
rect 34164 20525 34192 20556
rect 34149 20519 34207 20525
rect 34149 20485 34161 20519
rect 34195 20485 34207 20519
rect 34149 20479 34207 20485
rect 34333 20519 34391 20525
rect 34333 20485 34345 20519
rect 34379 20516 34391 20519
rect 35360 20516 35388 20556
rect 35710 20544 35716 20556
rect 35768 20544 35774 20596
rect 36630 20516 36636 20528
rect 34379 20488 35204 20516
rect 35360 20488 36636 20516
rect 34379 20485 34391 20488
rect 34333 20479 34391 20485
rect 25455 20451 25513 20457
rect 25455 20448 25467 20451
rect 25280 20420 25467 20448
rect 25280 20408 25286 20420
rect 25455 20417 25467 20420
rect 25501 20417 25513 20451
rect 25682 20448 25688 20460
rect 25643 20420 25688 20448
rect 25455 20411 25513 20417
rect 25682 20408 25688 20420
rect 25740 20408 25746 20460
rect 25774 20408 25780 20460
rect 25832 20457 25838 20460
rect 25832 20451 25871 20457
rect 25859 20417 25871 20451
rect 25832 20411 25871 20417
rect 25961 20451 26019 20457
rect 25961 20417 25973 20451
rect 26007 20417 26019 20451
rect 25961 20411 26019 20417
rect 27893 20451 27951 20457
rect 27893 20417 27905 20451
rect 27939 20417 27951 20451
rect 27893 20411 27951 20417
rect 28077 20451 28135 20457
rect 28077 20417 28089 20451
rect 28123 20448 28135 20451
rect 28994 20448 29000 20460
rect 28123 20420 29000 20448
rect 28123 20417 28135 20420
rect 28077 20411 28135 20417
rect 25832 20408 25838 20411
rect 25976 20380 26004 20411
rect 23860 20352 26004 20380
rect 27908 20380 27936 20411
rect 28994 20408 29000 20420
rect 29052 20408 29058 20460
rect 29270 20448 29276 20460
rect 29183 20420 29276 20448
rect 29270 20408 29276 20420
rect 29328 20448 29334 20460
rect 29914 20448 29920 20460
rect 29328 20420 29920 20448
rect 29328 20408 29334 20420
rect 29914 20408 29920 20420
rect 29972 20448 29978 20460
rect 31481 20451 31539 20457
rect 31481 20448 31493 20451
rect 29972 20420 31493 20448
rect 29972 20408 29978 20420
rect 31481 20417 31493 20420
rect 31527 20417 31539 20451
rect 31481 20411 31539 20417
rect 31754 20408 31760 20460
rect 31812 20448 31818 20460
rect 33238 20451 33296 20457
rect 33238 20448 33250 20451
rect 31812 20420 33250 20448
rect 31812 20408 31818 20420
rect 33238 20417 33250 20420
rect 33284 20417 33296 20451
rect 33238 20411 33296 20417
rect 33410 20408 33416 20460
rect 33468 20448 33474 20460
rect 33965 20451 34023 20457
rect 33965 20448 33977 20451
rect 33468 20420 33977 20448
rect 33468 20408 33474 20420
rect 33965 20417 33977 20420
rect 34011 20448 34023 20451
rect 34698 20448 34704 20460
rect 34011 20420 34704 20448
rect 34011 20417 34023 20420
rect 33965 20411 34023 20417
rect 34698 20408 34704 20420
rect 34756 20408 34762 20460
rect 34790 20408 34796 20460
rect 34848 20448 34854 20460
rect 35069 20451 35127 20457
rect 35069 20448 35081 20451
rect 34848 20420 35081 20448
rect 34848 20408 34854 20420
rect 35069 20417 35081 20420
rect 35115 20417 35127 20451
rect 35176 20451 35204 20488
rect 36630 20476 36636 20488
rect 36688 20476 36694 20528
rect 35253 20451 35311 20457
rect 35176 20423 35265 20451
rect 35069 20411 35127 20417
rect 35253 20417 35265 20423
rect 35299 20417 35311 20451
rect 35253 20411 35311 20417
rect 35345 20451 35403 20457
rect 35345 20417 35357 20451
rect 35391 20417 35403 20451
rect 35345 20411 35403 20417
rect 35437 20451 35495 20457
rect 35437 20417 35449 20451
rect 35483 20448 35495 20451
rect 35526 20448 35532 20460
rect 35483 20420 35532 20448
rect 35483 20417 35495 20420
rect 35437 20411 35495 20417
rect 28258 20380 28264 20392
rect 27908 20352 28264 20380
rect 23860 20321 23888 20352
rect 28258 20340 28264 20352
rect 28316 20340 28322 20392
rect 33505 20383 33563 20389
rect 33505 20349 33517 20383
rect 33551 20349 33563 20383
rect 35360 20380 35388 20411
rect 35526 20408 35532 20420
rect 35584 20448 35590 20460
rect 36173 20451 36231 20457
rect 36173 20448 36185 20451
rect 35584 20420 36185 20448
rect 35584 20408 35590 20420
rect 36173 20417 36185 20420
rect 36219 20417 36231 20451
rect 38194 20448 38200 20460
rect 38155 20420 38200 20448
rect 36173 20411 36231 20417
rect 38194 20408 38200 20420
rect 38252 20408 38258 20460
rect 38286 20408 38292 20460
rect 38344 20448 38350 20460
rect 38453 20451 38511 20457
rect 38453 20448 38465 20451
rect 38344 20420 38465 20448
rect 38344 20408 38350 20420
rect 38453 20417 38465 20420
rect 38499 20417 38511 20451
rect 38453 20411 38511 20417
rect 35360 20352 35480 20380
rect 33505 20343 33563 20349
rect 23716 20284 23796 20312
rect 23845 20315 23903 20321
rect 23716 20272 23722 20284
rect 23845 20281 23857 20315
rect 23891 20281 23903 20315
rect 23845 20275 23903 20281
rect 24670 20272 24676 20324
rect 24728 20312 24734 20324
rect 26878 20312 26884 20324
rect 24728 20284 26884 20312
rect 24728 20272 24734 20284
rect 26878 20272 26884 20284
rect 26936 20272 26942 20324
rect 31110 20312 31116 20324
rect 30392 20284 31116 20312
rect 12802 20244 12808 20256
rect 10428 20216 12808 20244
rect 9401 20207 9459 20213
rect 12802 20204 12808 20216
rect 12860 20204 12866 20256
rect 15746 20204 15752 20256
rect 15804 20244 15810 20256
rect 16206 20244 16212 20256
rect 15804 20216 16212 20244
rect 15804 20204 15810 20216
rect 16206 20204 16212 20216
rect 16264 20204 16270 20256
rect 16666 20244 16672 20256
rect 16627 20216 16672 20244
rect 16666 20204 16672 20216
rect 16724 20204 16730 20256
rect 18966 20204 18972 20256
rect 19024 20244 19030 20256
rect 19061 20247 19119 20253
rect 19061 20244 19073 20247
rect 19024 20216 19073 20244
rect 19024 20204 19030 20216
rect 19061 20213 19073 20216
rect 19107 20244 19119 20247
rect 19426 20244 19432 20256
rect 19107 20216 19432 20244
rect 19107 20213 19119 20216
rect 19061 20207 19119 20213
rect 19426 20204 19432 20216
rect 19484 20204 19490 20256
rect 19886 20244 19892 20256
rect 19847 20216 19892 20244
rect 19886 20204 19892 20216
rect 19944 20204 19950 20256
rect 21542 20204 21548 20256
rect 21600 20244 21606 20256
rect 21821 20247 21879 20253
rect 21821 20244 21833 20247
rect 21600 20216 21833 20244
rect 21600 20204 21606 20216
rect 21821 20213 21833 20216
rect 21867 20213 21879 20247
rect 21821 20207 21879 20213
rect 23934 20204 23940 20256
rect 23992 20244 23998 20256
rect 25317 20247 25375 20253
rect 25317 20244 25329 20247
rect 23992 20216 25329 20244
rect 23992 20204 23998 20216
rect 25317 20213 25329 20216
rect 25363 20213 25375 20247
rect 25317 20207 25375 20213
rect 25498 20204 25504 20256
rect 25556 20244 25562 20256
rect 30392 20244 30420 20284
rect 31110 20272 31116 20284
rect 31168 20272 31174 20324
rect 33520 20312 33548 20343
rect 35452 20324 35480 20352
rect 34146 20312 34152 20324
rect 33520 20284 34152 20312
rect 34146 20272 34152 20284
rect 34204 20312 34210 20324
rect 35342 20312 35348 20324
rect 34204 20284 35348 20312
rect 34204 20272 34210 20284
rect 35342 20272 35348 20284
rect 35400 20272 35406 20324
rect 35434 20272 35440 20324
rect 35492 20272 35498 20324
rect 37458 20312 37464 20324
rect 37371 20284 37464 20312
rect 37458 20272 37464 20284
rect 37516 20312 37522 20324
rect 38194 20312 38200 20324
rect 37516 20284 38200 20312
rect 37516 20272 37522 20284
rect 38194 20272 38200 20284
rect 38252 20272 38258 20324
rect 25556 20216 30420 20244
rect 25556 20204 25562 20216
rect 30466 20204 30472 20256
rect 30524 20244 30530 20256
rect 32125 20247 32183 20253
rect 32125 20244 32137 20247
rect 30524 20216 32137 20244
rect 30524 20204 30530 20216
rect 32125 20213 32137 20216
rect 32171 20213 32183 20247
rect 32125 20207 32183 20213
rect 37642 20204 37648 20256
rect 37700 20244 37706 20256
rect 39577 20247 39635 20253
rect 39577 20244 39589 20247
rect 37700 20216 39589 20244
rect 37700 20204 37706 20216
rect 39577 20213 39589 20216
rect 39623 20213 39635 20247
rect 39577 20207 39635 20213
rect 1104 20154 68816 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 65654 20154
rect 65706 20102 65718 20154
rect 65770 20102 65782 20154
rect 65834 20102 65846 20154
rect 65898 20102 65910 20154
rect 65962 20102 68816 20154
rect 1104 20080 68816 20102
rect 2501 20043 2559 20049
rect 2501 20009 2513 20043
rect 2547 20040 2559 20043
rect 3050 20040 3056 20052
rect 2547 20012 3056 20040
rect 2547 20009 2559 20012
rect 2501 20003 2559 20009
rect 3050 20000 3056 20012
rect 3108 20000 3114 20052
rect 3142 20000 3148 20052
rect 3200 20040 3206 20052
rect 8386 20040 8392 20052
rect 3200 20012 8392 20040
rect 3200 20000 3206 20012
rect 8386 20000 8392 20012
rect 8444 20000 8450 20052
rect 12434 20000 12440 20052
rect 12492 20040 12498 20052
rect 13081 20043 13139 20049
rect 13081 20040 13093 20043
rect 12492 20012 13093 20040
rect 12492 20000 12498 20012
rect 13081 20009 13093 20012
rect 13127 20009 13139 20043
rect 13081 20003 13139 20009
rect 15565 20043 15623 20049
rect 15565 20009 15577 20043
rect 15611 20040 15623 20043
rect 16022 20040 16028 20052
rect 15611 20012 16028 20040
rect 15611 20009 15623 20012
rect 15565 20003 15623 20009
rect 16022 20000 16028 20012
rect 16080 20000 16086 20052
rect 16114 20000 16120 20052
rect 16172 20040 16178 20052
rect 19245 20043 19303 20049
rect 16172 20012 18644 20040
rect 16172 20000 16178 20012
rect 2314 19972 2320 19984
rect 1872 19944 2320 19972
rect 1872 19848 1900 19944
rect 2314 19932 2320 19944
rect 2372 19972 2378 19984
rect 4338 19972 4344 19984
rect 2372 19944 4344 19972
rect 2372 19932 2378 19944
rect 4338 19932 4344 19944
rect 4396 19972 4402 19984
rect 5350 19972 5356 19984
rect 4396 19944 5356 19972
rect 4396 19932 4402 19944
rect 5350 19932 5356 19944
rect 5408 19932 5414 19984
rect 10597 19975 10655 19981
rect 10597 19941 10609 19975
rect 10643 19972 10655 19975
rect 16482 19972 16488 19984
rect 10643 19944 16488 19972
rect 10643 19941 10655 19944
rect 10597 19935 10655 19941
rect 2774 19864 2780 19916
rect 2832 19904 2838 19916
rect 2961 19907 3019 19913
rect 2961 19904 2973 19907
rect 2832 19876 2973 19904
rect 2832 19864 2838 19876
rect 2961 19873 2973 19876
rect 3007 19904 3019 19907
rect 3050 19904 3056 19916
rect 3007 19876 3056 19904
rect 3007 19873 3019 19876
rect 2961 19867 3019 19873
rect 3050 19864 3056 19876
rect 3108 19864 3114 19916
rect 4062 19864 4068 19916
rect 4120 19904 4126 19916
rect 5445 19907 5503 19913
rect 5445 19904 5457 19907
rect 4120 19876 5457 19904
rect 4120 19864 4126 19876
rect 5445 19873 5457 19876
rect 5491 19873 5503 19907
rect 5445 19867 5503 19873
rect 1854 19836 1860 19848
rect 1815 19808 1860 19836
rect 1854 19796 1860 19808
rect 1912 19796 1918 19848
rect 2038 19836 2044 19848
rect 1999 19808 2044 19836
rect 2038 19796 2044 19808
rect 2096 19796 2102 19848
rect 2133 19839 2191 19845
rect 2133 19805 2145 19839
rect 2179 19805 2191 19839
rect 2133 19799 2191 19805
rect 2225 19839 2283 19845
rect 2225 19805 2237 19839
rect 2271 19836 2283 19839
rect 2406 19836 2412 19848
rect 2271 19808 2412 19836
rect 2271 19805 2283 19808
rect 2225 19799 2283 19805
rect 2148 19768 2176 19799
rect 2406 19796 2412 19808
rect 2464 19796 2470 19848
rect 4338 19836 4344 19848
rect 4299 19808 4344 19836
rect 4338 19796 4344 19808
rect 4396 19796 4402 19848
rect 4522 19836 4528 19848
rect 4483 19808 4528 19836
rect 4522 19796 4528 19808
rect 4580 19796 4586 19848
rect 4617 19839 4675 19845
rect 4617 19805 4629 19839
rect 4663 19805 4675 19839
rect 4617 19799 4675 19805
rect 4709 19839 4767 19845
rect 4709 19805 4721 19839
rect 4755 19836 4767 19839
rect 5074 19836 5080 19848
rect 4755 19808 5080 19836
rect 4755 19805 4767 19808
rect 4709 19799 4767 19805
rect 4632 19768 4660 19799
rect 5074 19796 5080 19808
rect 5132 19836 5138 19848
rect 5132 19808 7604 19836
rect 5132 19796 5138 19808
rect 7576 19780 7604 19808
rect 8294 19796 8300 19848
rect 8352 19836 8358 19848
rect 9214 19836 9220 19848
rect 8352 19808 9220 19836
rect 8352 19796 8358 19808
rect 9214 19796 9220 19808
rect 9272 19796 9278 19848
rect 2148 19740 4660 19768
rect 4985 19771 5043 19777
rect 2240 19712 2268 19740
rect 4985 19737 4997 19771
rect 5031 19768 5043 19771
rect 5690 19771 5748 19777
rect 5690 19768 5702 19771
rect 5031 19740 5702 19768
rect 5031 19737 5043 19740
rect 4985 19731 5043 19737
rect 5690 19737 5702 19740
rect 5736 19737 5748 19771
rect 5690 19731 5748 19737
rect 7282 19728 7288 19780
rect 7340 19768 7346 19780
rect 7377 19771 7435 19777
rect 7377 19768 7389 19771
rect 7340 19740 7389 19768
rect 7340 19728 7346 19740
rect 7377 19737 7389 19740
rect 7423 19737 7435 19771
rect 7558 19768 7564 19780
rect 7519 19740 7564 19768
rect 7377 19731 7435 19737
rect 7558 19728 7564 19740
rect 7616 19728 7622 19780
rect 8018 19768 8024 19780
rect 7979 19740 8024 19768
rect 8018 19728 8024 19740
rect 8076 19728 8082 19780
rect 8205 19771 8263 19777
rect 8205 19737 8217 19771
rect 8251 19768 8263 19771
rect 8251 19740 9076 19768
rect 8251 19737 8263 19740
rect 8205 19731 8263 19737
rect 2222 19660 2228 19712
rect 2280 19660 2286 19712
rect 6730 19660 6736 19712
rect 6788 19700 6794 19712
rect 6825 19703 6883 19709
rect 6825 19700 6837 19703
rect 6788 19672 6837 19700
rect 6788 19660 6794 19672
rect 6825 19669 6837 19672
rect 6871 19669 6883 19703
rect 6825 19663 6883 19669
rect 8389 19703 8447 19709
rect 8389 19669 8401 19703
rect 8435 19700 8447 19703
rect 8478 19700 8484 19712
rect 8435 19672 8484 19700
rect 8435 19669 8447 19672
rect 8389 19663 8447 19669
rect 8478 19660 8484 19672
rect 8536 19660 8542 19712
rect 9048 19700 9076 19740
rect 9122 19728 9128 19780
rect 9180 19768 9186 19780
rect 9462 19771 9520 19777
rect 9462 19768 9474 19771
rect 9180 19740 9474 19768
rect 9180 19728 9186 19740
rect 9462 19737 9474 19740
rect 9508 19737 9520 19771
rect 9462 19731 9520 19737
rect 10612 19700 10640 19935
rect 16482 19932 16488 19944
rect 16540 19932 16546 19984
rect 18616 19972 18644 20012
rect 19245 20009 19257 20043
rect 19291 20040 19303 20043
rect 25682 20040 25688 20052
rect 19291 20012 25688 20040
rect 19291 20009 19303 20012
rect 19245 20003 19303 20009
rect 25682 20000 25688 20012
rect 25740 20000 25746 20052
rect 26418 20000 26424 20052
rect 26476 20040 26482 20052
rect 27522 20040 27528 20052
rect 26476 20012 27528 20040
rect 26476 20000 26482 20012
rect 27522 20000 27528 20012
rect 27580 20040 27586 20052
rect 30190 20040 30196 20052
rect 27580 20012 30196 20040
rect 27580 20000 27586 20012
rect 30190 20000 30196 20012
rect 30248 20000 30254 20052
rect 31754 20000 31760 20052
rect 31812 20040 31818 20052
rect 31812 20012 31857 20040
rect 31812 20000 31818 20012
rect 19886 19972 19892 19984
rect 18616 19944 19892 19972
rect 19886 19932 19892 19944
rect 19944 19972 19950 19984
rect 27801 19975 27859 19981
rect 27801 19972 27813 19975
rect 19944 19944 20668 19972
rect 19944 19932 19950 19944
rect 15470 19864 15476 19916
rect 15528 19904 15534 19916
rect 16853 19907 16911 19913
rect 16853 19904 16865 19907
rect 15528 19876 16865 19904
rect 15528 19864 15534 19876
rect 16853 19873 16865 19876
rect 16899 19873 16911 19907
rect 16853 19867 16911 19873
rect 19150 19864 19156 19916
rect 19208 19904 19214 19916
rect 19208 19876 20300 19904
rect 19208 19864 19214 19876
rect 20272 19848 20300 19876
rect 11330 19836 11336 19848
rect 11243 19808 11336 19836
rect 11330 19796 11336 19808
rect 11388 19836 11394 19848
rect 11793 19839 11851 19845
rect 11793 19836 11805 19839
rect 11388 19808 11805 19836
rect 11388 19796 11394 19808
rect 11793 19805 11805 19808
rect 11839 19836 11851 19839
rect 12342 19836 12348 19848
rect 11839 19808 12348 19836
rect 11839 19805 11851 19808
rect 11793 19799 11851 19805
rect 12342 19796 12348 19808
rect 12400 19796 12406 19848
rect 15010 19796 15016 19848
rect 15068 19836 15074 19848
rect 15381 19839 15439 19845
rect 15381 19836 15393 19839
rect 15068 19808 15393 19836
rect 15068 19796 15074 19808
rect 15381 19805 15393 19808
rect 15427 19805 15439 19839
rect 16206 19836 16212 19848
rect 16167 19808 16212 19836
rect 15381 19799 15439 19805
rect 16206 19796 16212 19808
rect 16264 19796 16270 19848
rect 16666 19796 16672 19848
rect 16724 19836 16730 19848
rect 17109 19839 17167 19845
rect 17109 19836 17121 19839
rect 16724 19808 17121 19836
rect 16724 19796 16730 19808
rect 17109 19805 17121 19808
rect 17155 19805 17167 19839
rect 19426 19836 19432 19848
rect 19387 19808 19432 19836
rect 17109 19799 17167 19805
rect 19426 19796 19432 19808
rect 19484 19796 19490 19848
rect 19518 19796 19524 19848
rect 19576 19836 19582 19848
rect 19794 19836 19800 19848
rect 19576 19808 19621 19836
rect 19755 19808 19800 19836
rect 19576 19796 19582 19808
rect 19794 19796 19800 19808
rect 19852 19796 19858 19848
rect 20254 19836 20260 19848
rect 20215 19808 20260 19836
rect 20254 19796 20260 19808
rect 20312 19796 20318 19848
rect 20438 19836 20444 19848
rect 20399 19808 20444 19836
rect 20438 19796 20444 19808
rect 20496 19796 20502 19848
rect 20640 19845 20668 19944
rect 23124 19944 27813 19972
rect 22741 19907 22799 19913
rect 22741 19873 22753 19907
rect 22787 19904 22799 19907
rect 22922 19904 22928 19916
rect 22787 19876 22928 19904
rect 22787 19873 22799 19876
rect 22741 19867 22799 19873
rect 22922 19864 22928 19876
rect 22980 19864 22986 19916
rect 20533 19839 20591 19845
rect 20533 19805 20545 19839
rect 20579 19805 20591 19839
rect 20533 19799 20591 19805
rect 20625 19839 20683 19845
rect 20625 19805 20637 19839
rect 20671 19836 20683 19839
rect 21174 19836 21180 19848
rect 20671 19808 21180 19836
rect 20671 19805 20683 19808
rect 20625 19799 20683 19805
rect 14918 19728 14924 19780
rect 14976 19768 14982 19780
rect 15197 19771 15255 19777
rect 15197 19768 15209 19771
rect 14976 19740 15209 19768
rect 14976 19728 14982 19740
rect 15197 19737 15209 19740
rect 15243 19768 15255 19771
rect 17586 19768 17592 19780
rect 15243 19740 17592 19768
rect 15243 19737 15255 19740
rect 15197 19731 15255 19737
rect 17586 19728 17592 19740
rect 17644 19728 17650 19780
rect 19150 19728 19156 19780
rect 19208 19768 19214 19780
rect 19613 19771 19671 19777
rect 19613 19768 19625 19771
rect 19208 19740 19625 19768
rect 19208 19728 19214 19740
rect 19613 19737 19625 19740
rect 19659 19737 19671 19771
rect 19613 19731 19671 19737
rect 20070 19728 20076 19780
rect 20128 19768 20134 19780
rect 20548 19768 20576 19799
rect 21174 19796 21180 19808
rect 21232 19796 21238 19848
rect 21266 19796 21272 19848
rect 21324 19836 21330 19848
rect 23124 19836 23152 19944
rect 27801 19941 27813 19944
rect 27847 19972 27859 19975
rect 27847 19944 28764 19972
rect 27847 19941 27859 19944
rect 27801 19935 27859 19941
rect 24762 19904 24768 19916
rect 23400 19876 24768 19904
rect 23400 19845 23428 19876
rect 24762 19864 24768 19876
rect 24820 19864 24826 19916
rect 25130 19864 25136 19916
rect 25188 19904 25194 19916
rect 25498 19904 25504 19916
rect 25188 19876 25504 19904
rect 25188 19864 25194 19876
rect 25498 19864 25504 19876
rect 25556 19864 25562 19916
rect 27430 19904 27436 19916
rect 26712 19876 27436 19904
rect 21324 19808 23152 19836
rect 23201 19839 23259 19845
rect 21324 19796 21330 19808
rect 23201 19805 23213 19839
rect 23247 19805 23259 19839
rect 23201 19799 23259 19805
rect 23385 19839 23443 19845
rect 23385 19805 23397 19839
rect 23431 19805 23443 19839
rect 23385 19799 23443 19805
rect 23477 19839 23535 19845
rect 23477 19805 23489 19839
rect 23523 19805 23535 19839
rect 23477 19799 23535 19805
rect 23569 19839 23627 19845
rect 23569 19805 23581 19839
rect 23615 19836 23627 19839
rect 23658 19836 23664 19848
rect 23615 19808 23664 19836
rect 23615 19805 23627 19808
rect 23569 19799 23627 19805
rect 20128 19740 20576 19768
rect 20901 19771 20959 19777
rect 20128 19728 20134 19740
rect 20901 19737 20913 19771
rect 20947 19768 20959 19771
rect 22474 19771 22532 19777
rect 22474 19768 22486 19771
rect 20947 19740 22486 19768
rect 20947 19737 20959 19740
rect 20901 19731 20959 19737
rect 22474 19737 22486 19740
rect 22520 19737 22532 19771
rect 22474 19731 22532 19737
rect 22646 19728 22652 19780
rect 22704 19768 22710 19780
rect 23216 19768 23244 19799
rect 22704 19740 23244 19768
rect 22704 19728 22710 19740
rect 9048 19672 10640 19700
rect 18138 19660 18144 19712
rect 18196 19700 18202 19712
rect 18233 19703 18291 19709
rect 18233 19700 18245 19703
rect 18196 19672 18245 19700
rect 18196 19660 18202 19672
rect 18233 19669 18245 19672
rect 18279 19669 18291 19703
rect 18233 19663 18291 19669
rect 20530 19660 20536 19712
rect 20588 19700 20594 19712
rect 21361 19703 21419 19709
rect 21361 19700 21373 19703
rect 20588 19672 21373 19700
rect 20588 19660 20594 19672
rect 21361 19669 21373 19672
rect 21407 19669 21419 19703
rect 21361 19663 21419 19669
rect 22370 19660 22376 19712
rect 22428 19700 22434 19712
rect 23492 19700 23520 19799
rect 23658 19796 23664 19808
rect 23716 19796 23722 19848
rect 24397 19839 24455 19845
rect 24397 19805 24409 19839
rect 24443 19836 24455 19839
rect 24486 19836 24492 19848
rect 24443 19808 24492 19836
rect 24443 19805 24455 19808
rect 24397 19799 24455 19805
rect 24486 19796 24492 19808
rect 24544 19796 24550 19848
rect 25222 19845 25228 19848
rect 25220 19836 25228 19845
rect 25183 19808 25228 19836
rect 25220 19799 25228 19808
rect 25222 19796 25228 19799
rect 25280 19796 25286 19848
rect 25406 19836 25412 19848
rect 25367 19808 25412 19836
rect 25406 19796 25412 19808
rect 25464 19796 25470 19848
rect 25592 19839 25650 19845
rect 25592 19805 25604 19839
rect 25638 19805 25650 19839
rect 25592 19799 25650 19805
rect 23845 19771 23903 19777
rect 23845 19737 23857 19771
rect 23891 19768 23903 19771
rect 24946 19768 24952 19780
rect 23891 19740 24952 19768
rect 23891 19737 23903 19740
rect 23845 19731 23903 19737
rect 24946 19728 24952 19740
rect 25004 19728 25010 19780
rect 25317 19771 25375 19777
rect 25317 19737 25329 19771
rect 25363 19737 25375 19771
rect 25608 19768 25636 19799
rect 25682 19796 25688 19848
rect 25740 19836 25746 19848
rect 26418 19836 26424 19848
rect 25740 19808 25785 19836
rect 26379 19808 26424 19836
rect 25740 19796 25746 19808
rect 26418 19796 26424 19808
rect 26476 19796 26482 19848
rect 26602 19836 26608 19848
rect 26563 19808 26608 19836
rect 26602 19796 26608 19808
rect 26660 19796 26666 19848
rect 26712 19845 26740 19876
rect 27430 19864 27436 19876
rect 27488 19904 27494 19916
rect 27488 19876 28672 19904
rect 27488 19864 27494 19876
rect 26697 19839 26755 19845
rect 26697 19805 26709 19839
rect 26743 19805 26755 19839
rect 26697 19799 26755 19805
rect 26789 19839 26847 19845
rect 26789 19805 26801 19839
rect 26835 19805 26847 19839
rect 26789 19799 26847 19805
rect 25958 19768 25964 19780
rect 25608 19740 25964 19768
rect 25317 19731 25375 19737
rect 22428 19672 23520 19700
rect 24581 19703 24639 19709
rect 22428 19660 22434 19672
rect 24581 19669 24593 19703
rect 24627 19700 24639 19703
rect 24670 19700 24676 19712
rect 24627 19672 24676 19700
rect 24627 19669 24639 19672
rect 24581 19663 24639 19669
rect 24670 19660 24676 19672
rect 24728 19660 24734 19712
rect 25038 19700 25044 19712
rect 24999 19672 25044 19700
rect 25038 19660 25044 19672
rect 25096 19660 25102 19712
rect 25332 19700 25360 19731
rect 25958 19728 25964 19740
rect 26016 19728 26022 19780
rect 26142 19728 26148 19780
rect 26200 19768 26206 19780
rect 26804 19768 26832 19799
rect 27522 19796 27528 19848
rect 27580 19836 27586 19848
rect 28353 19839 28411 19845
rect 28353 19836 28365 19839
rect 27580 19808 28365 19836
rect 27580 19796 27586 19808
rect 28353 19805 28365 19808
rect 28399 19805 28411 19839
rect 28534 19836 28540 19848
rect 28495 19808 28540 19836
rect 28353 19799 28411 19805
rect 28534 19796 28540 19808
rect 28592 19796 28598 19848
rect 28644 19845 28672 19876
rect 28736 19845 28764 19944
rect 28994 19932 29000 19984
rect 29052 19972 29058 19984
rect 29733 19975 29791 19981
rect 29733 19972 29745 19975
rect 29052 19944 29745 19972
rect 29052 19932 29058 19944
rect 29733 19941 29745 19944
rect 29779 19972 29791 19975
rect 30282 19972 30288 19984
rect 29779 19944 30288 19972
rect 29779 19941 29791 19944
rect 29733 19935 29791 19941
rect 30282 19932 30288 19944
rect 30340 19932 30346 19984
rect 35621 19975 35679 19981
rect 35621 19941 35633 19975
rect 35667 19941 35679 19975
rect 35621 19935 35679 19941
rect 35636 19904 35664 19935
rect 28920 19876 35664 19904
rect 28629 19839 28687 19845
rect 28629 19805 28641 19839
rect 28675 19805 28687 19839
rect 28629 19799 28687 19805
rect 28721 19839 28779 19845
rect 28721 19805 28733 19839
rect 28767 19805 28779 19839
rect 28721 19799 28779 19805
rect 26200 19740 26832 19768
rect 26896 19740 28488 19768
rect 26200 19728 26206 19740
rect 26896 19700 26924 19740
rect 27062 19700 27068 19712
rect 25332 19672 26924 19700
rect 27023 19672 27068 19700
rect 27062 19660 27068 19672
rect 27120 19660 27126 19712
rect 28460 19700 28488 19740
rect 28920 19700 28948 19876
rect 29086 19796 29092 19848
rect 29144 19836 29150 19848
rect 29549 19839 29607 19845
rect 29549 19836 29561 19839
rect 29144 19808 29561 19836
rect 29144 19796 29150 19808
rect 29549 19805 29561 19808
rect 29595 19805 29607 19839
rect 30282 19836 30288 19848
rect 30243 19808 30288 19836
rect 29549 19799 29607 19805
rect 30282 19796 30288 19808
rect 30340 19796 30346 19848
rect 31113 19839 31171 19845
rect 31113 19836 31125 19839
rect 30392 19808 31125 19836
rect 30190 19728 30196 19780
rect 30248 19768 30254 19780
rect 30392 19768 30420 19808
rect 31113 19805 31125 19808
rect 31159 19805 31171 19839
rect 31113 19799 31171 19805
rect 31297 19839 31355 19845
rect 31297 19805 31309 19839
rect 31343 19805 31355 19839
rect 31297 19799 31355 19805
rect 30248 19740 30420 19768
rect 30248 19728 30254 19740
rect 30466 19728 30472 19780
rect 30524 19768 30530 19780
rect 30653 19771 30711 19777
rect 30524 19740 30569 19768
rect 30524 19728 30530 19740
rect 30653 19737 30665 19771
rect 30699 19768 30711 19771
rect 31312 19768 31340 19799
rect 31386 19796 31392 19848
rect 31444 19836 31450 19848
rect 34900 19845 34928 19876
rect 31527 19839 31585 19845
rect 31444 19808 31489 19836
rect 31444 19796 31450 19808
rect 31527 19805 31539 19839
rect 31573 19836 31585 19839
rect 32217 19839 32275 19845
rect 32217 19836 32229 19839
rect 31573 19808 32229 19836
rect 31573 19805 31585 19808
rect 31527 19799 31585 19805
rect 30699 19740 31340 19768
rect 30699 19737 30711 19740
rect 30653 19731 30711 19737
rect 28460 19672 28948 19700
rect 28997 19703 29055 19709
rect 28997 19669 29009 19703
rect 29043 19700 29055 19703
rect 29178 19700 29184 19712
rect 29043 19672 29184 19700
rect 29043 19669 29055 19672
rect 28997 19663 29055 19669
rect 29178 19660 29184 19672
rect 29236 19660 29242 19712
rect 30374 19660 30380 19712
rect 30432 19700 30438 19712
rect 31726 19700 31754 19808
rect 32217 19805 32229 19808
rect 32263 19805 32275 19839
rect 32217 19799 32275 19805
rect 34885 19839 34943 19845
rect 34885 19805 34897 19839
rect 34931 19805 34943 19839
rect 34885 19799 34943 19805
rect 35342 19796 35348 19848
rect 35400 19836 35406 19848
rect 37001 19839 37059 19845
rect 37001 19836 37013 19839
rect 35400 19808 37013 19836
rect 35400 19796 35406 19808
rect 37001 19805 37013 19808
rect 37047 19836 37059 19839
rect 39022 19836 39028 19848
rect 37047 19808 39028 19836
rect 37047 19805 37059 19808
rect 37001 19799 37059 19805
rect 39022 19796 39028 19808
rect 39080 19796 39086 19848
rect 68094 19836 68100 19848
rect 68055 19808 68100 19836
rect 68094 19796 68100 19808
rect 68152 19796 68158 19848
rect 34698 19768 34704 19780
rect 34659 19740 34704 19768
rect 34698 19728 34704 19740
rect 34756 19728 34762 19780
rect 35802 19728 35808 19780
rect 35860 19768 35866 19780
rect 36734 19771 36792 19777
rect 36734 19768 36746 19771
rect 35860 19740 36746 19768
rect 35860 19728 35866 19740
rect 36734 19737 36746 19740
rect 36780 19737 36792 19771
rect 37458 19768 37464 19780
rect 37419 19740 37464 19768
rect 36734 19731 36792 19737
rect 37458 19728 37464 19740
rect 37516 19728 37522 19780
rect 37642 19768 37648 19780
rect 37603 19740 37648 19768
rect 37642 19728 37648 19740
rect 37700 19728 37706 19780
rect 30432 19672 31754 19700
rect 34149 19703 34207 19709
rect 30432 19660 30438 19672
rect 34149 19669 34161 19703
rect 34195 19700 34207 19703
rect 34790 19700 34796 19712
rect 34195 19672 34796 19700
rect 34195 19669 34207 19672
rect 34149 19663 34207 19669
rect 34790 19660 34796 19672
rect 34848 19660 34854 19712
rect 35069 19703 35127 19709
rect 35069 19669 35081 19703
rect 35115 19700 35127 19703
rect 35250 19700 35256 19712
rect 35115 19672 35256 19700
rect 35115 19669 35127 19672
rect 35069 19663 35127 19669
rect 35250 19660 35256 19672
rect 35308 19660 35314 19712
rect 37734 19660 37740 19712
rect 37792 19700 37798 19712
rect 37829 19703 37887 19709
rect 37829 19700 37841 19703
rect 37792 19672 37841 19700
rect 37792 19660 37798 19672
rect 37829 19669 37841 19672
rect 37875 19669 37887 19703
rect 37829 19663 37887 19669
rect 1104 19610 68816 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 68816 19610
rect 1104 19536 68816 19558
rect 1673 19499 1731 19505
rect 1673 19465 1685 19499
rect 1719 19496 1731 19499
rect 2406 19496 2412 19508
rect 1719 19468 2412 19496
rect 1719 19465 1731 19468
rect 1673 19459 1731 19465
rect 2406 19456 2412 19468
rect 2464 19456 2470 19508
rect 2682 19456 2688 19508
rect 2740 19496 2746 19508
rect 5626 19496 5632 19508
rect 2740 19468 5632 19496
rect 2740 19456 2746 19468
rect 5626 19456 5632 19468
rect 5684 19456 5690 19508
rect 8478 19456 8484 19508
rect 8536 19456 8542 19508
rect 9122 19496 9128 19508
rect 9083 19468 9128 19496
rect 9122 19456 9128 19468
rect 9180 19456 9186 19508
rect 16761 19499 16819 19505
rect 16761 19496 16773 19499
rect 15580 19468 16773 19496
rect 2222 19388 2228 19440
rect 2280 19428 2286 19440
rect 2777 19431 2835 19437
rect 2280 19400 2452 19428
rect 2280 19388 2286 19400
rect 1854 19320 1860 19372
rect 1912 19360 1918 19372
rect 2133 19363 2191 19369
rect 2133 19360 2145 19363
rect 1912 19332 2145 19360
rect 1912 19320 1918 19332
rect 2133 19329 2145 19332
rect 2179 19329 2191 19363
rect 2314 19360 2320 19372
rect 2275 19332 2320 19360
rect 2133 19323 2191 19329
rect 2314 19320 2320 19332
rect 2372 19320 2378 19372
rect 2424 19369 2452 19400
rect 2777 19397 2789 19431
rect 2823 19428 2835 19431
rect 3666 19431 3724 19437
rect 3666 19428 3678 19431
rect 2823 19400 3678 19428
rect 2823 19397 2835 19400
rect 2777 19391 2835 19397
rect 3666 19397 3678 19400
rect 3712 19397 3724 19431
rect 8496 19428 8524 19456
rect 8496 19400 8616 19428
rect 3666 19391 3724 19397
rect 2409 19363 2467 19369
rect 2409 19329 2421 19363
rect 2455 19329 2467 19363
rect 2409 19323 2467 19329
rect 2501 19363 2559 19369
rect 2501 19329 2513 19363
rect 2547 19360 2559 19363
rect 3234 19360 3240 19372
rect 2547 19332 3240 19360
rect 2547 19329 2559 19332
rect 2501 19323 2559 19329
rect 3234 19320 3240 19332
rect 3292 19320 3298 19372
rect 3418 19320 3424 19372
rect 3476 19360 3482 19372
rect 4062 19360 4068 19372
rect 3476 19332 4068 19360
rect 3476 19320 3482 19332
rect 4062 19320 4068 19332
rect 4120 19320 4126 19372
rect 7098 19320 7104 19372
rect 7156 19360 7162 19372
rect 7285 19363 7343 19369
rect 7285 19360 7297 19363
rect 7156 19332 7297 19360
rect 7156 19320 7162 19332
rect 7285 19329 7297 19332
rect 7331 19329 7343 19363
rect 8478 19360 8484 19372
rect 8439 19332 8484 19360
rect 7285 19323 7343 19329
rect 8478 19320 8484 19332
rect 8536 19320 8542 19372
rect 8588 19360 8616 19400
rect 9214 19388 9220 19440
rect 9272 19428 9278 19440
rect 10318 19428 10324 19440
rect 9272 19400 10324 19428
rect 9272 19388 9278 19400
rect 10318 19388 10324 19400
rect 10376 19428 10382 19440
rect 12158 19428 12164 19440
rect 10376 19400 12164 19428
rect 10376 19388 10382 19400
rect 12158 19388 12164 19400
rect 12216 19428 12222 19440
rect 14918 19428 14924 19440
rect 12216 19400 12388 19428
rect 14879 19400 14924 19428
rect 12216 19388 12222 19400
rect 8644 19363 8702 19369
rect 8644 19360 8656 19363
rect 8588 19332 8656 19360
rect 8644 19329 8656 19332
rect 8690 19329 8702 19363
rect 8644 19323 8702 19329
rect 8754 19320 8760 19372
rect 8812 19360 8818 19372
rect 12360 19369 12388 19400
rect 14918 19388 14924 19400
rect 14976 19388 14982 19440
rect 8895 19363 8953 19369
rect 8812 19332 8857 19360
rect 8812 19320 8818 19332
rect 8895 19329 8907 19363
rect 8941 19329 8953 19363
rect 8895 19323 8953 19329
rect 12345 19363 12403 19369
rect 12345 19329 12357 19363
rect 12391 19329 12403 19363
rect 12345 19323 12403 19329
rect 6549 19295 6607 19301
rect 6549 19261 6561 19295
rect 6595 19292 6607 19295
rect 7006 19292 7012 19304
rect 6595 19264 7012 19292
rect 6595 19261 6607 19264
rect 6549 19255 6607 19261
rect 7006 19252 7012 19264
rect 7064 19252 7070 19304
rect 7466 19252 7472 19304
rect 7524 19292 7530 19304
rect 8386 19292 8392 19304
rect 7524 19264 8392 19292
rect 7524 19252 7530 19264
rect 8386 19252 8392 19264
rect 8444 19292 8450 19304
rect 8910 19292 8938 19323
rect 14458 19320 14464 19372
rect 14516 19360 14522 19372
rect 14737 19363 14795 19369
rect 14737 19360 14749 19363
rect 14516 19332 14749 19360
rect 14516 19320 14522 19332
rect 14737 19329 14749 19332
rect 14783 19329 14795 19363
rect 15580 19363 15608 19468
rect 16761 19465 16773 19468
rect 16807 19496 16819 19499
rect 16850 19496 16856 19508
rect 16807 19468 16856 19496
rect 16807 19465 16819 19468
rect 16761 19459 16819 19465
rect 16850 19456 16856 19468
rect 16908 19496 16914 19508
rect 17494 19496 17500 19508
rect 16908 19468 17500 19496
rect 16908 19456 16914 19468
rect 17494 19456 17500 19468
rect 17552 19456 17558 19508
rect 20254 19456 20260 19508
rect 20312 19496 20318 19508
rect 20312 19468 20759 19496
rect 20312 19456 20318 19468
rect 16482 19388 16488 19440
rect 16540 19428 16546 19440
rect 19245 19431 19303 19437
rect 19245 19428 19257 19431
rect 16540 19400 19257 19428
rect 16540 19388 16546 19400
rect 19245 19397 19257 19400
rect 19291 19397 19303 19431
rect 19245 19391 19303 19397
rect 20349 19431 20407 19437
rect 20349 19397 20361 19431
rect 20395 19428 20407 19431
rect 20622 19428 20628 19440
rect 20395 19400 20628 19428
rect 20395 19397 20407 19400
rect 20349 19391 20407 19397
rect 20622 19388 20628 19400
rect 20680 19388 20686 19440
rect 20731 19428 20759 19468
rect 22738 19456 22744 19508
rect 22796 19496 22802 19508
rect 22971 19499 23029 19505
rect 22971 19496 22983 19499
rect 22796 19468 22983 19496
rect 22796 19456 22802 19468
rect 22971 19465 22983 19468
rect 23017 19465 23029 19499
rect 22971 19459 23029 19465
rect 26142 19456 26148 19508
rect 26200 19496 26206 19508
rect 26237 19499 26295 19505
rect 26237 19496 26249 19499
rect 26200 19468 26249 19496
rect 26200 19456 26206 19468
rect 26237 19465 26249 19468
rect 26283 19465 26295 19499
rect 26237 19459 26295 19465
rect 28534 19456 28540 19508
rect 28592 19496 28598 19508
rect 29454 19496 29460 19508
rect 28592 19468 29460 19496
rect 28592 19456 28598 19468
rect 29454 19456 29460 19468
rect 29512 19456 29518 19508
rect 30190 19456 30196 19508
rect 30248 19496 30254 19508
rect 30469 19499 30527 19505
rect 30469 19496 30481 19499
rect 30248 19468 30481 19496
rect 30248 19456 30254 19468
rect 30469 19465 30481 19468
rect 30515 19465 30527 19499
rect 35802 19496 35808 19508
rect 35763 19468 35808 19496
rect 30469 19459 30527 19465
rect 35802 19456 35808 19468
rect 35860 19456 35866 19508
rect 38197 19499 38255 19505
rect 38197 19465 38209 19499
rect 38243 19496 38255 19499
rect 38286 19496 38292 19508
rect 38243 19468 38292 19496
rect 38243 19465 38255 19468
rect 38197 19459 38255 19465
rect 38286 19456 38292 19468
rect 38344 19456 38350 19508
rect 30926 19428 30932 19440
rect 20731 19400 24716 19428
rect 15657 19363 15715 19369
rect 15580 19335 15669 19363
rect 14737 19323 14795 19329
rect 15657 19329 15669 19335
rect 15703 19329 15715 19363
rect 15657 19323 15715 19329
rect 15749 19363 15807 19369
rect 15841 19366 15899 19372
rect 15841 19363 15853 19366
rect 15749 19329 15761 19363
rect 15795 19329 15807 19363
rect 15749 19323 15807 19329
rect 15837 19332 15853 19363
rect 15887 19332 15899 19366
rect 15837 19326 15899 19332
rect 16025 19363 16083 19369
rect 16025 19329 16037 19363
rect 16071 19360 16083 19363
rect 16390 19360 16396 19372
rect 16071 19332 16396 19360
rect 16071 19329 16083 19332
rect 9677 19295 9735 19301
rect 9677 19292 9689 19295
rect 8444 19264 9689 19292
rect 8444 19252 8450 19264
rect 9677 19261 9689 19264
rect 9723 19261 9735 19295
rect 9677 19255 9735 19261
rect 12621 19295 12679 19301
rect 12621 19261 12633 19295
rect 12667 19292 12679 19295
rect 14553 19295 14611 19301
rect 12667 19264 13124 19292
rect 12667 19261 12679 19264
rect 12621 19255 12679 19261
rect 9030 19184 9036 19236
rect 9088 19224 9094 19236
rect 10229 19227 10287 19233
rect 10229 19224 10241 19227
rect 9088 19196 10241 19224
rect 9088 19184 9094 19196
rect 10229 19193 10241 19196
rect 10275 19224 10287 19227
rect 12986 19224 12992 19236
rect 10275 19196 12992 19224
rect 10275 19193 10287 19196
rect 10229 19187 10287 19193
rect 12986 19184 12992 19196
rect 13044 19184 13050 19236
rect 13096 19168 13124 19264
rect 14553 19261 14565 19295
rect 14599 19292 14611 19295
rect 14599 19264 15194 19292
rect 14599 19261 14611 19264
rect 14553 19255 14611 19261
rect 15166 19224 15194 19264
rect 15562 19252 15568 19304
rect 15620 19292 15626 19304
rect 15764 19292 15792 19323
rect 15620 19264 15792 19292
rect 15620 19252 15626 19264
rect 15837 19224 15865 19326
rect 16025 19323 16083 19329
rect 16390 19320 16396 19332
rect 16448 19320 16454 19372
rect 18966 19360 18972 19372
rect 18927 19332 18972 19360
rect 18966 19320 18972 19332
rect 19024 19320 19030 19372
rect 19150 19360 19156 19372
rect 19111 19332 19156 19360
rect 19150 19320 19156 19332
rect 19208 19320 19214 19372
rect 19337 19363 19395 19369
rect 19337 19329 19349 19363
rect 19383 19360 19395 19363
rect 19426 19360 19432 19372
rect 19383 19332 19432 19360
rect 19383 19329 19395 19332
rect 19337 19323 19395 19329
rect 19426 19320 19432 19332
rect 19484 19320 19490 19372
rect 20530 19360 20536 19372
rect 19996 19332 20536 19360
rect 17310 19292 17316 19304
rect 17271 19264 17316 19292
rect 17310 19252 17316 19264
rect 17368 19252 17374 19304
rect 18046 19252 18052 19304
rect 18104 19292 18110 19304
rect 19996 19292 20024 19332
rect 20530 19320 20536 19332
rect 20588 19320 20594 19372
rect 24688 19369 24716 19400
rect 26988 19400 30932 19428
rect 26988 19372 27016 19400
rect 24673 19363 24731 19369
rect 24673 19329 24685 19363
rect 24719 19329 24731 19363
rect 26970 19360 26976 19372
rect 26883 19332 26976 19360
rect 24673 19323 24731 19329
rect 26970 19320 26976 19332
rect 27028 19320 27034 19372
rect 27062 19320 27068 19372
rect 27120 19360 27126 19372
rect 29104 19369 29132 19400
rect 30926 19388 30932 19400
rect 30984 19388 30990 19440
rect 31110 19388 31116 19440
rect 31168 19428 31174 19440
rect 31297 19431 31355 19437
rect 31297 19428 31309 19431
rect 31168 19400 31309 19428
rect 31168 19388 31174 19400
rect 31297 19397 31309 19400
rect 31343 19428 31355 19431
rect 31343 19400 31754 19428
rect 31343 19397 31355 19400
rect 31297 19391 31355 19397
rect 27229 19363 27287 19369
rect 27229 19360 27241 19363
rect 27120 19332 27241 19360
rect 27120 19320 27126 19332
rect 27229 19329 27241 19332
rect 27275 19329 27287 19363
rect 27229 19323 27287 19329
rect 29089 19363 29147 19369
rect 29089 19329 29101 19363
rect 29135 19329 29147 19363
rect 29089 19323 29147 19329
rect 29178 19320 29184 19372
rect 29236 19360 29242 19372
rect 29345 19363 29403 19369
rect 29345 19360 29357 19363
rect 29236 19332 29357 19360
rect 29236 19320 29242 19332
rect 29345 19329 29357 19332
rect 29391 19329 29403 19363
rect 29345 19323 29403 19329
rect 18104 19264 20024 19292
rect 18104 19252 18110 19264
rect 20438 19252 20444 19304
rect 20496 19292 20502 19304
rect 20717 19295 20775 19301
rect 20717 19292 20729 19295
rect 20496 19264 20729 19292
rect 20496 19252 20502 19264
rect 20717 19261 20729 19264
rect 20763 19261 20775 19295
rect 21174 19292 21180 19304
rect 21135 19264 21180 19292
rect 20717 19255 20775 19261
rect 21174 19252 21180 19264
rect 21232 19252 21238 19304
rect 21358 19252 21364 19304
rect 21416 19292 21422 19304
rect 22741 19295 22799 19301
rect 22741 19292 22753 19295
rect 21416 19264 22753 19292
rect 21416 19252 21422 19264
rect 22741 19261 22753 19264
rect 22787 19261 22799 19295
rect 22741 19255 22799 19261
rect 24949 19295 25007 19301
rect 24949 19261 24961 19295
rect 24995 19292 25007 19295
rect 25130 19292 25136 19304
rect 24995 19264 25136 19292
rect 24995 19261 25007 19264
rect 24949 19255 25007 19261
rect 25130 19252 25136 19264
rect 25188 19252 25194 19304
rect 31726 19292 31754 19400
rect 33502 19388 33508 19440
rect 33560 19428 33566 19440
rect 33560 19400 35480 19428
rect 33560 19388 33566 19400
rect 33870 19320 33876 19372
rect 33928 19360 33934 19372
rect 34434 19363 34492 19369
rect 34434 19360 34446 19363
rect 33928 19332 34446 19360
rect 33928 19320 33934 19332
rect 34434 19329 34446 19332
rect 34480 19329 34492 19363
rect 34434 19323 34492 19329
rect 34790 19320 34796 19372
rect 34848 19360 34854 19372
rect 35158 19360 35164 19372
rect 34848 19332 35164 19360
rect 34848 19320 34854 19332
rect 35158 19320 35164 19332
rect 35216 19320 35222 19372
rect 35250 19320 35256 19372
rect 35308 19360 35314 19372
rect 35452 19369 35480 19400
rect 35345 19363 35403 19369
rect 35345 19360 35357 19363
rect 35308 19332 35357 19360
rect 35308 19320 35314 19332
rect 35345 19329 35357 19332
rect 35391 19329 35403 19363
rect 35345 19323 35403 19329
rect 35437 19363 35495 19369
rect 35437 19329 35449 19363
rect 35483 19329 35495 19363
rect 35437 19323 35495 19329
rect 35529 19363 35587 19369
rect 35529 19329 35541 19363
rect 35575 19360 35587 19363
rect 35710 19360 35716 19372
rect 35575 19332 35716 19360
rect 35575 19329 35587 19332
rect 35529 19323 35587 19329
rect 35710 19320 35716 19332
rect 35768 19320 35774 19372
rect 37550 19360 37556 19372
rect 37511 19332 37556 19360
rect 37550 19320 37556 19332
rect 37608 19320 37614 19372
rect 37734 19360 37740 19372
rect 37695 19332 37740 19360
rect 37734 19320 37740 19332
rect 37792 19320 37798 19372
rect 37829 19363 37887 19369
rect 37829 19329 37841 19363
rect 37875 19329 37887 19363
rect 37829 19323 37887 19329
rect 37921 19363 37979 19369
rect 37921 19329 37933 19363
rect 37967 19360 37979 19363
rect 38194 19360 38200 19372
rect 37967 19332 38200 19360
rect 37967 19329 37979 19332
rect 37921 19323 37979 19329
rect 33134 19292 33140 19304
rect 31726 19264 33140 19292
rect 33134 19252 33140 19264
rect 33192 19252 33198 19304
rect 34701 19295 34759 19301
rect 34701 19261 34713 19295
rect 34747 19292 34759 19295
rect 34747 19264 35388 19292
rect 34747 19261 34759 19264
rect 34701 19255 34759 19261
rect 35360 19236 35388 19264
rect 37366 19252 37372 19304
rect 37424 19292 37430 19304
rect 37844 19292 37872 19323
rect 38194 19320 38200 19332
rect 38252 19320 38258 19372
rect 39206 19320 39212 19372
rect 39264 19360 39270 19372
rect 39373 19363 39431 19369
rect 39373 19360 39385 19363
rect 39264 19332 39385 19360
rect 39264 19320 39270 19332
rect 39373 19329 39385 19332
rect 39419 19329 39431 19363
rect 39373 19323 39431 19329
rect 37424 19264 37872 19292
rect 37424 19252 37430 19264
rect 39022 19252 39028 19304
rect 39080 19292 39086 19304
rect 39117 19295 39175 19301
rect 39117 19292 39129 19295
rect 39080 19264 39129 19292
rect 39080 19252 39086 19264
rect 39117 19261 39129 19264
rect 39163 19261 39175 19295
rect 39117 19255 39175 19261
rect 15166 19196 15865 19224
rect 16390 19184 16396 19236
rect 16448 19224 16454 19236
rect 22830 19224 22836 19236
rect 16448 19196 22836 19224
rect 16448 19184 16454 19196
rect 22830 19184 22836 19196
rect 22888 19184 22894 19236
rect 31481 19227 31539 19233
rect 31481 19193 31493 19227
rect 31527 19224 31539 19227
rect 33686 19224 33692 19236
rect 31527 19196 33692 19224
rect 31527 19193 31539 19196
rect 31481 19187 31539 19193
rect 33686 19184 33692 19196
rect 33744 19184 33750 19236
rect 35342 19184 35348 19236
rect 35400 19184 35406 19236
rect 4801 19159 4859 19165
rect 4801 19125 4813 19159
rect 4847 19156 4859 19159
rect 5166 19156 5172 19168
rect 4847 19128 5172 19156
rect 4847 19125 4859 19128
rect 4801 19119 4859 19125
rect 5166 19116 5172 19128
rect 5224 19116 5230 19168
rect 13078 19156 13084 19168
rect 13039 19128 13084 19156
rect 13078 19116 13084 19128
rect 13136 19116 13142 19168
rect 15378 19156 15384 19168
rect 15339 19128 15384 19156
rect 15378 19116 15384 19128
rect 15436 19116 15442 19168
rect 19521 19159 19579 19165
rect 19521 19125 19533 19159
rect 19567 19156 19579 19159
rect 20622 19156 20628 19168
rect 19567 19128 20628 19156
rect 19567 19125 19579 19128
rect 19521 19119 19579 19125
rect 20622 19116 20628 19128
rect 20680 19116 20686 19168
rect 22281 19159 22339 19165
rect 22281 19125 22293 19159
rect 22327 19156 22339 19159
rect 23658 19156 23664 19168
rect 22327 19128 23664 19156
rect 22327 19125 22339 19128
rect 22281 19119 22339 19125
rect 23658 19116 23664 19128
rect 23716 19116 23722 19168
rect 28350 19156 28356 19168
rect 28311 19128 28356 19156
rect 28350 19116 28356 19128
rect 28408 19116 28414 19168
rect 33318 19156 33324 19168
rect 33279 19128 33324 19156
rect 33318 19116 33324 19128
rect 33376 19116 33382 19168
rect 35158 19116 35164 19168
rect 35216 19156 35222 19168
rect 35618 19156 35624 19168
rect 35216 19128 35624 19156
rect 35216 19116 35222 19128
rect 35618 19116 35624 19128
rect 35676 19156 35682 19168
rect 36265 19159 36323 19165
rect 36265 19156 36277 19159
rect 35676 19128 36277 19156
rect 35676 19116 35682 19128
rect 36265 19125 36277 19128
rect 36311 19125 36323 19159
rect 36265 19119 36323 19125
rect 37918 19116 37924 19168
rect 37976 19156 37982 19168
rect 40497 19159 40555 19165
rect 40497 19156 40509 19159
rect 37976 19128 40509 19156
rect 37976 19116 37982 19128
rect 40497 19125 40509 19128
rect 40543 19125 40555 19159
rect 40497 19119 40555 19125
rect 1104 19066 68816 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 65654 19066
rect 65706 19014 65718 19066
rect 65770 19014 65782 19066
rect 65834 19014 65846 19066
rect 65898 19014 65910 19066
rect 65962 19014 68816 19066
rect 1104 18992 68816 19014
rect 2314 18912 2320 18964
rect 2372 18952 2378 18964
rect 2501 18955 2559 18961
rect 2501 18952 2513 18955
rect 2372 18924 2513 18952
rect 2372 18912 2378 18924
rect 2501 18921 2513 18924
rect 2547 18921 2559 18955
rect 2501 18915 2559 18921
rect 3053 18955 3111 18961
rect 3053 18921 3065 18955
rect 3099 18952 3111 18955
rect 3234 18952 3240 18964
rect 3099 18924 3240 18952
rect 3099 18921 3111 18924
rect 3053 18915 3111 18921
rect 3234 18912 3240 18924
rect 3292 18912 3298 18964
rect 7006 18912 7012 18964
rect 7064 18952 7070 18964
rect 7064 18924 12940 18952
rect 7064 18912 7070 18924
rect 12912 18884 12940 18924
rect 12986 18912 12992 18964
rect 13044 18952 13050 18964
rect 15838 18952 15844 18964
rect 13044 18924 15844 18952
rect 13044 18912 13050 18924
rect 15838 18912 15844 18924
rect 15896 18952 15902 18964
rect 20714 18952 20720 18964
rect 15896 18924 20720 18952
rect 15896 18912 15902 18924
rect 20714 18912 20720 18924
rect 20772 18912 20778 18964
rect 20993 18955 21051 18961
rect 20993 18921 21005 18955
rect 21039 18952 21051 18955
rect 21266 18952 21272 18964
rect 21039 18924 21272 18952
rect 21039 18921 21051 18924
rect 20993 18915 21051 18921
rect 21266 18912 21272 18924
rect 21324 18952 21330 18964
rect 24486 18952 24492 18964
rect 21324 18924 24492 18952
rect 21324 18912 21330 18924
rect 24486 18912 24492 18924
rect 24544 18912 24550 18964
rect 26602 18912 26608 18964
rect 26660 18952 26666 18964
rect 27341 18955 27399 18961
rect 27341 18952 27353 18955
rect 26660 18924 27353 18952
rect 26660 18912 26666 18924
rect 27341 18921 27353 18924
rect 27387 18921 27399 18955
rect 27341 18915 27399 18921
rect 29454 18912 29460 18964
rect 29512 18952 29518 18964
rect 29549 18955 29607 18961
rect 29549 18952 29561 18955
rect 29512 18924 29561 18952
rect 29512 18912 29518 18924
rect 29549 18921 29561 18924
rect 29595 18921 29607 18955
rect 29549 18915 29607 18921
rect 34514 18912 34520 18964
rect 34572 18952 34578 18964
rect 37090 18952 37096 18964
rect 34572 18924 37096 18952
rect 34572 18912 34578 18924
rect 37090 18912 37096 18924
rect 37148 18952 37154 18964
rect 38930 18952 38936 18964
rect 37148 18924 38936 18952
rect 37148 18912 37154 18924
rect 38930 18912 38936 18924
rect 38988 18912 38994 18964
rect 39206 18952 39212 18964
rect 39167 18924 39212 18952
rect 39206 18912 39212 18924
rect 39264 18912 39270 18964
rect 14366 18884 14372 18896
rect 12912 18856 14372 18884
rect 14366 18844 14372 18856
rect 14424 18844 14430 18896
rect 18322 18844 18328 18896
rect 18380 18884 18386 18896
rect 19150 18884 19156 18896
rect 18380 18856 19156 18884
rect 18380 18844 18386 18856
rect 19150 18844 19156 18856
rect 19208 18884 19214 18896
rect 19208 18856 19564 18884
rect 19208 18844 19214 18856
rect 6641 18819 6699 18825
rect 6641 18785 6653 18819
rect 6687 18816 6699 18819
rect 7098 18816 7104 18828
rect 6687 18788 7104 18816
rect 6687 18785 6699 18788
rect 6641 18779 6699 18785
rect 7098 18776 7104 18788
rect 7156 18776 7162 18828
rect 7469 18819 7527 18825
rect 7469 18785 7481 18819
rect 7515 18816 7527 18819
rect 8941 18819 8999 18825
rect 8941 18816 8953 18819
rect 7515 18788 8953 18816
rect 7515 18785 7527 18788
rect 7469 18779 7527 18785
rect 8941 18785 8953 18788
rect 8987 18816 8999 18819
rect 9674 18816 9680 18828
rect 8987 18788 9680 18816
rect 8987 18785 8999 18788
rect 8941 18779 8999 18785
rect 9674 18776 9680 18788
rect 9732 18776 9738 18828
rect 18690 18816 18696 18828
rect 15580 18788 18460 18816
rect 2130 18748 2136 18760
rect 2091 18720 2136 18748
rect 2130 18708 2136 18720
rect 2188 18708 2194 18760
rect 4982 18708 4988 18760
rect 5040 18748 5046 18760
rect 6365 18751 6423 18757
rect 6365 18748 6377 18751
rect 5040 18720 6377 18748
rect 5040 18708 5046 18720
rect 6365 18717 6377 18720
rect 6411 18717 6423 18751
rect 6365 18711 6423 18717
rect 7377 18751 7435 18757
rect 7377 18717 7389 18751
rect 7423 18717 7435 18751
rect 7377 18711 7435 18717
rect 7561 18751 7619 18757
rect 7561 18717 7573 18751
rect 7607 18748 7619 18751
rect 7834 18748 7840 18760
rect 7607 18720 7840 18748
rect 7607 18717 7619 18720
rect 7561 18711 7619 18717
rect 2317 18683 2375 18689
rect 2317 18649 2329 18683
rect 2363 18680 2375 18683
rect 5166 18680 5172 18692
rect 2363 18652 5172 18680
rect 2363 18649 2375 18652
rect 2317 18643 2375 18649
rect 5166 18640 5172 18652
rect 5224 18640 5230 18692
rect 5353 18683 5411 18689
rect 5353 18649 5365 18683
rect 5399 18680 5411 18683
rect 7392 18680 7420 18711
rect 7834 18708 7840 18720
rect 7892 18708 7898 18760
rect 7926 18708 7932 18760
rect 7984 18748 7990 18760
rect 8021 18751 8079 18757
rect 8021 18748 8033 18751
rect 7984 18720 8033 18748
rect 7984 18708 7990 18720
rect 8021 18717 8033 18720
rect 8067 18717 8079 18751
rect 8021 18711 8079 18717
rect 8205 18751 8263 18757
rect 8205 18717 8217 18751
rect 8251 18717 8263 18751
rect 8205 18711 8263 18717
rect 8220 18680 8248 18711
rect 8754 18708 8760 18760
rect 8812 18748 8818 18760
rect 9217 18751 9275 18757
rect 9217 18748 9229 18751
rect 8812 18720 9229 18748
rect 8812 18708 8818 18720
rect 9217 18717 9229 18720
rect 9263 18717 9275 18751
rect 9217 18711 9275 18717
rect 10229 18751 10287 18757
rect 10229 18717 10241 18751
rect 10275 18717 10287 18751
rect 10962 18748 10968 18760
rect 10923 18720 10968 18748
rect 10229 18711 10287 18717
rect 5399 18652 8248 18680
rect 5399 18649 5411 18652
rect 5353 18643 5411 18649
rect 8220 18612 8248 18652
rect 8389 18683 8447 18689
rect 8389 18649 8401 18683
rect 8435 18680 8447 18683
rect 8846 18680 8852 18692
rect 8435 18652 8852 18680
rect 8435 18649 8447 18652
rect 8389 18643 8447 18649
rect 8846 18640 8852 18652
rect 8904 18680 8910 18692
rect 10244 18680 10272 18711
rect 10962 18708 10968 18720
rect 11020 18708 11026 18760
rect 12434 18708 12440 18760
rect 12492 18748 12498 18760
rect 15470 18748 15476 18760
rect 12492 18720 15476 18748
rect 12492 18708 12498 18720
rect 15470 18708 15476 18720
rect 15528 18708 15534 18760
rect 8904 18652 10272 18680
rect 11232 18683 11290 18689
rect 8904 18640 8910 18652
rect 11232 18649 11244 18683
rect 11278 18680 11290 18683
rect 11514 18680 11520 18692
rect 11278 18652 11520 18680
rect 11278 18649 11290 18652
rect 11232 18643 11290 18649
rect 11514 18640 11520 18652
rect 11572 18640 11578 18692
rect 12618 18680 12624 18692
rect 11624 18652 12624 18680
rect 9030 18612 9036 18624
rect 8220 18584 9036 18612
rect 9030 18572 9036 18584
rect 9088 18572 9094 18624
rect 10413 18615 10471 18621
rect 10413 18581 10425 18615
rect 10459 18612 10471 18615
rect 10502 18612 10508 18624
rect 10459 18584 10508 18612
rect 10459 18581 10471 18584
rect 10413 18575 10471 18581
rect 10502 18572 10508 18584
rect 10560 18612 10566 18624
rect 11624 18612 11652 18652
rect 12618 18640 12624 18652
rect 12676 18680 12682 18692
rect 12805 18683 12863 18689
rect 12805 18680 12817 18683
rect 12676 18652 12817 18680
rect 12676 18640 12682 18652
rect 12805 18649 12817 18652
rect 12851 18649 12863 18683
rect 12805 18643 12863 18649
rect 12989 18683 13047 18689
rect 12989 18649 13001 18683
rect 13035 18680 13047 18683
rect 15228 18683 15286 18689
rect 13035 18652 14596 18680
rect 13035 18649 13047 18652
rect 12989 18643 13047 18649
rect 10560 18584 11652 18612
rect 12345 18615 12403 18621
rect 10560 18572 10566 18584
rect 12345 18581 12357 18615
rect 12391 18612 12403 18615
rect 13004 18612 13032 18643
rect 13170 18612 13176 18624
rect 12391 18584 13032 18612
rect 13131 18584 13176 18612
rect 12391 18581 12403 18584
rect 12345 18575 12403 18581
rect 13170 18572 13176 18584
rect 13228 18572 13234 18624
rect 14093 18615 14151 18621
rect 14093 18581 14105 18615
rect 14139 18612 14151 18615
rect 14458 18612 14464 18624
rect 14139 18584 14464 18612
rect 14139 18581 14151 18584
rect 14093 18575 14151 18581
rect 14458 18572 14464 18584
rect 14516 18572 14522 18624
rect 14568 18612 14596 18652
rect 15228 18649 15240 18683
rect 15274 18680 15286 18683
rect 15378 18680 15384 18692
rect 15274 18652 15384 18680
rect 15274 18649 15286 18652
rect 15228 18643 15286 18649
rect 15378 18640 15384 18652
rect 15436 18640 15442 18692
rect 15580 18612 15608 18788
rect 16390 18748 16396 18760
rect 16351 18720 16396 18748
rect 16390 18708 16396 18720
rect 16448 18708 16454 18760
rect 16666 18748 16672 18760
rect 16627 18720 16672 18748
rect 16666 18708 16672 18720
rect 16724 18708 16730 18760
rect 16758 18708 16764 18760
rect 16816 18748 16822 18760
rect 16816 18720 16861 18748
rect 16816 18708 16822 18720
rect 17310 18708 17316 18760
rect 17368 18748 17374 18760
rect 17494 18748 17500 18760
rect 17368 18720 17500 18748
rect 17368 18708 17374 18720
rect 17494 18708 17500 18720
rect 17552 18708 17558 18760
rect 18046 18708 18052 18760
rect 18104 18748 18110 18760
rect 18141 18751 18199 18757
rect 18141 18748 18153 18751
rect 18104 18720 18153 18748
rect 18104 18708 18110 18720
rect 18141 18717 18153 18720
rect 18187 18717 18199 18751
rect 18322 18748 18328 18760
rect 18283 18720 18328 18748
rect 18141 18711 18199 18717
rect 18322 18708 18328 18720
rect 18380 18708 18386 18760
rect 18432 18757 18460 18788
rect 18524 18788 18696 18816
rect 18524 18757 18552 18788
rect 18690 18776 18696 18788
rect 18748 18816 18754 18828
rect 19426 18816 19432 18828
rect 18748 18788 19432 18816
rect 18748 18776 18754 18788
rect 19426 18776 19432 18788
rect 19484 18776 19490 18828
rect 19536 18825 19564 18856
rect 34606 18844 34612 18896
rect 34664 18884 34670 18896
rect 35069 18887 35127 18893
rect 35069 18884 35081 18887
rect 34664 18856 35081 18884
rect 34664 18844 34670 18856
rect 35069 18853 35081 18856
rect 35115 18884 35127 18887
rect 35710 18884 35716 18896
rect 35115 18856 35716 18884
rect 35115 18853 35127 18856
rect 35069 18847 35127 18853
rect 35710 18844 35716 18856
rect 35768 18884 35774 18896
rect 37274 18884 37280 18896
rect 35768 18856 37280 18884
rect 35768 18844 35774 18856
rect 37274 18844 37280 18856
rect 37332 18844 37338 18896
rect 19521 18819 19579 18825
rect 19521 18785 19533 18819
rect 19567 18785 19579 18819
rect 19521 18779 19579 18785
rect 20254 18776 20260 18828
rect 20312 18816 20318 18828
rect 21358 18816 21364 18828
rect 20312 18788 21364 18816
rect 20312 18776 20318 18788
rect 18417 18751 18475 18757
rect 18417 18717 18429 18751
rect 18463 18717 18475 18751
rect 18417 18711 18475 18717
rect 18509 18751 18567 18757
rect 18509 18717 18521 18751
rect 18555 18717 18567 18751
rect 18509 18711 18567 18717
rect 19245 18751 19303 18757
rect 19245 18717 19257 18751
rect 19291 18748 19303 18751
rect 19334 18748 19340 18760
rect 19291 18720 19340 18748
rect 19291 18717 19303 18720
rect 19245 18711 19303 18717
rect 15746 18640 15752 18692
rect 15804 18680 15810 18692
rect 16577 18683 16635 18689
rect 16577 18680 16589 18683
rect 15804 18652 16589 18680
rect 15804 18640 15810 18652
rect 16577 18649 16589 18652
rect 16623 18680 16635 18683
rect 19260 18680 19288 18711
rect 19334 18708 19340 18720
rect 19392 18708 19398 18760
rect 19978 18708 19984 18760
rect 20036 18748 20042 18760
rect 20438 18748 20444 18760
rect 20036 18720 20444 18748
rect 20036 18708 20042 18720
rect 20438 18708 20444 18720
rect 20496 18748 20502 18760
rect 20824 18757 20852 18788
rect 21358 18776 21364 18788
rect 21416 18776 21422 18828
rect 21634 18776 21640 18828
rect 21692 18816 21698 18828
rect 22833 18819 22891 18825
rect 22833 18816 22845 18819
rect 21692 18788 22845 18816
rect 21692 18776 21698 18788
rect 20625 18751 20683 18757
rect 20625 18748 20637 18751
rect 20496 18720 20637 18748
rect 20496 18708 20502 18720
rect 20625 18717 20637 18720
rect 20671 18717 20683 18751
rect 20625 18711 20683 18717
rect 20809 18751 20867 18757
rect 20809 18717 20821 18751
rect 20855 18717 20867 18751
rect 20809 18711 20867 18717
rect 21174 18708 21180 18760
rect 21232 18748 21238 18760
rect 21836 18757 21864 18788
rect 22833 18785 22845 18788
rect 22879 18785 22891 18819
rect 22833 18779 22891 18785
rect 25961 18819 26019 18825
rect 25961 18785 25973 18819
rect 26007 18816 26019 18819
rect 26970 18816 26976 18828
rect 26007 18788 26976 18816
rect 26007 18785 26019 18788
rect 25961 18779 26019 18785
rect 26970 18776 26976 18788
rect 27028 18776 27034 18828
rect 28905 18819 28963 18825
rect 28905 18785 28917 18819
rect 28951 18816 28963 18819
rect 32309 18819 32367 18825
rect 28951 18788 30328 18816
rect 28951 18785 28963 18788
rect 28905 18779 28963 18785
rect 21729 18751 21787 18757
rect 21729 18748 21741 18751
rect 21232 18720 21741 18748
rect 21232 18708 21238 18720
rect 21729 18717 21741 18720
rect 21775 18717 21787 18751
rect 21729 18711 21787 18717
rect 21821 18751 21879 18757
rect 21821 18717 21833 18751
rect 21867 18717 21879 18751
rect 21821 18711 21879 18717
rect 21913 18751 21971 18757
rect 21913 18717 21925 18751
rect 21959 18750 21971 18751
rect 22002 18750 22008 18760
rect 21959 18722 22008 18750
rect 21959 18717 21971 18722
rect 21913 18711 21971 18717
rect 22002 18708 22008 18722
rect 22060 18708 22066 18760
rect 22094 18708 22100 18760
rect 22152 18748 22158 18760
rect 22152 18720 22197 18748
rect 22152 18708 22158 18720
rect 22462 18708 22468 18760
rect 22520 18748 22526 18760
rect 22557 18751 22615 18757
rect 22557 18748 22569 18751
rect 22520 18720 22569 18748
rect 22520 18708 22526 18720
rect 22557 18717 22569 18720
rect 22603 18717 22615 18751
rect 22557 18711 22615 18717
rect 24946 18708 24952 18760
rect 25004 18748 25010 18760
rect 25694 18751 25752 18757
rect 25694 18748 25706 18751
rect 25004 18720 25706 18748
rect 25004 18708 25010 18720
rect 25694 18717 25706 18720
rect 25740 18717 25752 18751
rect 25694 18711 25752 18717
rect 27525 18751 27583 18757
rect 27525 18717 27537 18751
rect 27571 18748 27583 18751
rect 28350 18748 28356 18760
rect 27571 18720 28356 18748
rect 27571 18717 27583 18720
rect 27525 18711 27583 18717
rect 28350 18708 28356 18720
rect 28408 18708 28414 18760
rect 28810 18748 28816 18760
rect 28771 18720 28816 18748
rect 28810 18708 28816 18720
rect 28868 18708 28874 18760
rect 28997 18751 29055 18757
rect 28997 18717 29009 18751
rect 29043 18748 29055 18751
rect 29546 18748 29552 18760
rect 29043 18720 29552 18748
rect 29043 18717 29055 18720
rect 28997 18711 29055 18717
rect 29546 18708 29552 18720
rect 29604 18708 29610 18760
rect 29733 18751 29791 18757
rect 29733 18717 29745 18751
rect 29779 18748 29791 18751
rect 30190 18748 30196 18760
rect 29779 18720 30196 18748
rect 29779 18717 29791 18720
rect 29733 18711 29791 18717
rect 30190 18708 30196 18720
rect 30248 18708 30254 18760
rect 30300 18748 30328 18788
rect 32309 18785 32321 18819
rect 32355 18816 32367 18819
rect 35342 18816 35348 18828
rect 32355 18788 35348 18816
rect 32355 18785 32367 18788
rect 32309 18779 32367 18785
rect 35342 18776 35348 18788
rect 35400 18776 35406 18828
rect 38105 18819 38163 18825
rect 38105 18785 38117 18819
rect 38151 18816 38163 18819
rect 39022 18816 39028 18828
rect 38151 18788 39028 18816
rect 38151 18785 38163 18788
rect 38105 18779 38163 18785
rect 39022 18776 39028 18788
rect 39080 18776 39086 18828
rect 32950 18748 32956 18760
rect 30300 18720 32956 18748
rect 32950 18708 32956 18720
rect 33008 18708 33014 18760
rect 33134 18748 33140 18760
rect 33095 18720 33140 18748
rect 33134 18708 33140 18720
rect 33192 18708 33198 18760
rect 33413 18751 33471 18757
rect 33413 18717 33425 18751
rect 33459 18748 33471 18751
rect 33594 18748 33600 18760
rect 33459 18720 33600 18748
rect 33459 18717 33471 18720
rect 33413 18711 33471 18717
rect 33594 18708 33600 18720
rect 33652 18748 33658 18760
rect 37550 18748 37556 18760
rect 33652 18720 37556 18748
rect 33652 18708 33658 18720
rect 37550 18708 37556 18720
rect 37608 18748 37614 18760
rect 37826 18748 37832 18760
rect 37608 18720 37832 18748
rect 37608 18708 37614 18720
rect 37826 18708 37832 18720
rect 37884 18748 37890 18760
rect 38565 18751 38623 18757
rect 38565 18748 38577 18751
rect 37884 18720 38577 18748
rect 37884 18708 37890 18720
rect 38565 18717 38577 18720
rect 38611 18717 38623 18751
rect 38744 18751 38802 18757
rect 38744 18748 38756 18751
rect 38565 18711 38623 18717
rect 38672 18720 38756 18748
rect 16623 18652 19288 18680
rect 21453 18683 21511 18689
rect 16623 18649 16635 18652
rect 16577 18643 16635 18649
rect 21453 18649 21465 18683
rect 21499 18680 21511 18683
rect 24118 18680 24124 18692
rect 21499 18652 24124 18680
rect 21499 18649 21511 18652
rect 21453 18643 21511 18649
rect 24118 18640 24124 18652
rect 24176 18640 24182 18692
rect 27709 18683 27767 18689
rect 27709 18649 27721 18683
rect 27755 18680 27767 18683
rect 29917 18683 29975 18689
rect 27755 18652 29040 18680
rect 27755 18649 27767 18652
rect 27709 18643 27767 18649
rect 29012 18624 29040 18652
rect 29917 18649 29929 18683
rect 29963 18649 29975 18683
rect 29917 18643 29975 18649
rect 30469 18683 30527 18689
rect 30469 18649 30481 18683
rect 30515 18680 30527 18683
rect 31478 18680 31484 18692
rect 30515 18652 31484 18680
rect 30515 18649 30527 18652
rect 30469 18643 30527 18649
rect 16942 18612 16948 18624
rect 14568 18584 15608 18612
rect 16903 18584 16948 18612
rect 16942 18572 16948 18584
rect 17000 18572 17006 18624
rect 17402 18572 17408 18624
rect 17460 18612 17466 18624
rect 17589 18615 17647 18621
rect 17589 18612 17601 18615
rect 17460 18584 17601 18612
rect 17460 18572 17466 18584
rect 17589 18581 17601 18584
rect 17635 18581 17647 18615
rect 17589 18575 17647 18581
rect 18693 18615 18751 18621
rect 18693 18581 18705 18615
rect 18739 18612 18751 18615
rect 20806 18612 20812 18624
rect 18739 18584 20812 18612
rect 18739 18581 18751 18584
rect 18693 18575 18751 18581
rect 20806 18572 20812 18584
rect 20864 18572 20870 18624
rect 20898 18572 20904 18624
rect 20956 18612 20962 18624
rect 24578 18612 24584 18624
rect 20956 18584 24584 18612
rect 20956 18572 20962 18584
rect 24578 18572 24584 18584
rect 24636 18572 24642 18624
rect 28166 18572 28172 18624
rect 28224 18612 28230 18624
rect 28353 18615 28411 18621
rect 28353 18612 28365 18615
rect 28224 18584 28365 18612
rect 28224 18572 28230 18584
rect 28353 18581 28365 18584
rect 28399 18612 28411 18615
rect 28810 18612 28816 18624
rect 28399 18584 28816 18612
rect 28399 18581 28411 18584
rect 28353 18575 28411 18581
rect 28810 18572 28816 18584
rect 28868 18572 28874 18624
rect 28994 18572 29000 18624
rect 29052 18612 29058 18624
rect 29932 18612 29960 18643
rect 31478 18640 31484 18652
rect 31536 18640 31542 18692
rect 31938 18640 31944 18692
rect 31996 18680 32002 18692
rect 32042 18683 32100 18689
rect 32042 18680 32054 18683
rect 31996 18652 32054 18680
rect 31996 18640 32002 18652
rect 32042 18649 32054 18652
rect 32088 18649 32100 18683
rect 36357 18683 36415 18689
rect 36357 18680 36369 18683
rect 32042 18643 32100 18649
rect 35912 18652 36369 18680
rect 35912 18624 35940 18652
rect 36357 18649 36369 18652
rect 36403 18649 36415 18683
rect 36357 18643 36415 18649
rect 38102 18640 38108 18692
rect 38160 18680 38166 18692
rect 38672 18680 38700 18720
rect 38744 18717 38756 18720
rect 38790 18717 38802 18751
rect 38744 18711 38802 18717
rect 38841 18751 38899 18757
rect 38841 18717 38853 18751
rect 38887 18717 38899 18751
rect 38841 18711 38899 18717
rect 38160 18652 38700 18680
rect 38160 18640 38166 18652
rect 29052 18584 29960 18612
rect 30929 18615 30987 18621
rect 29052 18572 29058 18584
rect 30929 18581 30941 18615
rect 30975 18612 30987 18615
rect 31018 18612 31024 18624
rect 30975 18584 31024 18612
rect 30975 18581 30987 18584
rect 30929 18575 30987 18581
rect 31018 18572 31024 18584
rect 31076 18572 31082 18624
rect 35894 18612 35900 18624
rect 35855 18584 35900 18612
rect 35894 18572 35900 18584
rect 35952 18572 35958 18624
rect 37366 18572 37372 18624
rect 37424 18612 37430 18624
rect 38856 18612 38884 18711
rect 38930 18708 38936 18760
rect 38988 18748 38994 18760
rect 39853 18751 39911 18757
rect 39853 18748 39865 18751
rect 38988 18720 39865 18748
rect 38988 18708 38994 18720
rect 39853 18717 39865 18720
rect 39899 18717 39911 18751
rect 68094 18748 68100 18760
rect 68055 18720 68100 18748
rect 39853 18711 39911 18717
rect 68094 18708 68100 18720
rect 68152 18708 68158 18760
rect 37424 18584 38884 18612
rect 37424 18572 37430 18584
rect 1104 18522 68816 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 68816 18522
rect 1104 18448 68816 18470
rect 8018 18368 8024 18420
rect 8076 18408 8082 18420
rect 8205 18411 8263 18417
rect 8205 18408 8217 18411
rect 8076 18380 8217 18408
rect 8076 18368 8082 18380
rect 8205 18377 8217 18380
rect 8251 18377 8263 18411
rect 11514 18408 11520 18420
rect 11475 18380 11520 18408
rect 8205 18371 8263 18377
rect 11514 18368 11520 18380
rect 11572 18368 11578 18420
rect 14093 18411 14151 18417
rect 14093 18408 14105 18411
rect 11900 18380 14105 18408
rect 2501 18343 2559 18349
rect 2501 18309 2513 18343
rect 2547 18340 2559 18343
rect 3418 18340 3424 18352
rect 2547 18312 2912 18340
rect 2547 18309 2559 18312
rect 2501 18303 2559 18309
rect 1854 18272 1860 18284
rect 1815 18244 1860 18272
rect 1854 18232 1860 18244
rect 1912 18232 1918 18284
rect 2038 18281 2044 18284
rect 2036 18272 2044 18281
rect 1999 18244 2044 18272
rect 2036 18235 2044 18244
rect 2038 18232 2044 18235
rect 2096 18232 2102 18284
rect 2130 18232 2136 18284
rect 2188 18272 2194 18284
rect 2271 18275 2329 18281
rect 2188 18244 2233 18272
rect 2188 18232 2194 18244
rect 2271 18241 2283 18275
rect 2317 18272 2329 18275
rect 2682 18272 2688 18284
rect 2317 18244 2688 18272
rect 2317 18241 2329 18244
rect 2271 18235 2329 18241
rect 2682 18232 2688 18244
rect 2740 18232 2746 18284
rect 2884 18204 2912 18312
rect 2976 18312 3424 18340
rect 2976 18281 3004 18312
rect 3418 18300 3424 18312
rect 3476 18300 3482 18352
rect 8846 18340 8852 18352
rect 8807 18312 8852 18340
rect 8846 18300 8852 18312
rect 8904 18300 8910 18352
rect 9033 18343 9091 18349
rect 9033 18309 9045 18343
rect 9079 18340 9091 18343
rect 11900 18340 11928 18380
rect 14093 18377 14105 18380
rect 14139 18408 14151 18411
rect 16666 18408 16672 18420
rect 14139 18380 16672 18408
rect 14139 18377 14151 18380
rect 14093 18371 14151 18377
rect 16666 18368 16672 18380
rect 16724 18368 16730 18420
rect 20898 18408 20904 18420
rect 18340 18380 20904 18408
rect 13170 18340 13176 18352
rect 9079 18312 11928 18340
rect 11992 18312 13176 18340
rect 9079 18309 9091 18312
rect 9033 18303 9091 18309
rect 2961 18275 3019 18281
rect 2961 18241 2973 18275
rect 3007 18241 3019 18275
rect 3217 18275 3275 18281
rect 3217 18272 3229 18275
rect 2961 18235 3019 18241
rect 3068 18244 3229 18272
rect 3068 18204 3096 18244
rect 3217 18241 3229 18244
rect 3263 18241 3275 18275
rect 3217 18235 3275 18241
rect 6914 18232 6920 18284
rect 6972 18272 6978 18284
rect 7478 18275 7536 18281
rect 7478 18272 7490 18275
rect 6972 18244 7490 18272
rect 6972 18232 6978 18244
rect 7478 18241 7490 18244
rect 7524 18241 7536 18275
rect 7478 18235 7536 18241
rect 7745 18275 7803 18281
rect 7745 18241 7757 18275
rect 7791 18272 7803 18275
rect 8018 18272 8024 18284
rect 7791 18244 8024 18272
rect 7791 18241 7803 18244
rect 7745 18235 7803 18241
rect 8018 18232 8024 18244
rect 8076 18272 8082 18284
rect 8294 18272 8300 18284
rect 8076 18244 8300 18272
rect 8076 18232 8082 18244
rect 8294 18232 8300 18244
rect 8352 18232 8358 18284
rect 8389 18275 8447 18281
rect 8389 18241 8401 18275
rect 8435 18272 8447 18275
rect 8864 18272 8892 18300
rect 8435 18244 8892 18272
rect 8435 18241 8447 18244
rect 8389 18235 8447 18241
rect 9674 18232 9680 18284
rect 9732 18272 9738 18284
rect 11790 18272 11796 18284
rect 9732 18244 9777 18272
rect 11751 18244 11796 18272
rect 9732 18232 9738 18244
rect 11790 18232 11796 18244
rect 11848 18232 11854 18284
rect 11992 18281 12020 18312
rect 13170 18300 13176 18312
rect 13228 18300 13234 18352
rect 15838 18340 15844 18352
rect 15799 18312 15844 18340
rect 15838 18300 15844 18312
rect 15896 18300 15902 18352
rect 16114 18300 16120 18352
rect 16172 18340 16178 18352
rect 16172 18312 16620 18340
rect 16172 18300 16178 18312
rect 11885 18275 11943 18281
rect 11885 18241 11897 18275
rect 11931 18241 11943 18275
rect 11885 18235 11943 18241
rect 11977 18275 12035 18281
rect 11977 18241 11989 18275
rect 12023 18241 12035 18275
rect 12158 18272 12164 18284
rect 12119 18244 12164 18272
rect 11977 18235 12035 18241
rect 2884 18176 3096 18204
rect 9953 18207 10011 18213
rect 9953 18173 9965 18207
rect 9999 18204 10011 18207
rect 10594 18204 10600 18216
rect 9999 18176 10600 18204
rect 9999 18173 10011 18176
rect 9953 18167 10011 18173
rect 10594 18164 10600 18176
rect 10652 18204 10658 18216
rect 11900 18204 11928 18235
rect 12158 18232 12164 18244
rect 12216 18232 12222 18284
rect 12250 18232 12256 18284
rect 12308 18272 12314 18284
rect 12969 18275 13027 18281
rect 12969 18272 12981 18275
rect 12308 18244 12981 18272
rect 12308 18232 12314 18244
rect 12969 18241 12981 18244
rect 13015 18241 13027 18275
rect 12969 18235 13027 18241
rect 15286 18232 15292 18284
rect 15344 18272 15350 18284
rect 16025 18275 16083 18281
rect 16025 18272 16037 18275
rect 15344 18244 16037 18272
rect 15344 18232 15350 18244
rect 16025 18241 16037 18244
rect 16071 18272 16083 18275
rect 16482 18272 16488 18284
rect 16071 18244 16488 18272
rect 16071 18241 16083 18244
rect 16025 18235 16083 18241
rect 16482 18232 16488 18244
rect 16540 18232 16546 18284
rect 16592 18272 16620 18312
rect 16942 18300 16948 18352
rect 17000 18340 17006 18352
rect 17000 18312 17724 18340
rect 17000 18300 17006 18312
rect 17126 18272 17132 18284
rect 16592 18244 17132 18272
rect 17126 18232 17132 18244
rect 17184 18281 17190 18284
rect 17184 18275 17233 18281
rect 17184 18241 17187 18275
rect 17221 18241 17233 18275
rect 17310 18272 17316 18284
rect 17271 18244 17316 18272
rect 17184 18235 17233 18241
rect 17184 18232 17190 18235
rect 17310 18232 17316 18244
rect 17368 18232 17374 18284
rect 17696 18281 17724 18312
rect 17405 18275 17463 18281
rect 17405 18241 17417 18275
rect 17451 18241 17463 18275
rect 17405 18235 17463 18241
rect 17588 18275 17646 18281
rect 17588 18241 17600 18275
rect 17634 18241 17646 18275
rect 17588 18235 17646 18241
rect 17681 18275 17739 18281
rect 17681 18241 17693 18275
rect 17727 18241 17739 18275
rect 17681 18235 17739 18241
rect 10652 18176 11928 18204
rect 10652 18164 10658 18176
rect 4341 18071 4399 18077
rect 4341 18037 4353 18071
rect 4387 18068 4399 18071
rect 4614 18068 4620 18080
rect 4387 18040 4620 18068
rect 4387 18037 4399 18040
rect 4341 18031 4399 18037
rect 4614 18028 4620 18040
rect 4672 18028 4678 18080
rect 6362 18068 6368 18080
rect 6323 18040 6368 18068
rect 6362 18028 6368 18040
rect 6420 18028 6426 18080
rect 9217 18071 9275 18077
rect 9217 18037 9229 18071
rect 9263 18068 9275 18071
rect 9490 18068 9496 18080
rect 9263 18040 9496 18068
rect 9263 18037 9275 18040
rect 9217 18031 9275 18037
rect 9490 18028 9496 18040
rect 9548 18028 9554 18080
rect 11900 18068 11928 18176
rect 12434 18164 12440 18216
rect 12492 18204 12498 18216
rect 12713 18207 12771 18213
rect 12713 18204 12725 18207
rect 12492 18176 12725 18204
rect 12492 18164 12498 18176
rect 12713 18173 12725 18176
rect 12759 18173 12771 18207
rect 12713 18167 12771 18173
rect 16390 18164 16396 18216
rect 16448 18204 16454 18216
rect 17420 18204 17448 18235
rect 16448 18176 17448 18204
rect 17604 18204 17632 18235
rect 18340 18204 18368 18380
rect 20898 18368 20904 18380
rect 20956 18368 20962 18420
rect 21910 18368 21916 18420
rect 21968 18408 21974 18420
rect 22189 18411 22247 18417
rect 22189 18408 22201 18411
rect 21968 18380 22201 18408
rect 21968 18368 21974 18380
rect 22189 18377 22201 18380
rect 22235 18377 22247 18411
rect 22189 18371 22247 18377
rect 22278 18368 22284 18420
rect 22336 18408 22342 18420
rect 27709 18411 27767 18417
rect 27709 18408 27721 18411
rect 22336 18380 27721 18408
rect 22336 18368 22342 18380
rect 27709 18377 27721 18380
rect 27755 18408 27767 18411
rect 28718 18408 28724 18420
rect 27755 18380 28724 18408
rect 27755 18377 27767 18380
rect 27709 18371 27767 18377
rect 28718 18368 28724 18380
rect 28776 18368 28782 18420
rect 28810 18368 28816 18420
rect 28868 18408 28874 18420
rect 38102 18408 38108 18420
rect 28868 18380 29868 18408
rect 38063 18380 38108 18408
rect 28868 18368 28874 18380
rect 20257 18343 20315 18349
rect 20257 18309 20269 18343
rect 20303 18340 20315 18343
rect 21082 18340 21088 18352
rect 20303 18312 21088 18340
rect 20303 18309 20315 18312
rect 20257 18303 20315 18309
rect 21082 18300 21088 18312
rect 21140 18300 21146 18352
rect 21174 18300 21180 18352
rect 21232 18340 21238 18352
rect 22005 18343 22063 18349
rect 22005 18340 22017 18343
rect 21232 18312 22017 18340
rect 21232 18300 21238 18312
rect 22005 18309 22017 18312
rect 22051 18309 22063 18343
rect 22005 18303 22063 18309
rect 18690 18272 18696 18284
rect 18651 18244 18696 18272
rect 18690 18232 18696 18244
rect 18748 18232 18754 18284
rect 20070 18232 20076 18284
rect 20128 18281 20134 18284
rect 20128 18275 20177 18281
rect 20128 18241 20131 18275
rect 20165 18241 20177 18275
rect 20128 18235 20177 18241
rect 20349 18275 20407 18281
rect 20349 18241 20361 18275
rect 20395 18241 20407 18275
rect 20530 18272 20536 18284
rect 20491 18244 20536 18272
rect 20349 18235 20407 18241
rect 20128 18232 20134 18235
rect 17604 18176 18368 18204
rect 18417 18207 18475 18213
rect 16448 18164 16454 18176
rect 18417 18173 18429 18207
rect 18463 18173 18475 18207
rect 18417 18167 18475 18173
rect 16758 18096 16764 18148
rect 16816 18136 16822 18148
rect 18432 18136 18460 18167
rect 16816 18108 18460 18136
rect 16816 18096 16822 18108
rect 19426 18096 19432 18148
rect 19484 18136 19490 18148
rect 20364 18136 20392 18235
rect 20530 18232 20536 18244
rect 20588 18232 20594 18284
rect 20622 18232 20628 18284
rect 20680 18272 20686 18284
rect 21266 18272 21272 18284
rect 20680 18244 20725 18272
rect 21227 18244 21272 18272
rect 20680 18232 20686 18244
rect 21266 18232 21272 18244
rect 21324 18232 21330 18284
rect 21821 18275 21879 18281
rect 21821 18241 21833 18275
rect 21867 18241 21879 18275
rect 21821 18235 21879 18241
rect 21836 18204 21864 18235
rect 21100 18176 21864 18204
rect 20714 18136 20720 18148
rect 19484 18108 20116 18136
rect 20364 18108 20720 18136
rect 19484 18096 19490 18108
rect 12710 18068 12716 18080
rect 11900 18040 12716 18068
rect 12710 18028 12716 18040
rect 12768 18028 12774 18080
rect 17037 18071 17095 18077
rect 17037 18037 17049 18071
rect 17083 18068 17095 18071
rect 17126 18068 17132 18080
rect 17083 18040 17132 18068
rect 17083 18037 17095 18040
rect 17037 18031 17095 18037
rect 17126 18028 17132 18040
rect 17184 18028 17190 18080
rect 19978 18068 19984 18080
rect 19939 18040 19984 18068
rect 19978 18028 19984 18040
rect 20036 18028 20042 18080
rect 20088 18068 20116 18108
rect 20714 18096 20720 18108
rect 20772 18096 20778 18148
rect 21100 18077 21128 18176
rect 21085 18071 21143 18077
rect 21085 18068 21097 18071
rect 20088 18040 21097 18068
rect 21085 18037 21097 18040
rect 21131 18037 21143 18071
rect 22020 18068 22048 18303
rect 24118 18300 24124 18352
rect 24176 18349 24182 18352
rect 24176 18340 24188 18349
rect 24176 18312 24221 18340
rect 24176 18303 24188 18312
rect 24176 18300 24182 18303
rect 28442 18300 28448 18352
rect 28500 18340 28506 18352
rect 28500 18312 29684 18340
rect 28500 18300 28506 18312
rect 26326 18272 26332 18284
rect 26287 18244 26332 18272
rect 26326 18232 26332 18244
rect 26384 18272 26390 18284
rect 29656 18281 29684 18312
rect 29840 18281 29868 18380
rect 38102 18368 38108 18380
rect 38160 18368 38166 18420
rect 30282 18300 30288 18352
rect 30340 18340 30346 18352
rect 30837 18343 30895 18349
rect 30837 18340 30849 18343
rect 30340 18312 30849 18340
rect 30340 18300 30346 18312
rect 30837 18309 30849 18312
rect 30883 18340 30895 18343
rect 30883 18312 31754 18340
rect 30883 18309 30895 18312
rect 30837 18303 30895 18309
rect 28997 18275 29055 18281
rect 28997 18272 29009 18275
rect 26384 18270 28304 18272
rect 28460 18270 29009 18272
rect 26384 18244 29009 18270
rect 26384 18232 26390 18244
rect 28276 18242 28488 18244
rect 28997 18241 29009 18244
rect 29043 18241 29055 18275
rect 28997 18235 29055 18241
rect 29641 18275 29699 18281
rect 29641 18241 29653 18275
rect 29687 18241 29699 18275
rect 29641 18235 29699 18241
rect 29825 18275 29883 18281
rect 29825 18241 29837 18275
rect 29871 18241 29883 18275
rect 31018 18272 31024 18284
rect 30979 18244 31024 18272
rect 29825 18235 29883 18241
rect 31018 18232 31024 18244
rect 31076 18232 31082 18284
rect 31726 18272 31754 18312
rect 33318 18300 33324 18352
rect 33376 18340 33382 18352
rect 34241 18343 34299 18349
rect 34241 18340 34253 18343
rect 33376 18312 34253 18340
rect 33376 18300 33382 18312
rect 34241 18309 34253 18312
rect 34287 18309 34299 18343
rect 34241 18303 34299 18309
rect 37458 18300 37464 18352
rect 37516 18340 37522 18352
rect 37737 18343 37795 18349
rect 37737 18340 37749 18343
rect 37516 18312 37749 18340
rect 37516 18300 37522 18312
rect 37737 18309 37749 18312
rect 37783 18309 37795 18343
rect 37737 18303 37795 18309
rect 32125 18275 32183 18281
rect 32125 18272 32137 18275
rect 31726 18244 32137 18272
rect 32125 18241 32137 18244
rect 32171 18241 32183 18275
rect 32125 18235 32183 18241
rect 34425 18275 34483 18281
rect 34425 18241 34437 18275
rect 34471 18272 34483 18275
rect 34698 18272 34704 18284
rect 34471 18244 34704 18272
rect 34471 18241 34483 18244
rect 34425 18235 34483 18241
rect 24394 18204 24400 18216
rect 24355 18176 24400 18204
rect 24394 18164 24400 18176
rect 24452 18164 24458 18216
rect 25222 18164 25228 18216
rect 25280 18204 25286 18216
rect 26053 18207 26111 18213
rect 26053 18204 26065 18207
rect 25280 18176 26065 18204
rect 25280 18164 25286 18176
rect 26053 18173 26065 18176
rect 26099 18173 26111 18207
rect 26053 18167 26111 18173
rect 23017 18139 23075 18145
rect 23017 18105 23029 18139
rect 23063 18105 23075 18139
rect 26068 18136 26096 18167
rect 27614 18164 27620 18216
rect 27672 18204 27678 18216
rect 28166 18204 28172 18216
rect 27672 18176 28172 18204
rect 27672 18164 27678 18176
rect 28166 18164 28172 18176
rect 28224 18204 28230 18216
rect 28261 18207 28319 18213
rect 28261 18204 28273 18207
rect 28224 18176 28273 18204
rect 28224 18164 28230 18176
rect 28261 18173 28273 18176
rect 28307 18173 28319 18207
rect 28261 18167 28319 18173
rect 28718 18164 28724 18216
rect 28776 18204 28782 18216
rect 28813 18207 28871 18213
rect 28813 18204 28825 18207
rect 28776 18176 28825 18204
rect 28776 18164 28782 18176
rect 28813 18173 28825 18176
rect 28859 18173 28871 18207
rect 29730 18204 29736 18216
rect 29643 18176 29736 18204
rect 28813 18167 28871 18173
rect 28442 18136 28448 18148
rect 26068 18108 28448 18136
rect 23017 18099 23075 18105
rect 23032 18068 23060 18099
rect 28442 18096 28448 18108
rect 28500 18096 28506 18148
rect 22020 18040 23060 18068
rect 28828 18068 28856 18167
rect 29730 18164 29736 18176
rect 29788 18204 29794 18216
rect 31110 18204 31116 18216
rect 29788 18176 31116 18204
rect 29788 18164 29794 18176
rect 31110 18164 31116 18176
rect 31168 18204 31174 18216
rect 32769 18207 32827 18213
rect 32769 18204 32781 18207
rect 31168 18176 32781 18204
rect 31168 18164 31174 18176
rect 32769 18173 32781 18176
rect 32815 18173 32827 18207
rect 32769 18167 32827 18173
rect 33045 18207 33103 18213
rect 33045 18173 33057 18207
rect 33091 18204 33103 18207
rect 33502 18204 33508 18216
rect 33091 18176 33508 18204
rect 33091 18173 33103 18176
rect 33045 18167 33103 18173
rect 33502 18164 33508 18176
rect 33560 18164 33566 18216
rect 29178 18096 29184 18148
rect 29236 18136 29242 18148
rect 30282 18136 30288 18148
rect 29236 18108 30288 18136
rect 29236 18096 29242 18108
rect 30282 18096 30288 18108
rect 30340 18096 30346 18148
rect 31386 18136 31392 18148
rect 30392 18108 31392 18136
rect 30392 18077 30420 18108
rect 31386 18096 31392 18108
rect 31444 18096 31450 18148
rect 32309 18139 32367 18145
rect 32309 18105 32321 18139
rect 32355 18136 32367 18139
rect 34440 18136 34468 18235
rect 34698 18232 34704 18244
rect 34756 18232 34762 18284
rect 35342 18272 35348 18284
rect 35303 18244 35348 18272
rect 35342 18232 35348 18244
rect 35400 18232 35406 18284
rect 35434 18232 35440 18284
rect 35492 18272 35498 18284
rect 35601 18275 35659 18281
rect 35601 18272 35613 18275
rect 35492 18244 35613 18272
rect 35492 18232 35498 18244
rect 35601 18241 35613 18244
rect 35647 18241 35659 18275
rect 37918 18272 37924 18284
rect 37879 18244 37924 18272
rect 35601 18235 35659 18241
rect 37918 18232 37924 18244
rect 37976 18232 37982 18284
rect 38654 18232 38660 18284
rect 38712 18272 38718 18284
rect 39281 18275 39339 18281
rect 39281 18272 39293 18275
rect 38712 18244 39293 18272
rect 38712 18232 38718 18244
rect 39281 18241 39293 18244
rect 39327 18241 39339 18275
rect 39281 18235 39339 18241
rect 39022 18204 39028 18216
rect 38983 18176 39028 18204
rect 39022 18164 39028 18176
rect 39080 18164 39086 18216
rect 32355 18108 34468 18136
rect 32355 18105 32367 18108
rect 32309 18099 32367 18105
rect 30377 18071 30435 18077
rect 30377 18068 30389 18071
rect 28828 18040 30389 18068
rect 21085 18031 21143 18037
rect 30377 18037 30389 18040
rect 30423 18037 30435 18071
rect 30377 18031 30435 18037
rect 31018 18028 31024 18080
rect 31076 18068 31082 18080
rect 31205 18071 31263 18077
rect 31205 18068 31217 18071
rect 31076 18040 31217 18068
rect 31076 18028 31082 18040
rect 31205 18037 31217 18040
rect 31251 18037 31263 18071
rect 31205 18031 31263 18037
rect 33410 18028 33416 18080
rect 33468 18068 33474 18080
rect 34057 18071 34115 18077
rect 34057 18068 34069 18071
rect 33468 18040 34069 18068
rect 33468 18028 33474 18040
rect 34057 18037 34069 18040
rect 34103 18037 34115 18071
rect 36722 18068 36728 18080
rect 36683 18040 36728 18068
rect 34057 18031 34115 18037
rect 36722 18028 36728 18040
rect 36780 18028 36786 18080
rect 40402 18068 40408 18080
rect 40363 18040 40408 18068
rect 40402 18028 40408 18040
rect 40460 18028 40466 18080
rect 1104 17978 68816 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 65654 17978
rect 65706 17926 65718 17978
rect 65770 17926 65782 17978
rect 65834 17926 65846 17978
rect 65898 17926 65910 17978
rect 65962 17926 68816 17978
rect 1104 17904 68816 17926
rect 2682 17864 2688 17876
rect 2643 17836 2688 17864
rect 2682 17824 2688 17836
rect 2740 17824 2746 17876
rect 10045 17867 10103 17873
rect 10045 17833 10057 17867
rect 10091 17864 10103 17867
rect 12250 17864 12256 17876
rect 10091 17836 12256 17864
rect 10091 17833 10103 17836
rect 10045 17827 10103 17833
rect 12250 17824 12256 17836
rect 12308 17824 12314 17876
rect 20530 17824 20536 17876
rect 20588 17864 20594 17876
rect 22278 17864 22284 17876
rect 20588 17836 22284 17864
rect 20588 17824 20594 17836
rect 22278 17824 22284 17836
rect 22336 17824 22342 17876
rect 24762 17864 24768 17876
rect 24723 17836 24768 17864
rect 24762 17824 24768 17836
rect 24820 17824 24826 17876
rect 26970 17824 26976 17876
rect 27028 17864 27034 17876
rect 27028 17836 27936 17864
rect 27028 17824 27034 17836
rect 20898 17796 20904 17808
rect 9646 17768 9996 17796
rect 2038 17688 2044 17740
rect 2096 17728 2102 17740
rect 4157 17731 4215 17737
rect 4157 17728 4169 17731
rect 2096 17700 4169 17728
rect 2096 17688 2102 17700
rect 4157 17697 4169 17700
rect 4203 17697 4215 17731
rect 4157 17691 4215 17697
rect 7009 17731 7067 17737
rect 7009 17697 7021 17731
rect 7055 17728 7067 17731
rect 7098 17728 7104 17740
rect 7055 17700 7104 17728
rect 7055 17697 7067 17700
rect 7009 17691 7067 17697
rect 7098 17688 7104 17700
rect 7156 17688 7162 17740
rect 7374 17688 7380 17740
rect 7432 17728 7438 17740
rect 8202 17728 8208 17740
rect 7432 17700 8208 17728
rect 7432 17688 7438 17700
rect 8202 17688 8208 17700
rect 8260 17728 8266 17740
rect 9646 17728 9674 17768
rect 8260 17700 9674 17728
rect 8260 17688 8266 17700
rect 4341 17663 4399 17669
rect 4341 17629 4353 17663
rect 4387 17660 4399 17663
rect 4614 17660 4620 17672
rect 4387 17632 4620 17660
rect 4387 17629 4399 17632
rect 4341 17623 4399 17629
rect 4614 17620 4620 17632
rect 4672 17660 4678 17672
rect 5350 17660 5356 17672
rect 4672 17632 5356 17660
rect 4672 17620 4678 17632
rect 5350 17620 5356 17632
rect 5408 17620 5414 17672
rect 7285 17663 7343 17669
rect 7285 17629 7297 17663
rect 7331 17629 7343 17663
rect 9398 17660 9404 17672
rect 9359 17632 9404 17660
rect 7285 17623 7343 17629
rect 4525 17595 4583 17601
rect 4525 17561 4537 17595
rect 4571 17592 4583 17595
rect 4798 17592 4804 17604
rect 4571 17564 4804 17592
rect 4571 17561 4583 17564
rect 4525 17555 4583 17561
rect 4798 17552 4804 17564
rect 4856 17552 4862 17604
rect 7098 17552 7104 17604
rect 7156 17592 7162 17604
rect 7300 17592 7328 17623
rect 9398 17620 9404 17632
rect 9456 17620 9462 17672
rect 9490 17620 9496 17672
rect 9548 17660 9554 17672
rect 9585 17660 9643 17666
rect 9548 17632 9597 17660
rect 9548 17620 9554 17632
rect 9585 17626 9597 17632
rect 9631 17626 9643 17660
rect 9585 17620 9643 17626
rect 9674 17620 9680 17672
rect 9732 17660 9738 17672
rect 9815 17663 9873 17669
rect 9732 17632 9777 17660
rect 9732 17620 9738 17632
rect 9815 17629 9827 17663
rect 9861 17660 9873 17663
rect 9968 17660 9996 17768
rect 19536 17768 20904 17796
rect 12434 17688 12440 17740
rect 12492 17728 12498 17740
rect 14553 17731 14611 17737
rect 14553 17728 14565 17731
rect 12492 17700 14565 17728
rect 12492 17688 12498 17700
rect 14553 17697 14565 17700
rect 14599 17697 14611 17731
rect 17402 17728 17408 17740
rect 14553 17691 14611 17697
rect 16960 17700 17408 17728
rect 9861 17632 9996 17660
rect 12989 17663 13047 17669
rect 9861 17629 9873 17632
rect 9815 17623 9873 17629
rect 12989 17629 13001 17663
rect 13035 17660 13047 17663
rect 16022 17660 16028 17672
rect 13035 17632 16028 17660
rect 13035 17629 13047 17632
rect 12989 17623 13047 17629
rect 16022 17620 16028 17632
rect 16080 17620 16086 17672
rect 16850 17660 16856 17672
rect 16811 17632 16856 17660
rect 16850 17620 16856 17632
rect 16908 17620 16914 17672
rect 16960 17669 16988 17700
rect 17402 17688 17408 17700
rect 17460 17688 17466 17740
rect 16942 17663 17000 17669
rect 16942 17629 16954 17663
rect 16988 17629 17000 17663
rect 16942 17623 17000 17629
rect 17034 17620 17040 17672
rect 17092 17660 17098 17672
rect 17221 17663 17279 17669
rect 17092 17632 17137 17660
rect 17092 17620 17098 17632
rect 17221 17629 17233 17663
rect 17267 17660 17279 17663
rect 17310 17660 17316 17672
rect 17267 17632 17316 17660
rect 17267 17629 17279 17632
rect 17221 17623 17279 17629
rect 17310 17620 17316 17632
rect 17368 17620 17374 17672
rect 18138 17660 18144 17672
rect 18099 17632 18144 17660
rect 18138 17620 18144 17632
rect 18196 17620 18202 17672
rect 18322 17660 18328 17672
rect 18283 17632 18328 17660
rect 18322 17620 18328 17632
rect 18380 17620 18386 17672
rect 18509 17663 18567 17669
rect 18509 17629 18521 17663
rect 18555 17660 18567 17663
rect 18690 17660 18696 17672
rect 18555 17632 18696 17660
rect 18555 17629 18567 17632
rect 18509 17623 18567 17629
rect 18690 17620 18696 17632
rect 18748 17620 18754 17672
rect 19536 17669 19564 17768
rect 20898 17756 20904 17768
rect 20956 17756 20962 17808
rect 24302 17728 24308 17740
rect 20456 17700 24308 17728
rect 19521 17663 19579 17669
rect 19521 17629 19533 17663
rect 19567 17629 19579 17663
rect 19521 17623 19579 17629
rect 20070 17620 20076 17672
rect 20128 17660 20134 17672
rect 20456 17669 20484 17700
rect 24302 17688 24308 17700
rect 24360 17688 24366 17740
rect 27908 17737 27936 17836
rect 27982 17824 27988 17876
rect 28040 17864 28046 17876
rect 33870 17864 33876 17876
rect 28040 17836 33640 17864
rect 33831 17836 33876 17864
rect 28040 17824 28046 17836
rect 27893 17731 27951 17737
rect 27893 17697 27905 17731
rect 27939 17697 27951 17731
rect 27893 17691 27951 17697
rect 29641 17731 29699 17737
rect 29641 17697 29653 17731
rect 29687 17728 29699 17731
rect 29730 17728 29736 17740
rect 29687 17700 29736 17728
rect 29687 17697 29699 17700
rect 29641 17691 29699 17697
rect 29730 17688 29736 17700
rect 29788 17688 29794 17740
rect 30929 17731 30987 17737
rect 30929 17697 30941 17731
rect 30975 17728 30987 17731
rect 31754 17728 31760 17740
rect 30975 17700 31760 17728
rect 30975 17697 30987 17700
rect 30929 17691 30987 17697
rect 31754 17688 31760 17700
rect 31812 17688 31818 17740
rect 32769 17731 32827 17737
rect 32769 17697 32781 17731
rect 32815 17728 32827 17731
rect 33134 17728 33140 17740
rect 32815 17700 33140 17728
rect 32815 17697 32827 17700
rect 32769 17691 32827 17697
rect 33134 17688 33140 17700
rect 33192 17688 33198 17740
rect 33612 17728 33640 17836
rect 33870 17824 33876 17836
rect 33928 17824 33934 17876
rect 35345 17867 35403 17873
rect 35345 17833 35357 17867
rect 35391 17864 35403 17867
rect 35434 17864 35440 17876
rect 35391 17836 35440 17864
rect 35391 17833 35403 17836
rect 35345 17827 35403 17833
rect 35434 17824 35440 17836
rect 35492 17824 35498 17876
rect 37274 17864 37280 17876
rect 37235 17836 37280 17864
rect 37274 17824 37280 17836
rect 37332 17864 37338 17876
rect 38286 17864 38292 17876
rect 37332 17836 38292 17864
rect 37332 17824 37338 17836
rect 33778 17756 33784 17808
rect 33836 17796 33842 17808
rect 33836 17768 35940 17796
rect 33836 17756 33842 17768
rect 34606 17728 34612 17740
rect 33612 17700 34612 17728
rect 34606 17688 34612 17700
rect 34664 17688 34670 17740
rect 35912 17728 35940 17768
rect 37366 17756 37372 17808
rect 37424 17796 37430 17808
rect 37424 17768 38151 17796
rect 37424 17756 37430 17768
rect 35912 17700 36032 17728
rect 20303 17663 20361 17669
rect 20303 17660 20315 17663
rect 20128 17632 20315 17660
rect 20128 17620 20134 17632
rect 20303 17629 20315 17632
rect 20349 17629 20361 17663
rect 20303 17623 20361 17629
rect 20441 17663 20499 17669
rect 20441 17629 20453 17663
rect 20487 17629 20499 17663
rect 20441 17623 20499 17629
rect 20716 17663 20774 17669
rect 20716 17629 20728 17663
rect 20762 17629 20774 17663
rect 20716 17623 20774 17629
rect 7156 17564 7328 17592
rect 7156 17552 7162 17564
rect 7926 17552 7932 17604
rect 7984 17592 7990 17604
rect 8294 17592 8300 17604
rect 7984 17564 8300 17592
rect 7984 17552 7990 17564
rect 8294 17552 8300 17564
rect 8352 17552 8358 17604
rect 12618 17552 12624 17604
rect 12676 17592 12682 17604
rect 12805 17595 12863 17601
rect 12805 17592 12817 17595
rect 12676 17564 12817 17592
rect 12676 17552 12682 17564
rect 12805 17561 12817 17564
rect 12851 17561 12863 17595
rect 12805 17555 12863 17561
rect 14820 17595 14878 17601
rect 14820 17561 14832 17595
rect 14866 17592 14878 17595
rect 16577 17595 16635 17601
rect 16577 17592 16589 17595
rect 14866 17564 16589 17592
rect 14866 17561 14878 17564
rect 14820 17555 14878 17561
rect 16577 17561 16589 17564
rect 16623 17561 16635 17595
rect 16577 17555 16635 17561
rect 18417 17595 18475 17601
rect 18417 17561 18429 17595
rect 18463 17561 18475 17595
rect 18417 17555 18475 17561
rect 19337 17595 19395 17601
rect 19337 17561 19349 17595
rect 19383 17592 19395 17595
rect 19426 17592 19432 17604
rect 19383 17564 19432 17592
rect 19383 17561 19395 17564
rect 19337 17555 19395 17561
rect 6181 17527 6239 17533
rect 6181 17493 6193 17527
rect 6227 17524 6239 17527
rect 6638 17524 6644 17536
rect 6227 17496 6644 17524
rect 6227 17493 6239 17496
rect 6181 17487 6239 17493
rect 6638 17484 6644 17496
rect 6696 17484 6702 17536
rect 8110 17484 8116 17536
rect 8168 17524 8174 17536
rect 11333 17527 11391 17533
rect 11333 17524 11345 17527
rect 8168 17496 11345 17524
rect 8168 17484 8174 17496
rect 11333 17493 11345 17496
rect 11379 17524 11391 17527
rect 11790 17524 11796 17536
rect 11379 17496 11796 17524
rect 11379 17493 11391 17496
rect 11333 17487 11391 17493
rect 11790 17484 11796 17496
rect 11848 17484 11854 17536
rect 13173 17527 13231 17533
rect 13173 17493 13185 17527
rect 13219 17524 13231 17527
rect 13538 17524 13544 17536
rect 13219 17496 13544 17524
rect 13219 17493 13231 17496
rect 13173 17487 13231 17493
rect 13538 17484 13544 17496
rect 13596 17484 13602 17536
rect 15930 17524 15936 17536
rect 15891 17496 15936 17524
rect 15930 17484 15936 17496
rect 15988 17484 15994 17536
rect 16022 17484 16028 17536
rect 16080 17524 16086 17536
rect 18432 17524 18460 17555
rect 19426 17552 19432 17564
rect 19484 17552 19490 17604
rect 19705 17595 19763 17601
rect 19705 17561 19717 17595
rect 19751 17592 19763 17595
rect 20533 17595 20591 17601
rect 19751 17564 20484 17592
rect 19751 17561 19763 17564
rect 19705 17555 19763 17561
rect 18690 17524 18696 17536
rect 16080 17496 18460 17524
rect 18651 17496 18696 17524
rect 16080 17484 16086 17496
rect 18690 17484 18696 17496
rect 18748 17484 18754 17536
rect 18966 17484 18972 17536
rect 19024 17524 19030 17536
rect 20165 17527 20223 17533
rect 20165 17524 20177 17527
rect 19024 17496 20177 17524
rect 19024 17484 19030 17496
rect 20165 17493 20177 17496
rect 20211 17493 20223 17527
rect 20456 17524 20484 17564
rect 20533 17561 20545 17595
rect 20579 17592 20591 17595
rect 20622 17592 20628 17604
rect 20579 17564 20628 17592
rect 20579 17561 20591 17564
rect 20533 17555 20591 17561
rect 20622 17552 20628 17564
rect 20680 17552 20686 17604
rect 20732 17592 20760 17623
rect 20806 17620 20812 17672
rect 20864 17660 20870 17672
rect 24578 17660 24584 17672
rect 20864 17632 20909 17660
rect 24539 17632 24584 17660
rect 20864 17620 20870 17632
rect 24578 17620 24584 17632
rect 24636 17620 24642 17672
rect 25130 17620 25136 17672
rect 25188 17660 25194 17672
rect 28997 17663 29055 17669
rect 25188 17632 28856 17660
rect 25188 17620 25194 17632
rect 21174 17592 21180 17604
rect 20732 17564 21180 17592
rect 21174 17552 21180 17564
rect 21232 17552 21238 17604
rect 21358 17592 21364 17604
rect 21319 17564 21364 17592
rect 21358 17552 21364 17564
rect 21416 17592 21422 17604
rect 21913 17595 21971 17601
rect 21913 17592 21925 17595
rect 21416 17564 21925 17592
rect 21416 17552 21422 17564
rect 21913 17561 21925 17564
rect 21959 17561 21971 17595
rect 21913 17555 21971 17561
rect 24397 17595 24455 17601
rect 24397 17561 24409 17595
rect 24443 17592 24455 17595
rect 24486 17592 24492 17604
rect 24443 17564 24492 17592
rect 24443 17561 24455 17564
rect 24397 17555 24455 17561
rect 24486 17552 24492 17564
rect 24544 17552 24550 17604
rect 24670 17552 24676 17604
rect 24728 17592 24734 17604
rect 25317 17595 25375 17601
rect 25317 17592 25329 17595
rect 24728 17564 25329 17592
rect 24728 17552 24734 17564
rect 25317 17561 25329 17564
rect 25363 17592 25375 17595
rect 25866 17592 25872 17604
rect 25363 17564 25872 17592
rect 25363 17561 25375 17564
rect 25317 17555 25375 17561
rect 25866 17552 25872 17564
rect 25924 17552 25930 17604
rect 26053 17595 26111 17601
rect 26053 17561 26065 17595
rect 26099 17592 26111 17595
rect 27062 17592 27068 17604
rect 26099 17564 27068 17592
rect 26099 17561 26111 17564
rect 26053 17555 26111 17561
rect 27062 17552 27068 17564
rect 27120 17592 27126 17604
rect 27246 17592 27252 17604
rect 27120 17564 27252 17592
rect 27120 17552 27126 17564
rect 27246 17552 27252 17564
rect 27304 17552 27310 17604
rect 27338 17552 27344 17604
rect 27396 17592 27402 17604
rect 27626 17595 27684 17601
rect 27626 17592 27638 17595
rect 27396 17564 27638 17592
rect 27396 17552 27402 17564
rect 27626 17561 27638 17564
rect 27672 17561 27684 17595
rect 27626 17555 27684 17561
rect 21266 17524 21272 17536
rect 20456 17496 21272 17524
rect 20165 17487 20223 17493
rect 21266 17484 21272 17496
rect 21324 17484 21330 17536
rect 23198 17524 23204 17536
rect 23159 17496 23204 17524
rect 23198 17484 23204 17496
rect 23256 17484 23262 17536
rect 26510 17524 26516 17536
rect 26471 17496 26516 17524
rect 26510 17484 26516 17496
rect 26568 17484 26574 17536
rect 26602 17484 26608 17536
rect 26660 17524 26666 17536
rect 27982 17524 27988 17536
rect 26660 17496 27988 17524
rect 26660 17484 26666 17496
rect 27982 17484 27988 17496
rect 28040 17484 28046 17536
rect 28828 17533 28856 17632
rect 28997 17629 29009 17663
rect 29043 17660 29055 17663
rect 29178 17660 29184 17672
rect 29043 17632 29184 17660
rect 29043 17629 29055 17632
rect 28997 17623 29055 17629
rect 29178 17620 29184 17632
rect 29236 17620 29242 17672
rect 29270 17620 29276 17672
rect 29328 17660 29334 17672
rect 29917 17663 29975 17669
rect 29917 17660 29929 17663
rect 29328 17632 29929 17660
rect 29328 17620 29334 17632
rect 29917 17629 29929 17632
rect 29963 17629 29975 17663
rect 29917 17623 29975 17629
rect 30834 17620 30840 17672
rect 30892 17660 30898 17672
rect 31113 17663 31171 17669
rect 31113 17660 31125 17663
rect 30892 17632 31125 17660
rect 30892 17620 30898 17632
rect 31113 17629 31125 17632
rect 31159 17629 31171 17663
rect 31113 17623 31171 17629
rect 31297 17663 31355 17669
rect 31297 17629 31309 17663
rect 31343 17660 31355 17663
rect 31386 17660 31392 17672
rect 31343 17632 31392 17660
rect 31343 17629 31355 17632
rect 31297 17623 31355 17629
rect 31386 17620 31392 17632
rect 31444 17620 31450 17672
rect 32306 17620 32312 17672
rect 32364 17660 32370 17672
rect 32493 17663 32551 17669
rect 32493 17660 32505 17663
rect 32364 17632 32505 17660
rect 32364 17620 32370 17632
rect 32493 17629 32505 17632
rect 32539 17629 32551 17663
rect 33226 17660 33232 17672
rect 33187 17632 33232 17660
rect 32493 17623 32551 17629
rect 33226 17620 33232 17632
rect 33284 17620 33290 17672
rect 33410 17660 33416 17672
rect 33371 17632 33416 17660
rect 33410 17620 33416 17632
rect 33468 17620 33474 17672
rect 33502 17620 33508 17672
rect 33560 17660 33566 17672
rect 33643 17663 33701 17669
rect 33560 17632 33605 17660
rect 33560 17620 33566 17632
rect 33643 17629 33655 17663
rect 33689 17660 33701 17663
rect 34790 17660 34796 17672
rect 33689 17632 34796 17660
rect 33689 17629 33701 17632
rect 33643 17623 33701 17629
rect 34790 17620 34796 17632
rect 34848 17620 34854 17672
rect 35621 17663 35679 17669
rect 35621 17629 35633 17663
rect 35667 17629 35679 17663
rect 35621 17623 35679 17629
rect 35713 17663 35771 17669
rect 35713 17629 35725 17663
rect 35759 17629 35771 17663
rect 35713 17623 35771 17629
rect 35526 17592 35532 17604
rect 34808 17564 35532 17592
rect 28813 17527 28871 17533
rect 28813 17493 28825 17527
rect 28859 17524 28871 17527
rect 29086 17524 29092 17536
rect 28859 17496 29092 17524
rect 28859 17493 28871 17496
rect 28813 17487 28871 17493
rect 29086 17484 29092 17496
rect 29144 17484 29150 17536
rect 31386 17484 31392 17536
rect 31444 17524 31450 17536
rect 33962 17524 33968 17536
rect 31444 17496 33968 17524
rect 31444 17484 31450 17496
rect 33962 17484 33968 17496
rect 34020 17484 34026 17536
rect 34698 17484 34704 17536
rect 34756 17524 34762 17536
rect 34808 17533 34836 17564
rect 35526 17552 35532 17564
rect 35584 17592 35590 17604
rect 35636 17592 35664 17623
rect 35584 17564 35664 17592
rect 35584 17552 35590 17564
rect 34793 17527 34851 17533
rect 34793 17524 34805 17527
rect 34756 17496 34805 17524
rect 34756 17484 34762 17496
rect 34793 17493 34805 17496
rect 34839 17493 34851 17527
rect 34793 17487 34851 17493
rect 35618 17484 35624 17536
rect 35676 17524 35682 17536
rect 35728 17524 35756 17623
rect 35802 17620 35808 17672
rect 35860 17660 35866 17672
rect 36004 17669 36032 17700
rect 35989 17663 36047 17669
rect 35860 17632 35905 17660
rect 35860 17620 35866 17632
rect 35989 17629 36001 17663
rect 36035 17629 36047 17663
rect 35989 17623 36047 17629
rect 36817 17663 36875 17669
rect 36817 17629 36829 17663
rect 36863 17660 36875 17663
rect 37458 17660 37464 17672
rect 36863 17632 37464 17660
rect 36863 17629 36875 17632
rect 36817 17623 36875 17629
rect 37458 17620 37464 17632
rect 37516 17620 37522 17672
rect 37826 17660 37832 17672
rect 37787 17632 37832 17660
rect 37826 17620 37832 17632
rect 37884 17620 37890 17672
rect 38010 17660 38016 17672
rect 37971 17632 38016 17660
rect 38010 17620 38016 17632
rect 38068 17620 38074 17672
rect 38123 17669 38151 17768
rect 38212 17669 38240 17836
rect 38286 17824 38292 17836
rect 38344 17824 38350 17876
rect 38473 17867 38531 17873
rect 38473 17833 38485 17867
rect 38519 17864 38531 17867
rect 38654 17864 38660 17876
rect 38519 17836 38660 17864
rect 38519 17833 38531 17836
rect 38473 17827 38531 17833
rect 38654 17824 38660 17836
rect 38712 17824 38718 17876
rect 38108 17663 38166 17669
rect 38108 17629 38120 17663
rect 38154 17629 38166 17663
rect 38108 17623 38166 17629
rect 38197 17663 38255 17669
rect 38197 17629 38209 17663
rect 38243 17629 38255 17663
rect 38197 17623 38255 17629
rect 38746 17620 38752 17672
rect 38804 17660 38810 17672
rect 39117 17663 39175 17669
rect 39117 17660 39129 17663
rect 38804 17632 39129 17660
rect 38804 17620 38810 17632
rect 39117 17629 39129 17632
rect 39163 17660 39175 17663
rect 40402 17660 40408 17672
rect 39163 17632 40408 17660
rect 39163 17629 39175 17632
rect 39117 17623 39175 17629
rect 40402 17620 40408 17632
rect 40460 17620 40466 17672
rect 36630 17592 36636 17604
rect 36591 17564 36636 17592
rect 36630 17552 36636 17564
rect 36688 17552 36694 17604
rect 37476 17592 37504 17620
rect 37734 17592 37740 17604
rect 37476 17564 37740 17592
rect 37734 17552 37740 17564
rect 37792 17552 37798 17604
rect 38838 17552 38844 17604
rect 38896 17592 38902 17604
rect 38933 17595 38991 17601
rect 38933 17592 38945 17595
rect 38896 17564 38945 17592
rect 38896 17552 38902 17564
rect 38933 17561 38945 17564
rect 38979 17561 38991 17595
rect 39298 17592 39304 17604
rect 39259 17564 39304 17592
rect 38933 17555 38991 17561
rect 39298 17552 39304 17564
rect 39356 17552 39362 17604
rect 35676 17496 35756 17524
rect 35676 17484 35682 17496
rect 35802 17484 35808 17536
rect 35860 17524 35866 17536
rect 36449 17527 36507 17533
rect 36449 17524 36461 17527
rect 35860 17496 36461 17524
rect 35860 17484 35866 17496
rect 36449 17493 36461 17496
rect 36495 17493 36507 17527
rect 36449 17487 36507 17493
rect 1104 17434 68816 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 68816 17434
rect 1104 17360 68816 17382
rect 2406 17280 2412 17332
rect 2464 17320 2470 17332
rect 4617 17323 4675 17329
rect 4617 17320 4629 17323
rect 2464 17292 4629 17320
rect 2464 17280 2470 17292
rect 4617 17289 4629 17292
rect 4663 17320 4675 17323
rect 5813 17323 5871 17329
rect 4663 17292 5580 17320
rect 4663 17289 4675 17292
rect 4617 17283 4675 17289
rect 2314 17212 2320 17264
rect 2372 17252 2378 17264
rect 2372 17224 5491 17252
rect 2372 17212 2378 17224
rect 1854 17184 1860 17196
rect 1815 17156 1860 17184
rect 1854 17144 1860 17156
rect 1912 17144 1918 17196
rect 2041 17187 2099 17193
rect 2041 17153 2053 17187
rect 2087 17184 2099 17187
rect 5074 17184 5080 17196
rect 2087 17156 5080 17184
rect 2087 17153 2099 17156
rect 2041 17147 2099 17153
rect 5074 17144 5080 17156
rect 5132 17144 5138 17196
rect 5463 17193 5491 17224
rect 5552 17193 5580 17292
rect 5813 17289 5825 17323
rect 5859 17320 5871 17323
rect 6914 17320 6920 17332
rect 5859 17292 6920 17320
rect 5859 17289 5871 17292
rect 5813 17283 5871 17289
rect 6914 17280 6920 17292
rect 6972 17280 6978 17332
rect 14550 17320 14556 17332
rect 7024 17292 14556 17320
rect 6362 17212 6368 17264
rect 6420 17252 6426 17264
rect 6549 17255 6607 17261
rect 6549 17252 6561 17255
rect 6420 17224 6561 17252
rect 6420 17212 6426 17224
rect 6549 17221 6561 17224
rect 6595 17221 6607 17255
rect 6549 17215 6607 17221
rect 6638 17212 6644 17264
rect 6696 17252 6702 17264
rect 7024 17252 7052 17292
rect 14550 17280 14556 17292
rect 14608 17320 14614 17332
rect 15657 17323 15715 17329
rect 14608 17292 15148 17320
rect 14608 17280 14614 17292
rect 10962 17252 10968 17264
rect 6696 17224 7052 17252
rect 8312 17224 10968 17252
rect 6696 17212 6702 17224
rect 5169 17187 5227 17193
rect 5332 17187 5390 17193
rect 5169 17153 5181 17187
rect 5215 17153 5227 17187
rect 5169 17147 5227 17153
rect 5276 17159 5344 17187
rect 4982 17076 4988 17128
rect 5040 17116 5046 17128
rect 5184 17116 5212 17147
rect 5040 17088 5212 17116
rect 5040 17076 5046 17088
rect 5276 17048 5304 17159
rect 5332 17153 5344 17159
rect 5378 17153 5390 17187
rect 5332 17147 5390 17153
rect 5445 17187 5503 17193
rect 5445 17153 5457 17187
rect 5491 17153 5503 17187
rect 5445 17147 5503 17153
rect 5537 17187 5595 17193
rect 5537 17153 5549 17187
rect 5583 17153 5595 17187
rect 5537 17147 5595 17153
rect 5463 17116 5491 17147
rect 6270 17144 6276 17196
rect 6328 17184 6334 17196
rect 6733 17187 6791 17193
rect 6733 17184 6745 17187
rect 6328 17156 6745 17184
rect 6328 17144 6334 17156
rect 6733 17153 6745 17156
rect 6779 17184 6791 17187
rect 6914 17184 6920 17196
rect 6779 17156 6920 17184
rect 6779 17153 6791 17156
rect 6733 17147 6791 17153
rect 6914 17144 6920 17156
rect 6972 17144 6978 17196
rect 7098 17144 7104 17196
rect 7156 17184 7162 17196
rect 7193 17187 7251 17193
rect 7193 17184 7205 17187
rect 7156 17156 7205 17184
rect 7156 17144 7162 17156
rect 7193 17153 7205 17156
rect 7239 17153 7251 17187
rect 7374 17184 7380 17196
rect 7335 17156 7380 17184
rect 7193 17147 7251 17153
rect 7374 17144 7380 17156
rect 7432 17144 7438 17196
rect 7469 17187 7527 17193
rect 7469 17153 7481 17187
rect 7515 17153 7527 17187
rect 7469 17147 7527 17153
rect 5463 17088 6914 17116
rect 6365 17051 6423 17057
rect 6365 17048 6377 17051
rect 5276 17020 6377 17048
rect 6365 17017 6377 17020
rect 6411 17017 6423 17051
rect 6365 17011 6423 17017
rect 2222 16980 2228 16992
rect 2183 16952 2228 16980
rect 2222 16940 2228 16952
rect 2280 16940 2286 16992
rect 6886 16980 6914 17088
rect 7484 16980 7512 17147
rect 7558 17144 7564 17196
rect 7616 17184 7622 17196
rect 7616 17156 7661 17184
rect 7616 17144 7622 17156
rect 8018 17144 8024 17196
rect 8076 17184 8082 17196
rect 8312 17193 8340 17224
rect 10962 17212 10968 17224
rect 11020 17252 11026 17264
rect 12434 17252 12440 17264
rect 11020 17224 12440 17252
rect 11020 17212 11026 17224
rect 8304 17187 8362 17193
rect 8304 17184 8316 17187
rect 8076 17156 8316 17184
rect 8076 17144 8082 17156
rect 8304 17153 8316 17156
rect 8350 17153 8362 17187
rect 8553 17187 8611 17193
rect 8553 17184 8565 17187
rect 8304 17147 8362 17153
rect 8404 17156 8565 17184
rect 7837 17119 7895 17125
rect 7837 17085 7849 17119
rect 7883 17116 7895 17119
rect 8404 17116 8432 17156
rect 8553 17153 8565 17156
rect 8599 17153 8611 17187
rect 10502 17184 10508 17196
rect 10463 17156 10508 17184
rect 8553 17147 8611 17153
rect 10502 17144 10508 17156
rect 10560 17144 10566 17196
rect 11532 17193 11560 17224
rect 12434 17212 12440 17224
rect 12492 17212 12498 17264
rect 12894 17212 12900 17264
rect 12952 17252 12958 17264
rect 13446 17252 13452 17264
rect 12952 17224 13452 17252
rect 12952 17212 12958 17224
rect 13446 17212 13452 17224
rect 13504 17252 13510 17264
rect 13504 17224 13768 17252
rect 13504 17212 13510 17224
rect 10689 17187 10747 17193
rect 10689 17153 10701 17187
rect 10735 17153 10747 17187
rect 10689 17147 10747 17153
rect 11517 17187 11575 17193
rect 11517 17153 11529 17187
rect 11563 17153 11575 17187
rect 11517 17147 11575 17153
rect 7883 17088 8432 17116
rect 7883 17085 7895 17088
rect 7837 17079 7895 17085
rect 10704 17048 10732 17147
rect 11606 17144 11612 17196
rect 11664 17184 11670 17196
rect 11773 17187 11831 17193
rect 11773 17184 11785 17187
rect 11664 17156 11785 17184
rect 11664 17144 11670 17156
rect 11773 17153 11785 17156
rect 11819 17153 11831 17187
rect 11773 17147 11831 17153
rect 13262 17144 13268 17196
rect 13320 17184 13326 17196
rect 13357 17187 13415 17193
rect 13357 17184 13369 17187
rect 13320 17156 13369 17184
rect 13320 17144 13326 17156
rect 13357 17153 13369 17156
rect 13403 17153 13415 17187
rect 13538 17184 13544 17196
rect 13499 17156 13544 17184
rect 13357 17147 13415 17153
rect 13538 17144 13544 17156
rect 13596 17144 13602 17196
rect 13740 17193 13768 17224
rect 15120 17193 15148 17292
rect 15657 17289 15669 17323
rect 15703 17320 15715 17323
rect 15838 17320 15844 17332
rect 15703 17292 15844 17320
rect 15703 17289 15715 17292
rect 15657 17283 15715 17289
rect 15838 17280 15844 17292
rect 15896 17280 15902 17332
rect 17034 17320 17040 17332
rect 16995 17292 17040 17320
rect 17034 17280 17040 17292
rect 17092 17280 17098 17332
rect 24486 17280 24492 17332
rect 24544 17320 24550 17332
rect 25314 17320 25320 17332
rect 24544 17292 25320 17320
rect 24544 17280 24550 17292
rect 25314 17280 25320 17292
rect 25372 17280 25378 17332
rect 27338 17320 27344 17332
rect 27299 17292 27344 17320
rect 27338 17280 27344 17292
rect 27396 17280 27402 17332
rect 27706 17320 27712 17332
rect 27641 17292 27712 17320
rect 15930 17212 15936 17264
rect 15988 17252 15994 17264
rect 16853 17255 16911 17261
rect 16853 17252 16865 17255
rect 15988 17224 16865 17252
rect 15988 17212 15994 17224
rect 16853 17221 16865 17224
rect 16899 17221 16911 17255
rect 16853 17215 16911 17221
rect 18782 17212 18788 17264
rect 18840 17252 18846 17264
rect 20717 17255 20775 17261
rect 18840 17224 19288 17252
rect 18840 17212 18846 17224
rect 13633 17187 13691 17193
rect 13633 17153 13645 17187
rect 13679 17153 13691 17187
rect 13633 17147 13691 17153
rect 13725 17187 13783 17193
rect 13725 17153 13737 17187
rect 13771 17184 13783 17187
rect 14461 17187 14519 17193
rect 14461 17184 14473 17187
rect 13771 17156 14473 17184
rect 13771 17153 13783 17156
rect 13725 17147 13783 17153
rect 14461 17153 14473 17156
rect 14507 17153 14519 17187
rect 14461 17147 14519 17153
rect 15105 17187 15163 17193
rect 15105 17153 15117 17187
rect 15151 17184 15163 17187
rect 15838 17184 15844 17196
rect 15151 17156 15844 17184
rect 15151 17153 15163 17156
rect 15105 17147 15163 17153
rect 12710 17076 12716 17128
rect 12768 17116 12774 17128
rect 13648 17116 13676 17147
rect 15838 17144 15844 17156
rect 15896 17144 15902 17196
rect 16666 17184 16672 17196
rect 16627 17156 16672 17184
rect 16666 17144 16672 17156
rect 16724 17144 16730 17196
rect 18874 17184 18880 17196
rect 18835 17156 18880 17184
rect 18874 17144 18880 17156
rect 18932 17144 18938 17196
rect 19260 17193 19288 17224
rect 20717 17221 20729 17255
rect 20763 17252 20775 17255
rect 26510 17252 26516 17264
rect 20763 17224 26516 17252
rect 20763 17221 20775 17224
rect 20717 17215 20775 17221
rect 26510 17212 26516 17224
rect 26568 17212 26574 17264
rect 27641 17252 27669 17292
rect 27706 17280 27712 17292
rect 27764 17280 27770 17332
rect 27798 17280 27804 17332
rect 27856 17320 27862 17332
rect 29270 17320 29276 17332
rect 27856 17292 29276 17320
rect 27856 17280 27862 17292
rect 29270 17280 29276 17292
rect 29328 17280 29334 17332
rect 31481 17323 31539 17329
rect 31481 17289 31493 17323
rect 31527 17320 31539 17323
rect 31938 17320 31944 17332
rect 31527 17292 31944 17320
rect 31527 17289 31539 17292
rect 31481 17283 31539 17289
rect 31938 17280 31944 17292
rect 31996 17280 32002 17332
rect 33045 17323 33103 17329
rect 33045 17320 33057 17323
rect 32324 17292 33057 17320
rect 27641 17224 27752 17252
rect 27724 17196 27752 17224
rect 27890 17212 27896 17264
rect 27948 17252 27954 17264
rect 28445 17255 28503 17261
rect 28445 17252 28457 17255
rect 27948 17224 28457 17252
rect 27948 17212 27954 17224
rect 28445 17221 28457 17224
rect 28491 17221 28503 17255
rect 28626 17252 28632 17264
rect 28587 17224 28632 17252
rect 28445 17215 28503 17221
rect 28626 17212 28632 17224
rect 28684 17212 28690 17264
rect 29638 17252 29644 17264
rect 29599 17224 29644 17252
rect 29638 17212 29644 17224
rect 29696 17212 29702 17264
rect 31386 17212 31392 17264
rect 31444 17252 31450 17264
rect 31754 17252 31760 17264
rect 31444 17224 31760 17252
rect 31444 17212 31450 17224
rect 31754 17212 31760 17224
rect 31812 17252 31818 17264
rect 32324 17261 32352 17292
rect 33045 17289 33057 17292
rect 33091 17289 33103 17323
rect 33045 17283 33103 17289
rect 37734 17280 37740 17332
rect 37792 17320 37798 17332
rect 38838 17320 38844 17332
rect 37792 17292 38844 17320
rect 37792 17280 37798 17292
rect 38838 17280 38844 17292
rect 38896 17280 38902 17332
rect 32125 17255 32183 17261
rect 32125 17252 32137 17255
rect 31812 17224 32137 17252
rect 31812 17212 31818 17224
rect 32125 17221 32137 17224
rect 32171 17221 32183 17255
rect 32125 17215 32183 17221
rect 32309 17255 32367 17261
rect 32309 17221 32321 17255
rect 32355 17221 32367 17255
rect 32309 17215 32367 17221
rect 19061 17187 19119 17193
rect 19061 17153 19073 17187
rect 19107 17153 19119 17187
rect 19061 17147 19119 17153
rect 19153 17187 19211 17193
rect 19153 17153 19165 17187
rect 19199 17153 19211 17187
rect 19153 17147 19211 17153
rect 19245 17187 19303 17193
rect 19245 17153 19257 17187
rect 19291 17153 19303 17187
rect 19245 17147 19303 17153
rect 12768 17088 13676 17116
rect 12768 17076 12774 17088
rect 16850 17076 16856 17128
rect 16908 17116 16914 17128
rect 17497 17119 17555 17125
rect 17497 17116 17509 17119
rect 16908 17088 17509 17116
rect 16908 17076 16914 17088
rect 17497 17085 17509 17088
rect 17543 17085 17555 17119
rect 17497 17079 17555 17085
rect 18322 17076 18328 17128
rect 18380 17116 18386 17128
rect 19076 17116 19104 17147
rect 18380 17088 19104 17116
rect 18380 17076 18386 17088
rect 12897 17051 12955 17057
rect 10704 17020 11560 17048
rect 7834 16980 7840 16992
rect 6886 16952 7840 16980
rect 7834 16940 7840 16952
rect 7892 16940 7898 16992
rect 9677 16983 9735 16989
rect 9677 16949 9689 16983
rect 9723 16980 9735 16983
rect 9858 16980 9864 16992
rect 9723 16952 9864 16980
rect 9723 16949 9735 16952
rect 9677 16943 9735 16949
rect 9858 16940 9864 16952
rect 9916 16940 9922 16992
rect 10410 16940 10416 16992
rect 10468 16980 10474 16992
rect 10873 16983 10931 16989
rect 10873 16980 10885 16983
rect 10468 16952 10885 16980
rect 10468 16940 10474 16952
rect 10873 16949 10885 16952
rect 10919 16949 10931 16983
rect 11532 16980 11560 17020
rect 12897 17017 12909 17051
rect 12943 17048 12955 17051
rect 19168 17048 19196 17147
rect 20070 17144 20076 17196
rect 20128 17184 20134 17196
rect 20579 17187 20637 17193
rect 20579 17184 20591 17187
rect 20128 17156 20591 17184
rect 20128 17144 20134 17156
rect 20579 17153 20591 17156
rect 20625 17153 20637 17187
rect 20806 17184 20812 17196
rect 20767 17156 20812 17184
rect 20579 17147 20637 17153
rect 20806 17144 20812 17156
rect 20864 17144 20870 17196
rect 20898 17144 20904 17196
rect 20956 17193 20962 17196
rect 20956 17187 20995 17193
rect 20983 17153 20995 17187
rect 20956 17147 20995 17153
rect 21085 17187 21143 17193
rect 21085 17153 21097 17187
rect 21131 17153 21143 17187
rect 21085 17147 21143 17153
rect 20956 17144 20962 17147
rect 21100 17116 21128 17147
rect 22094 17144 22100 17196
rect 22152 17184 22158 17196
rect 23302 17187 23360 17193
rect 23302 17184 23314 17187
rect 22152 17156 23314 17184
rect 22152 17144 22158 17156
rect 23302 17153 23314 17156
rect 23348 17153 23360 17187
rect 24486 17184 24492 17196
rect 24447 17156 24492 17184
rect 23302 17147 23360 17153
rect 24486 17144 24492 17156
rect 24544 17144 24550 17196
rect 25130 17184 25136 17196
rect 25091 17156 25136 17184
rect 25130 17144 25136 17156
rect 25188 17144 25194 17196
rect 25317 17187 25375 17193
rect 25317 17153 25329 17187
rect 25363 17153 25375 17187
rect 25317 17147 25375 17153
rect 26421 17187 26479 17193
rect 26421 17153 26433 17187
rect 26467 17184 26479 17187
rect 27522 17184 27528 17196
rect 26467 17156 27528 17184
rect 26467 17153 26479 17156
rect 26421 17147 26479 17153
rect 23566 17116 23572 17128
rect 19444 17088 21128 17116
rect 23527 17088 23572 17116
rect 19444 17057 19472 17088
rect 23566 17076 23572 17088
rect 23624 17076 23630 17128
rect 24302 17076 24308 17128
rect 24360 17116 24366 17128
rect 25332 17116 25360 17147
rect 27522 17144 27528 17156
rect 27580 17184 27586 17196
rect 27617 17187 27675 17193
rect 27617 17184 27629 17187
rect 27580 17156 27629 17184
rect 27580 17144 27586 17156
rect 27617 17153 27629 17156
rect 27663 17153 27675 17187
rect 27617 17147 27675 17153
rect 27706 17190 27764 17196
rect 27706 17156 27718 17190
rect 27752 17156 27764 17190
rect 27706 17150 27764 17156
rect 27798 17144 27804 17196
rect 27856 17184 27862 17196
rect 27985 17187 28043 17193
rect 27856 17156 27901 17184
rect 27856 17144 27862 17156
rect 27985 17153 27997 17187
rect 28031 17153 28043 17187
rect 27985 17147 28043 17153
rect 28813 17187 28871 17193
rect 28813 17153 28825 17187
rect 28859 17184 28871 17187
rect 29086 17184 29092 17196
rect 28859 17156 29092 17184
rect 28859 17153 28871 17156
rect 28813 17147 28871 17153
rect 24360 17088 25360 17116
rect 24360 17076 24366 17088
rect 12943 17020 19196 17048
rect 19429 17051 19487 17057
rect 12943 17017 12955 17020
rect 12897 17011 12955 17017
rect 19429 17017 19441 17051
rect 19475 17017 19487 17051
rect 19429 17011 19487 17017
rect 12912 16980 12940 17011
rect 20898 17008 20904 17060
rect 20956 17048 20962 17060
rect 22189 17051 22247 17057
rect 22189 17048 22201 17051
rect 20956 17020 22201 17048
rect 20956 17008 20962 17020
rect 22189 17017 22201 17020
rect 22235 17017 22247 17051
rect 22189 17011 22247 17017
rect 24673 17051 24731 17057
rect 24673 17017 24685 17051
rect 24719 17048 24731 17051
rect 25682 17048 25688 17060
rect 24719 17020 25688 17048
rect 24719 17017 24731 17020
rect 24673 17011 24731 17017
rect 25682 17008 25688 17020
rect 25740 17048 25746 17060
rect 26602 17048 26608 17060
rect 25740 17020 26608 17048
rect 25740 17008 25746 17020
rect 26602 17008 26608 17020
rect 26660 17008 26666 17060
rect 26786 17008 26792 17060
rect 26844 17048 26850 17060
rect 28000 17048 28028 17147
rect 29086 17144 29092 17156
rect 29144 17144 29150 17196
rect 29546 17184 29552 17196
rect 29507 17156 29552 17184
rect 29546 17144 29552 17156
rect 29604 17144 29610 17196
rect 29733 17187 29791 17193
rect 29733 17153 29745 17187
rect 29779 17153 29791 17187
rect 29733 17147 29791 17153
rect 29917 17187 29975 17193
rect 29917 17153 29929 17187
rect 29963 17184 29975 17187
rect 30006 17184 30012 17196
rect 29963 17156 30012 17184
rect 29963 17153 29975 17156
rect 29917 17147 29975 17153
rect 28902 17076 28908 17128
rect 28960 17116 28966 17128
rect 29748 17116 29776 17147
rect 30006 17144 30012 17156
rect 30064 17144 30070 17196
rect 30837 17187 30895 17193
rect 30837 17153 30849 17187
rect 30883 17153 30895 17187
rect 31018 17184 31024 17196
rect 30979 17156 31024 17184
rect 30837 17147 30895 17153
rect 28960 17088 29776 17116
rect 30852 17116 30880 17147
rect 31018 17144 31024 17156
rect 31076 17144 31082 17196
rect 31110 17144 31116 17196
rect 31168 17184 31174 17196
rect 31251 17187 31309 17193
rect 31168 17156 31213 17184
rect 31168 17144 31174 17156
rect 31251 17153 31263 17187
rect 31297 17184 31309 17187
rect 31478 17184 31484 17196
rect 31297 17156 31484 17184
rect 31297 17153 31309 17156
rect 31251 17147 31309 17153
rect 31478 17144 31484 17156
rect 31536 17144 31542 17196
rect 30926 17116 30932 17128
rect 30852 17088 30932 17116
rect 28960 17076 28966 17088
rect 30926 17076 30932 17088
rect 30984 17076 30990 17128
rect 26844 17020 29500 17048
rect 26844 17008 26850 17020
rect 13998 16980 14004 16992
rect 11532 16952 12940 16980
rect 13959 16952 14004 16980
rect 10873 16943 10931 16949
rect 13998 16940 14004 16952
rect 14056 16940 14062 16992
rect 20441 16983 20499 16989
rect 20441 16949 20453 16983
rect 20487 16980 20499 16983
rect 20622 16980 20628 16992
rect 20487 16952 20628 16980
rect 20487 16949 20499 16952
rect 20441 16943 20499 16949
rect 20622 16940 20628 16952
rect 20680 16940 20686 16992
rect 25501 16983 25559 16989
rect 25501 16949 25513 16983
rect 25547 16980 25559 16983
rect 26234 16980 26240 16992
rect 25547 16952 26240 16980
rect 25547 16949 25559 16952
rect 25501 16943 25559 16949
rect 26234 16940 26240 16952
rect 26292 16940 26298 16992
rect 29362 16980 29368 16992
rect 29323 16952 29368 16980
rect 29362 16940 29368 16952
rect 29420 16940 29426 16992
rect 29472 16980 29500 17020
rect 29730 17008 29736 17060
rect 29788 17048 29794 17060
rect 32324 17048 32352 17215
rect 32950 17212 32956 17264
rect 33008 17252 33014 17264
rect 38473 17255 38531 17261
rect 33008 17224 34376 17252
rect 33008 17212 33014 17224
rect 33134 17144 33140 17196
rect 33192 17184 33198 17196
rect 34158 17187 34216 17193
rect 34158 17184 34170 17187
rect 33192 17156 34170 17184
rect 33192 17144 33198 17156
rect 34158 17153 34170 17156
rect 34204 17153 34216 17187
rect 34158 17147 34216 17153
rect 34348 17116 34376 17224
rect 37384 17224 38151 17252
rect 37384 17196 37412 17224
rect 38123 17196 38151 17224
rect 38473 17221 38485 17255
rect 38519 17252 38531 17255
rect 39454 17255 39512 17261
rect 39454 17252 39466 17255
rect 38519 17224 39466 17252
rect 38519 17221 38531 17224
rect 38473 17215 38531 17221
rect 39454 17221 39466 17224
rect 39500 17221 39512 17255
rect 39454 17215 39512 17221
rect 34425 17187 34483 17193
rect 34425 17153 34437 17187
rect 34471 17184 34483 17187
rect 35342 17184 35348 17196
rect 34471 17156 35348 17184
rect 34471 17153 34483 17156
rect 34425 17147 34483 17153
rect 35342 17144 35348 17156
rect 35400 17144 35406 17196
rect 35529 17187 35587 17193
rect 35529 17153 35541 17187
rect 35575 17184 35587 17187
rect 35618 17184 35624 17196
rect 35575 17156 35624 17184
rect 35575 17153 35587 17156
rect 35529 17147 35587 17153
rect 35618 17144 35624 17156
rect 35676 17184 35682 17196
rect 37366 17184 37372 17196
rect 35676 17156 37372 17184
rect 35676 17144 35682 17156
rect 37366 17144 37372 17156
rect 37424 17144 37430 17196
rect 37826 17184 37832 17196
rect 37787 17156 37832 17184
rect 37826 17144 37832 17156
rect 37884 17144 37890 17196
rect 38013 17187 38071 17193
rect 38013 17153 38025 17187
rect 38059 17153 38071 17187
rect 38013 17147 38071 17153
rect 38108 17190 38166 17196
rect 38108 17156 38120 17190
rect 38154 17156 38166 17190
rect 38108 17150 38166 17156
rect 38217 17187 38275 17193
rect 38217 17153 38229 17187
rect 38263 17184 38275 17187
rect 38378 17184 38384 17196
rect 38263 17156 38384 17184
rect 38263 17153 38275 17156
rect 38217 17147 38275 17153
rect 35253 17119 35311 17125
rect 35253 17116 35265 17119
rect 34348 17088 35265 17116
rect 35253 17085 35265 17088
rect 35299 17085 35311 17119
rect 35253 17079 35311 17085
rect 29788 17020 32352 17048
rect 38028 17048 38056 17147
rect 38378 17144 38384 17156
rect 38436 17144 38442 17196
rect 39022 17144 39028 17196
rect 39080 17184 39086 17196
rect 39209 17187 39267 17193
rect 39209 17184 39221 17187
rect 39080 17156 39221 17184
rect 39080 17144 39086 17156
rect 39209 17153 39221 17156
rect 39255 17153 39267 17187
rect 39209 17147 39267 17153
rect 38102 17048 38108 17060
rect 38028 17020 38108 17048
rect 29788 17008 29794 17020
rect 38102 17008 38108 17020
rect 38160 17008 38166 17060
rect 67634 17048 67640 17060
rect 67595 17020 67640 17048
rect 67634 17008 67640 17020
rect 67692 17008 67698 17060
rect 31018 16980 31024 16992
rect 29472 16952 31024 16980
rect 31018 16940 31024 16952
rect 31076 16940 31082 16992
rect 32490 16980 32496 16992
rect 32451 16952 32496 16980
rect 32490 16940 32496 16952
rect 32548 16940 32554 16992
rect 37274 16980 37280 16992
rect 37235 16952 37280 16980
rect 37274 16940 37280 16952
rect 37332 16940 37338 16992
rect 40586 16980 40592 16992
rect 40547 16952 40592 16980
rect 40586 16940 40592 16952
rect 40644 16940 40650 16992
rect 1104 16890 68816 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 65654 16890
rect 65706 16838 65718 16890
rect 65770 16838 65782 16890
rect 65834 16838 65846 16890
rect 65898 16838 65910 16890
rect 65962 16838 68816 16890
rect 1104 16816 68816 16838
rect 3234 16776 3240 16788
rect 3195 16748 3240 16776
rect 3234 16736 3240 16748
rect 3292 16736 3298 16788
rect 5074 16736 5080 16788
rect 5132 16776 5138 16788
rect 5169 16779 5227 16785
rect 5169 16776 5181 16779
rect 5132 16748 5181 16776
rect 5132 16736 5138 16748
rect 5169 16745 5181 16748
rect 5215 16745 5227 16779
rect 5169 16739 5227 16745
rect 7374 16736 7380 16788
rect 7432 16776 7438 16788
rect 7837 16779 7895 16785
rect 7837 16776 7849 16779
rect 7432 16748 7849 16776
rect 7432 16736 7438 16748
rect 7837 16745 7849 16748
rect 7883 16745 7895 16779
rect 7837 16739 7895 16745
rect 10778 16736 10784 16788
rect 10836 16776 10842 16788
rect 11333 16779 11391 16785
rect 11333 16776 11345 16779
rect 10836 16748 11345 16776
rect 10836 16736 10842 16748
rect 11333 16745 11345 16748
rect 11379 16745 11391 16779
rect 15194 16776 15200 16788
rect 11333 16739 11391 16745
rect 14108 16748 15200 16776
rect 5905 16711 5963 16717
rect 5905 16677 5917 16711
rect 5951 16708 5963 16711
rect 5951 16680 6776 16708
rect 5951 16677 5963 16680
rect 5905 16671 5963 16677
rect 6638 16640 6644 16652
rect 5736 16612 6644 16640
rect 2038 16572 2044 16584
rect 1999 16544 2044 16572
rect 2038 16532 2044 16544
rect 2096 16532 2102 16584
rect 2222 16581 2228 16584
rect 2220 16572 2228 16581
rect 2183 16544 2228 16572
rect 2220 16535 2228 16544
rect 2222 16532 2228 16535
rect 2280 16532 2286 16584
rect 2455 16575 2513 16581
rect 2320 16569 2378 16575
rect 2320 16535 2332 16569
rect 2366 16535 2378 16569
rect 2455 16541 2467 16575
rect 2501 16572 2513 16575
rect 3234 16572 3240 16584
rect 2501 16544 3240 16572
rect 2501 16541 2513 16544
rect 2455 16535 2513 16541
rect 2320 16529 2378 16535
rect 3234 16532 3240 16544
rect 3292 16532 3298 16584
rect 3786 16572 3792 16584
rect 3747 16544 3792 16572
rect 3786 16532 3792 16544
rect 3844 16532 3850 16584
rect 5736 16581 5764 16612
rect 6638 16600 6644 16612
rect 6696 16600 6702 16652
rect 6748 16640 6776 16680
rect 7650 16668 7656 16720
rect 7708 16708 7714 16720
rect 8297 16711 8355 16717
rect 8297 16708 8309 16711
rect 7708 16680 8309 16708
rect 7708 16668 7714 16680
rect 8297 16677 8309 16680
rect 8343 16677 8355 16711
rect 8297 16671 8355 16677
rect 12406 16680 12664 16708
rect 8110 16640 8116 16652
rect 6748 16612 8116 16640
rect 8110 16600 8116 16612
rect 8168 16640 8174 16652
rect 8754 16640 8760 16652
rect 8168 16612 8760 16640
rect 8168 16600 8174 16612
rect 8754 16600 8760 16612
rect 8812 16600 8818 16652
rect 9398 16600 9404 16652
rect 9456 16640 9462 16652
rect 12406 16640 12434 16680
rect 9456 16612 12434 16640
rect 9456 16600 9462 16612
rect 5721 16575 5779 16581
rect 5721 16541 5733 16575
rect 5767 16541 5779 16575
rect 5721 16535 5779 16541
rect 6362 16532 6368 16584
rect 6420 16572 6426 16584
rect 6457 16575 6515 16581
rect 6457 16572 6469 16575
rect 6420 16544 6469 16572
rect 6420 16532 6426 16544
rect 6457 16541 6469 16544
rect 6503 16541 6515 16575
rect 6457 16535 6515 16541
rect 6546 16532 6552 16584
rect 6604 16572 6610 16584
rect 10244 16581 10272 16612
rect 6825 16575 6883 16581
rect 6825 16572 6837 16575
rect 6604 16544 6837 16572
rect 6604 16532 6610 16544
rect 6825 16541 6837 16544
rect 6871 16541 6883 16575
rect 6825 16535 6883 16541
rect 10229 16575 10287 16581
rect 10229 16541 10241 16575
rect 10275 16541 10287 16575
rect 10410 16572 10416 16584
rect 10371 16544 10416 16572
rect 10229 16535 10287 16541
rect 10410 16532 10416 16544
rect 10468 16532 10474 16584
rect 10502 16532 10508 16584
rect 10560 16572 10566 16584
rect 10643 16575 10701 16581
rect 10560 16544 10605 16572
rect 10560 16532 10566 16544
rect 10643 16541 10655 16575
rect 10689 16572 10701 16575
rect 10778 16572 10784 16584
rect 10689 16544 10784 16572
rect 10689 16541 10701 16544
rect 10643 16535 10701 16541
rect 10778 16532 10784 16544
rect 10836 16532 10842 16584
rect 12636 16581 12664 16680
rect 14108 16649 14136 16748
rect 15194 16736 15200 16748
rect 15252 16736 15258 16788
rect 15473 16779 15531 16785
rect 15473 16745 15485 16779
rect 15519 16776 15531 16779
rect 16022 16776 16028 16788
rect 15519 16748 16028 16776
rect 15519 16745 15531 16748
rect 15473 16739 15531 16745
rect 16022 16736 16028 16748
rect 16080 16736 16086 16788
rect 22094 16736 22100 16788
rect 22152 16776 22158 16788
rect 22152 16748 22197 16776
rect 22152 16736 22158 16748
rect 23566 16736 23572 16788
rect 23624 16776 23630 16788
rect 24394 16776 24400 16788
rect 23624 16748 24400 16776
rect 23624 16736 23630 16748
rect 24394 16736 24400 16748
rect 24452 16776 24458 16788
rect 24452 16748 25820 16776
rect 24452 16736 24458 16748
rect 16666 16668 16672 16720
rect 16724 16708 16730 16720
rect 19426 16708 19432 16720
rect 16724 16680 19432 16708
rect 16724 16668 16730 16680
rect 19426 16668 19432 16680
rect 19484 16708 19490 16720
rect 19610 16708 19616 16720
rect 19484 16680 19616 16708
rect 19484 16668 19490 16680
rect 19610 16668 19616 16680
rect 19668 16668 19674 16720
rect 20438 16668 20444 16720
rect 20496 16708 20502 16720
rect 20533 16711 20591 16717
rect 20533 16708 20545 16711
rect 20496 16680 20545 16708
rect 20496 16668 20502 16680
rect 20533 16677 20545 16680
rect 20579 16708 20591 16711
rect 21082 16708 21088 16720
rect 20579 16680 21088 16708
rect 20579 16677 20591 16680
rect 20533 16671 20591 16677
rect 21082 16668 21088 16680
rect 21140 16668 21146 16720
rect 21358 16668 21364 16720
rect 21416 16708 21422 16720
rect 23753 16711 23811 16717
rect 23753 16708 23765 16711
rect 21416 16680 23765 16708
rect 21416 16668 21422 16680
rect 23753 16677 23765 16680
rect 23799 16708 23811 16711
rect 24486 16708 24492 16720
rect 23799 16680 24492 16708
rect 23799 16677 23811 16680
rect 23753 16671 23811 16677
rect 24486 16668 24492 16680
rect 24544 16668 24550 16720
rect 14093 16643 14151 16649
rect 14093 16609 14105 16643
rect 14139 16609 14151 16643
rect 14093 16603 14151 16609
rect 15838 16600 15844 16652
rect 15896 16640 15902 16652
rect 16025 16643 16083 16649
rect 16025 16640 16037 16643
rect 15896 16612 16037 16640
rect 15896 16600 15902 16612
rect 16025 16609 16037 16612
rect 16071 16640 16083 16643
rect 16206 16640 16212 16652
rect 16071 16612 16212 16640
rect 16071 16609 16083 16612
rect 16025 16603 16083 16609
rect 16206 16600 16212 16612
rect 16264 16600 16270 16652
rect 17310 16640 17316 16652
rect 17144 16612 17316 16640
rect 12391 16575 12449 16581
rect 12391 16541 12403 16575
rect 12437 16541 12449 16575
rect 12391 16535 12449 16541
rect 12621 16575 12679 16581
rect 12621 16541 12633 16575
rect 12667 16572 12679 16575
rect 13262 16572 13268 16584
rect 12667 16544 13268 16572
rect 12667 16541 12679 16544
rect 12621 16535 12679 16541
rect 2332 16448 2360 16529
rect 2685 16507 2743 16513
rect 2685 16473 2697 16507
rect 2731 16504 2743 16507
rect 4034 16507 4092 16513
rect 4034 16504 4046 16507
rect 2731 16476 4046 16504
rect 2731 16473 2743 16476
rect 2685 16467 2743 16473
rect 4034 16473 4046 16476
rect 4080 16473 4092 16507
rect 4034 16467 4092 16473
rect 6270 16464 6276 16516
rect 6328 16504 6334 16516
rect 6641 16507 6699 16513
rect 6641 16504 6653 16507
rect 6328 16476 6653 16504
rect 6328 16464 6334 16476
rect 6641 16473 6653 16476
rect 6687 16473 6699 16507
rect 6641 16467 6699 16473
rect 6733 16507 6791 16513
rect 6733 16473 6745 16507
rect 6779 16504 6791 16507
rect 6779 16476 6868 16504
rect 6779 16473 6791 16476
rect 6733 16467 6791 16473
rect 2314 16396 2320 16448
rect 2372 16396 2378 16448
rect 5258 16396 5264 16448
rect 5316 16436 5322 16448
rect 6840 16436 6868 16476
rect 6914 16464 6920 16516
rect 6972 16504 6978 16516
rect 7469 16507 7527 16513
rect 7469 16504 7481 16507
rect 6972 16476 7481 16504
rect 6972 16464 6978 16476
rect 7469 16473 7481 16476
rect 7515 16504 7527 16507
rect 7558 16504 7564 16516
rect 7515 16476 7564 16504
rect 7515 16473 7527 16476
rect 7469 16467 7527 16473
rect 7558 16464 7564 16476
rect 7616 16464 7622 16516
rect 7653 16507 7711 16513
rect 7653 16473 7665 16507
rect 7699 16504 7711 16507
rect 9858 16504 9864 16516
rect 7699 16476 9864 16504
rect 7699 16473 7711 16476
rect 7653 16467 7711 16473
rect 9858 16464 9864 16476
rect 9916 16464 9922 16516
rect 10873 16507 10931 16513
rect 10873 16473 10885 16507
rect 10919 16504 10931 16507
rect 11606 16504 11612 16516
rect 10919 16476 11612 16504
rect 10919 16473 10931 16476
rect 10873 16467 10931 16473
rect 11606 16464 11612 16476
rect 11664 16464 11670 16516
rect 12406 16504 12434 16535
rect 13262 16532 13268 16544
rect 13320 16532 13326 16584
rect 13998 16532 14004 16584
rect 14056 16572 14062 16584
rect 14349 16575 14407 16581
rect 14349 16572 14361 16575
rect 14056 16544 14361 16572
rect 14056 16532 14062 16544
rect 14349 16541 14361 16544
rect 14395 16541 14407 16575
rect 16224 16572 16252 16600
rect 16761 16575 16819 16581
rect 16761 16572 16773 16575
rect 16224 16544 16773 16572
rect 14349 16535 14407 16541
rect 16761 16541 16773 16544
rect 16807 16541 16819 16575
rect 16761 16535 16819 16541
rect 16853 16575 16911 16581
rect 16853 16541 16865 16575
rect 16899 16541 16911 16575
rect 16853 16535 16911 16541
rect 16945 16575 17003 16581
rect 16945 16541 16957 16575
rect 16991 16569 17003 16575
rect 17034 16569 17040 16584
rect 16991 16541 17040 16569
rect 16945 16535 17003 16541
rect 13078 16504 13084 16516
rect 12406 16476 13084 16504
rect 13078 16464 13084 16476
rect 13136 16504 13142 16516
rect 13538 16504 13544 16516
rect 13136 16476 13544 16504
rect 13136 16464 13142 16476
rect 13538 16464 13544 16476
rect 13596 16464 13602 16516
rect 16868 16504 16896 16535
rect 17034 16532 17040 16541
rect 17092 16532 17098 16584
rect 17144 16581 17172 16612
rect 17310 16600 17316 16612
rect 17368 16640 17374 16652
rect 22646 16640 22652 16652
rect 17368 16612 22652 16640
rect 17368 16600 17374 16612
rect 17129 16575 17187 16581
rect 17129 16541 17141 16575
rect 17175 16541 17187 16575
rect 17129 16535 17187 16541
rect 18230 16532 18236 16584
rect 18288 16572 18294 16584
rect 18708 16581 18736 16612
rect 18325 16575 18383 16581
rect 18325 16572 18337 16575
rect 18288 16544 18337 16572
rect 18288 16532 18294 16544
rect 18325 16541 18337 16544
rect 18371 16541 18383 16575
rect 18325 16535 18383 16541
rect 18417 16575 18475 16581
rect 18417 16541 18429 16575
rect 18463 16541 18475 16575
rect 18417 16535 18475 16541
rect 18509 16575 18567 16581
rect 18509 16541 18521 16575
rect 18555 16541 18567 16575
rect 18509 16535 18567 16541
rect 18693 16575 18751 16581
rect 18693 16541 18705 16575
rect 18739 16541 18751 16575
rect 19610 16572 19616 16584
rect 19571 16544 19616 16572
rect 18693 16535 18751 16541
rect 17402 16504 17408 16516
rect 16868 16476 17408 16504
rect 17402 16464 17408 16476
rect 17460 16504 17466 16516
rect 18432 16504 18460 16535
rect 17460 16476 18460 16504
rect 18524 16504 18552 16535
rect 19610 16532 19616 16544
rect 19668 16532 19674 16584
rect 21468 16581 21496 16612
rect 22646 16600 22652 16612
rect 22704 16600 22710 16652
rect 25792 16649 25820 16748
rect 31018 16736 31024 16788
rect 31076 16776 31082 16788
rect 33226 16776 33232 16788
rect 31076 16748 33232 16776
rect 31076 16736 31082 16748
rect 33226 16736 33232 16748
rect 33284 16736 33290 16788
rect 34790 16776 34796 16788
rect 34703 16748 34796 16776
rect 34790 16736 34796 16748
rect 34848 16776 34854 16788
rect 37274 16776 37280 16788
rect 34848 16748 37280 16776
rect 34848 16736 34854 16748
rect 37274 16736 37280 16748
rect 37332 16736 37338 16788
rect 38102 16776 38108 16788
rect 38063 16748 38108 16776
rect 38102 16736 38108 16748
rect 38160 16736 38166 16788
rect 29546 16668 29552 16720
rect 29604 16668 29610 16720
rect 35253 16711 35311 16717
rect 35253 16677 35265 16711
rect 35299 16677 35311 16711
rect 37292 16708 37320 16736
rect 38378 16708 38384 16720
rect 37292 16680 38384 16708
rect 35253 16671 35311 16677
rect 25777 16643 25835 16649
rect 25777 16609 25789 16643
rect 25823 16640 25835 16643
rect 28537 16643 28595 16649
rect 28537 16640 28549 16643
rect 25823 16612 28549 16640
rect 25823 16609 25835 16612
rect 25777 16603 25835 16609
rect 28537 16609 28549 16612
rect 28583 16640 28595 16643
rect 28994 16640 29000 16652
rect 28583 16612 29000 16640
rect 28583 16609 28595 16612
rect 28537 16603 28595 16609
rect 28994 16600 29000 16612
rect 29052 16600 29058 16652
rect 29564 16640 29592 16668
rect 29825 16643 29883 16649
rect 29825 16640 29837 16643
rect 29564 16612 29837 16640
rect 29825 16609 29837 16612
rect 29871 16640 29883 16643
rect 30834 16640 30840 16652
rect 29871 16612 30840 16640
rect 29871 16609 29883 16612
rect 29825 16603 29883 16609
rect 30834 16600 30840 16612
rect 30892 16640 30898 16652
rect 30892 16612 31064 16640
rect 30892 16600 30898 16612
rect 21453 16575 21511 16581
rect 21453 16541 21465 16575
rect 21499 16541 21511 16575
rect 21616 16575 21674 16581
rect 21616 16572 21628 16575
rect 21453 16535 21511 16541
rect 21560 16544 21628 16572
rect 19245 16507 19303 16513
rect 19245 16504 19257 16507
rect 18524 16476 19257 16504
rect 17460 16464 17466 16476
rect 7006 16436 7012 16448
rect 5316 16408 6868 16436
rect 6967 16408 7012 16436
rect 5316 16396 5322 16408
rect 7006 16396 7012 16408
rect 7064 16396 7070 16448
rect 16485 16439 16543 16445
rect 16485 16405 16497 16439
rect 16531 16436 16543 16439
rect 16758 16436 16764 16448
rect 16531 16408 16764 16436
rect 16531 16405 16543 16408
rect 16485 16399 16543 16405
rect 16758 16396 16764 16408
rect 16816 16396 16822 16448
rect 18046 16436 18052 16448
rect 18007 16408 18052 16436
rect 18046 16396 18052 16408
rect 18104 16396 18110 16448
rect 18432 16436 18460 16476
rect 19245 16473 19257 16476
rect 19291 16473 19303 16507
rect 19426 16504 19432 16516
rect 19387 16476 19432 16504
rect 19245 16467 19303 16473
rect 19426 16464 19432 16476
rect 19484 16464 19490 16516
rect 21266 16464 21272 16516
rect 21324 16504 21330 16516
rect 21560 16504 21588 16544
rect 21616 16541 21628 16544
rect 21662 16541 21674 16575
rect 21616 16535 21674 16541
rect 21729 16575 21787 16581
rect 21729 16541 21741 16575
rect 21775 16541 21787 16575
rect 21729 16535 21787 16541
rect 21324 16476 21588 16504
rect 21324 16464 21330 16476
rect 21634 16436 21640 16448
rect 18432 16408 21640 16436
rect 21634 16396 21640 16408
rect 21692 16436 21698 16448
rect 21731 16436 21759 16535
rect 21818 16532 21824 16584
rect 21876 16572 21882 16584
rect 21876 16544 21921 16572
rect 21876 16532 21882 16544
rect 28166 16532 28172 16584
rect 28224 16572 28230 16584
rect 31036 16581 31064 16612
rect 32950 16600 32956 16652
rect 33008 16640 33014 16652
rect 33045 16643 33103 16649
rect 33045 16640 33057 16643
rect 33008 16612 33057 16640
rect 33008 16600 33014 16612
rect 33045 16609 33057 16612
rect 33091 16609 33103 16643
rect 33045 16603 33103 16609
rect 29549 16575 29607 16581
rect 29549 16572 29561 16575
rect 28224 16544 29561 16572
rect 28224 16532 28230 16544
rect 29549 16541 29561 16544
rect 29595 16541 29607 16575
rect 29549 16535 29607 16541
rect 31021 16575 31079 16581
rect 31021 16541 31033 16575
rect 31067 16541 31079 16575
rect 31021 16535 31079 16541
rect 31389 16575 31447 16581
rect 31389 16541 31401 16575
rect 31435 16572 31447 16575
rect 31570 16572 31576 16584
rect 31435 16544 31576 16572
rect 31435 16541 31447 16544
rect 31389 16535 31447 16541
rect 31570 16532 31576 16544
rect 31628 16532 31634 16584
rect 32769 16575 32827 16581
rect 32769 16541 32781 16575
rect 32815 16572 32827 16575
rect 32858 16572 32864 16584
rect 32815 16544 32864 16572
rect 32815 16541 32827 16544
rect 32769 16535 32827 16541
rect 32858 16532 32864 16544
rect 32916 16532 32922 16584
rect 33410 16532 33416 16584
rect 33468 16572 33474 16584
rect 33689 16575 33747 16581
rect 33689 16572 33701 16575
rect 33468 16544 33701 16572
rect 33468 16532 33474 16544
rect 33689 16541 33701 16544
rect 33735 16572 33747 16575
rect 35268 16572 35296 16671
rect 38378 16668 38384 16680
rect 38436 16668 38442 16720
rect 36630 16640 36636 16652
rect 36591 16612 36636 16640
rect 36630 16600 36636 16612
rect 36688 16600 36694 16652
rect 33735 16544 35296 16572
rect 33735 16541 33747 16544
rect 33689 16535 33747 16541
rect 25532 16507 25590 16513
rect 25532 16473 25544 16507
rect 25578 16504 25590 16507
rect 25774 16504 25780 16516
rect 25578 16476 25780 16504
rect 25578 16473 25590 16476
rect 25532 16467 25590 16473
rect 25774 16464 25780 16476
rect 25832 16464 25838 16516
rect 26789 16507 26847 16513
rect 26789 16473 26801 16507
rect 26835 16504 26847 16507
rect 28902 16504 28908 16516
rect 26835 16476 28908 16504
rect 26835 16473 26847 16476
rect 26789 16467 26847 16473
rect 28902 16464 28908 16476
rect 28960 16464 28966 16516
rect 31110 16504 31116 16516
rect 31071 16476 31116 16504
rect 31110 16464 31116 16476
rect 31168 16464 31174 16516
rect 31202 16464 31208 16516
rect 31260 16504 31266 16516
rect 31260 16476 31305 16504
rect 31260 16464 31266 16476
rect 32122 16464 32128 16516
rect 32180 16504 32186 16516
rect 33505 16507 33563 16513
rect 33505 16504 33517 16507
rect 32180 16476 33517 16504
rect 32180 16464 32186 16476
rect 33505 16473 33517 16476
rect 33551 16473 33563 16507
rect 33505 16467 33563 16473
rect 34514 16464 34520 16516
rect 34572 16504 34578 16516
rect 36366 16507 36424 16513
rect 36366 16504 36378 16507
rect 34572 16476 36378 16504
rect 34572 16464 34578 16476
rect 36366 16473 36378 16476
rect 36412 16473 36424 16507
rect 37734 16504 37740 16516
rect 37695 16476 37740 16504
rect 36366 16467 36424 16473
rect 37734 16464 37740 16476
rect 37792 16464 37798 16516
rect 37826 16464 37832 16516
rect 37884 16504 37890 16516
rect 37921 16507 37979 16513
rect 37921 16504 37933 16507
rect 37884 16476 37933 16504
rect 37884 16464 37890 16476
rect 37921 16473 37933 16476
rect 37967 16504 37979 16507
rect 40586 16504 40592 16516
rect 37967 16476 40592 16504
rect 37967 16473 37979 16476
rect 37921 16467 37979 16473
rect 40586 16464 40592 16476
rect 40644 16464 40650 16516
rect 21692 16408 21759 16436
rect 21692 16396 21698 16408
rect 24302 16396 24308 16448
rect 24360 16436 24366 16448
rect 24397 16439 24455 16445
rect 24397 16436 24409 16439
rect 24360 16408 24409 16436
rect 24360 16396 24366 16408
rect 24397 16405 24409 16408
rect 24443 16405 24455 16439
rect 26326 16436 26332 16448
rect 26287 16408 26332 16436
rect 24397 16399 24455 16405
rect 26326 16396 26332 16408
rect 26384 16396 26390 16448
rect 27338 16396 27344 16448
rect 27396 16436 27402 16448
rect 30837 16439 30895 16445
rect 30837 16436 30849 16439
rect 27396 16408 30849 16436
rect 27396 16396 27402 16408
rect 30837 16405 30849 16408
rect 30883 16405 30895 16439
rect 30837 16399 30895 16405
rect 31478 16396 31484 16448
rect 31536 16436 31542 16448
rect 32582 16436 32588 16448
rect 31536 16408 32588 16436
rect 31536 16396 31542 16408
rect 32582 16396 32588 16408
rect 32640 16396 32646 16448
rect 33873 16439 33931 16445
rect 33873 16405 33885 16439
rect 33919 16436 33931 16439
rect 34054 16436 34060 16448
rect 33919 16408 34060 16436
rect 33919 16405 33931 16408
rect 33873 16399 33931 16405
rect 34054 16396 34060 16408
rect 34112 16396 34118 16448
rect 1104 16346 68816 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 68816 16346
rect 1104 16272 68816 16294
rect 6822 16192 6828 16244
rect 6880 16232 6886 16244
rect 8665 16235 8723 16241
rect 8665 16232 8677 16235
rect 6880 16204 8677 16232
rect 6880 16192 6886 16204
rect 8665 16201 8677 16204
rect 8711 16232 8723 16235
rect 11330 16232 11336 16244
rect 8711 16204 11336 16232
rect 8711 16201 8723 16204
rect 8665 16195 8723 16201
rect 11330 16192 11336 16204
rect 11388 16192 11394 16244
rect 14366 16232 14372 16244
rect 14327 16204 14372 16232
rect 14366 16192 14372 16204
rect 14424 16192 14430 16244
rect 17034 16232 17040 16244
rect 16995 16204 17040 16232
rect 17034 16192 17040 16204
rect 17092 16192 17098 16244
rect 17957 16235 18015 16241
rect 17957 16201 17969 16235
rect 18003 16232 18015 16235
rect 18230 16232 18236 16244
rect 18003 16204 18236 16232
rect 18003 16201 18015 16204
rect 17957 16195 18015 16201
rect 18230 16192 18236 16204
rect 18288 16192 18294 16244
rect 21818 16232 21824 16244
rect 21779 16204 21824 16232
rect 21818 16192 21824 16204
rect 21876 16192 21882 16244
rect 23106 16192 23112 16244
rect 23164 16232 23170 16244
rect 23201 16235 23259 16241
rect 23201 16232 23213 16235
rect 23164 16204 23213 16232
rect 23164 16192 23170 16204
rect 23201 16201 23213 16204
rect 23247 16232 23259 16235
rect 25774 16232 25780 16244
rect 23247 16204 23888 16232
rect 25735 16204 25780 16232
rect 23247 16201 23259 16204
rect 23201 16195 23259 16201
rect 5166 16164 5172 16176
rect 5127 16136 5172 16164
rect 5166 16124 5172 16136
rect 5224 16124 5230 16176
rect 7377 16167 7435 16173
rect 6380 16136 6960 16164
rect 2038 16096 2044 16108
rect 1951 16068 2044 16096
rect 2038 16056 2044 16068
rect 2096 16056 2102 16108
rect 2222 16096 2228 16108
rect 2183 16068 2228 16096
rect 2222 16056 2228 16068
rect 2280 16056 2286 16108
rect 2314 16056 2320 16108
rect 2372 16096 2378 16108
rect 2455 16099 2513 16105
rect 2372 16068 2417 16096
rect 2372 16056 2378 16068
rect 2455 16065 2467 16099
rect 2501 16096 2513 16099
rect 2682 16096 2688 16108
rect 2501 16068 2688 16096
rect 2501 16065 2513 16068
rect 2455 16059 2513 16065
rect 2682 16056 2688 16068
rect 2740 16096 2746 16108
rect 3145 16099 3203 16105
rect 3145 16096 3157 16099
rect 2740 16068 3157 16096
rect 2740 16056 2746 16068
rect 3145 16065 3157 16068
rect 3191 16065 3203 16099
rect 3145 16059 3203 16065
rect 4893 16099 4951 16105
rect 4893 16065 4905 16099
rect 4939 16096 4951 16099
rect 4982 16096 4988 16108
rect 4939 16068 4988 16096
rect 4939 16065 4951 16068
rect 4893 16059 4951 16065
rect 4982 16056 4988 16068
rect 5040 16056 5046 16108
rect 6380 16105 6408 16136
rect 5077 16099 5135 16105
rect 5077 16065 5089 16099
rect 5123 16096 5135 16099
rect 5261 16099 5319 16105
rect 5123 16068 5212 16096
rect 5123 16065 5135 16068
rect 5077 16059 5135 16065
rect 2056 16028 2084 16056
rect 2056 16000 4936 16028
rect 4908 15972 4936 16000
rect 4890 15920 4896 15972
rect 4948 15920 4954 15972
rect 5184 15960 5212 16068
rect 5261 16065 5273 16099
rect 5307 16065 5319 16099
rect 5261 16059 5319 16065
rect 6365 16099 6423 16105
rect 6365 16065 6377 16099
rect 6411 16065 6423 16099
rect 6546 16096 6552 16108
rect 6507 16068 6552 16096
rect 6365 16059 6423 16065
rect 5276 16028 5304 16059
rect 6546 16056 6552 16068
rect 6604 16056 6610 16108
rect 6564 16028 6592 16056
rect 6932 16028 6960 16136
rect 7377 16133 7389 16167
rect 7423 16164 7435 16167
rect 10318 16164 10324 16176
rect 7423 16136 10324 16164
rect 7423 16133 7435 16136
rect 7377 16127 7435 16133
rect 10318 16124 10324 16136
rect 10376 16124 10382 16176
rect 12805 16167 12863 16173
rect 12805 16133 12817 16167
rect 12851 16164 12863 16167
rect 13906 16164 13912 16176
rect 12851 16136 13912 16164
rect 12851 16133 12863 16136
rect 12805 16127 12863 16133
rect 13906 16124 13912 16136
rect 13964 16164 13970 16176
rect 15289 16167 15347 16173
rect 15289 16164 15301 16167
rect 13964 16136 15301 16164
rect 13964 16124 13970 16136
rect 15289 16133 15301 16136
rect 15335 16133 15347 16167
rect 16666 16164 16672 16176
rect 16627 16136 16672 16164
rect 15289 16127 15347 16133
rect 16666 16124 16672 16136
rect 16724 16124 16730 16176
rect 19426 16124 19432 16176
rect 19484 16164 19490 16176
rect 19484 16136 19748 16164
rect 19484 16124 19490 16136
rect 19720 16108 19748 16136
rect 19794 16124 19800 16176
rect 19852 16164 19858 16176
rect 23860 16173 23888 16204
rect 25774 16192 25780 16204
rect 25832 16192 25838 16244
rect 25884 16204 26464 16232
rect 19889 16167 19947 16173
rect 19889 16164 19901 16167
rect 19852 16136 19901 16164
rect 19852 16124 19858 16136
rect 19889 16133 19901 16136
rect 19935 16133 19947 16167
rect 19889 16127 19947 16133
rect 19981 16167 20039 16173
rect 19981 16133 19993 16167
rect 20027 16164 20039 16167
rect 23845 16167 23903 16173
rect 20027 16136 22968 16164
rect 20027 16133 20039 16136
rect 19981 16127 20039 16133
rect 22940 16108 22968 16136
rect 23845 16133 23857 16167
rect 23891 16133 23903 16167
rect 23845 16127 23903 16133
rect 24029 16167 24087 16173
rect 24029 16133 24041 16167
rect 24075 16164 24087 16167
rect 24857 16167 24915 16173
rect 24075 16136 24808 16164
rect 24075 16133 24087 16136
rect 24029 16127 24087 16133
rect 7558 16096 7564 16108
rect 7519 16068 7564 16096
rect 7558 16056 7564 16068
rect 7616 16056 7622 16108
rect 12434 16056 12440 16108
rect 12492 16096 12498 16108
rect 12618 16096 12624 16108
rect 12492 16068 12624 16096
rect 12492 16056 12498 16068
rect 12618 16056 12624 16068
rect 12676 16056 12682 16108
rect 15010 16096 15016 16108
rect 14971 16068 15016 16096
rect 15010 16056 15016 16068
rect 15068 16056 15074 16108
rect 15197 16099 15255 16105
rect 15197 16065 15209 16099
rect 15243 16065 15255 16099
rect 15197 16059 15255 16065
rect 15381 16099 15439 16105
rect 15381 16065 15393 16099
rect 15427 16065 15439 16099
rect 15381 16059 15439 16065
rect 16853 16099 16911 16105
rect 16853 16065 16865 16099
rect 16899 16096 16911 16099
rect 17954 16096 17960 16108
rect 16899 16068 17960 16096
rect 16899 16065 16911 16068
rect 16853 16059 16911 16065
rect 7006 16028 7012 16040
rect 5276 16000 6592 16028
rect 6919 16000 7012 16028
rect 7006 15988 7012 16000
rect 7064 16028 7070 16040
rect 7742 16028 7748 16040
rect 7064 16000 7748 16028
rect 7064 15988 7070 16000
rect 7742 15988 7748 16000
rect 7800 15988 7806 16040
rect 5258 15960 5264 15972
rect 5184 15932 5264 15960
rect 5258 15920 5264 15932
rect 5316 15920 5322 15972
rect 5442 15960 5448 15972
rect 5403 15932 5448 15960
rect 5442 15920 5448 15932
rect 5500 15920 5506 15972
rect 6362 15920 6368 15972
rect 6420 15960 6426 15972
rect 7558 15960 7564 15972
rect 6420 15932 7564 15960
rect 6420 15920 6426 15932
rect 7558 15920 7564 15932
rect 7616 15960 7622 15972
rect 8021 15963 8079 15969
rect 8021 15960 8033 15963
rect 7616 15932 8033 15960
rect 7616 15920 7622 15932
rect 8021 15929 8033 15932
rect 8067 15929 8079 15963
rect 15212 15960 15240 16059
rect 15286 15988 15292 16040
rect 15344 16028 15350 16040
rect 15396 16028 15424 16059
rect 17954 16056 17960 16068
rect 18012 16056 18018 16108
rect 18690 16056 18696 16108
rect 18748 16096 18754 16108
rect 19613 16099 19671 16105
rect 19613 16096 19625 16099
rect 18748 16068 19625 16096
rect 18748 16056 18754 16068
rect 19613 16065 19625 16068
rect 19659 16065 19671 16099
rect 19613 16059 19671 16065
rect 19702 16056 19708 16108
rect 19760 16096 19766 16108
rect 19760 16068 19805 16096
rect 19760 16056 19766 16068
rect 20070 16056 20076 16108
rect 20128 16105 20134 16108
rect 20128 16096 20136 16105
rect 21269 16099 21327 16105
rect 20128 16068 20173 16096
rect 20128 16059 20136 16068
rect 21269 16065 21281 16099
rect 21315 16096 21327 16099
rect 21315 16068 22094 16096
rect 21315 16065 21327 16068
rect 21269 16059 21327 16065
rect 20128 16056 20134 16059
rect 15746 16028 15752 16040
rect 15344 16000 15424 16028
rect 15488 16000 15752 16028
rect 15344 15988 15350 16000
rect 15378 15960 15384 15972
rect 15212 15932 15384 15960
rect 8021 15923 8079 15929
rect 15378 15920 15384 15932
rect 15436 15960 15442 15972
rect 15488 15960 15516 16000
rect 15746 15988 15752 16000
rect 15804 15988 15810 16040
rect 16390 15988 16396 16040
rect 16448 16028 16454 16040
rect 20254 16028 20260 16040
rect 16448 16000 20260 16028
rect 16448 15988 16454 16000
rect 20254 15988 20260 16000
rect 20312 15988 20318 16040
rect 21177 16031 21235 16037
rect 21177 15997 21189 16031
rect 21223 16028 21235 16031
rect 21818 16028 21824 16040
rect 21223 16000 21824 16028
rect 21223 15997 21235 16000
rect 21177 15991 21235 15997
rect 21818 15988 21824 16000
rect 21876 15988 21882 16040
rect 22066 16028 22094 16068
rect 22922 16056 22928 16108
rect 22980 16096 22986 16108
rect 24673 16099 24731 16105
rect 24673 16096 24685 16099
rect 22980 16068 24685 16096
rect 22980 16056 22986 16068
rect 24673 16065 24685 16068
rect 24719 16065 24731 16099
rect 24780 16096 24808 16136
rect 24857 16133 24869 16167
rect 24903 16164 24915 16167
rect 25130 16164 25136 16176
rect 24903 16136 25136 16164
rect 24903 16133 24915 16136
rect 24857 16127 24915 16133
rect 25130 16124 25136 16136
rect 25188 16124 25194 16176
rect 25314 16124 25320 16176
rect 25372 16164 25378 16176
rect 25884 16164 25912 16204
rect 26326 16164 26332 16176
rect 25372 16136 25912 16164
rect 26068 16136 26332 16164
rect 25372 16124 25378 16136
rect 25958 16096 25964 16108
rect 24780 16068 25964 16096
rect 24673 16059 24731 16065
rect 25958 16056 25964 16068
rect 26016 16096 26022 16108
rect 26068 16105 26096 16136
rect 26326 16124 26332 16136
rect 26384 16124 26390 16176
rect 26053 16099 26111 16105
rect 26053 16096 26065 16099
rect 26016 16068 26065 16096
rect 26016 16056 26022 16068
rect 26053 16065 26065 16068
rect 26099 16065 26111 16099
rect 26053 16059 26111 16065
rect 26145 16099 26203 16105
rect 26145 16065 26157 16099
rect 26191 16065 26203 16099
rect 26145 16059 26203 16065
rect 24854 16028 24860 16040
rect 22066 16000 24860 16028
rect 24854 15988 24860 16000
rect 24912 15988 24918 16040
rect 25774 15988 25780 16040
rect 25832 16028 25838 16040
rect 26160 16028 26188 16059
rect 26234 16056 26240 16108
rect 26292 16096 26298 16108
rect 26436 16105 26464 16204
rect 28902 16192 28908 16244
rect 28960 16232 28966 16244
rect 29914 16232 29920 16244
rect 28960 16204 29920 16232
rect 28960 16192 28966 16204
rect 29914 16192 29920 16204
rect 29972 16192 29978 16244
rect 32953 16235 33011 16241
rect 32953 16201 32965 16235
rect 32999 16232 33011 16235
rect 33134 16232 33140 16244
rect 32999 16204 33140 16232
rect 32999 16201 33011 16204
rect 32953 16195 33011 16201
rect 33134 16192 33140 16204
rect 33192 16192 33198 16244
rect 34514 16232 34520 16244
rect 34475 16204 34520 16232
rect 34514 16192 34520 16204
rect 34572 16192 34578 16244
rect 35897 16235 35955 16241
rect 35897 16201 35909 16235
rect 35943 16232 35955 16235
rect 37734 16232 37740 16244
rect 35943 16204 37740 16232
rect 35943 16201 35955 16204
rect 35897 16195 35955 16201
rect 37734 16192 37740 16204
rect 37792 16192 37798 16244
rect 28626 16164 28632 16176
rect 28587 16136 28632 16164
rect 28626 16124 28632 16136
rect 28684 16124 28690 16176
rect 31113 16167 31171 16173
rect 31113 16133 31125 16167
rect 31159 16164 31171 16167
rect 31159 16136 32168 16164
rect 31159 16133 31171 16136
rect 31113 16127 31171 16133
rect 26421 16099 26479 16105
rect 26292 16068 26337 16096
rect 26292 16056 26298 16068
rect 26421 16065 26433 16099
rect 26467 16096 26479 16099
rect 26786 16096 26792 16108
rect 26467 16068 26792 16096
rect 26467 16065 26479 16068
rect 26421 16059 26479 16065
rect 26786 16056 26792 16068
rect 26844 16056 26850 16108
rect 27893 16099 27951 16105
rect 27893 16065 27905 16099
rect 27939 16096 27951 16099
rect 28810 16096 28816 16108
rect 27939 16068 28816 16096
rect 27939 16065 27951 16068
rect 27893 16059 27951 16065
rect 28810 16056 28816 16068
rect 28868 16056 28874 16108
rect 30834 16056 30840 16108
rect 30892 16096 30898 16108
rect 31021 16099 31079 16105
rect 31021 16096 31033 16099
rect 30892 16068 31033 16096
rect 30892 16056 30898 16068
rect 31021 16065 31033 16068
rect 31067 16065 31079 16099
rect 31021 16059 31079 16065
rect 31202 16056 31208 16108
rect 31260 16096 31266 16108
rect 31389 16099 31447 16105
rect 31260 16068 31353 16096
rect 31260 16056 31266 16068
rect 31389 16065 31401 16099
rect 31435 16096 31447 16099
rect 31662 16096 31668 16108
rect 31435 16068 31668 16096
rect 31435 16065 31447 16068
rect 31389 16059 31447 16065
rect 31662 16056 31668 16068
rect 31720 16056 31726 16108
rect 27706 16028 27712 16040
rect 25832 16000 27712 16028
rect 25832 15988 25838 16000
rect 27706 15988 27712 16000
rect 27764 15988 27770 16040
rect 28169 16031 28227 16037
rect 28169 15997 28181 16031
rect 28215 16028 28227 16031
rect 28534 16028 28540 16040
rect 28215 16000 28540 16028
rect 28215 15997 28227 16000
rect 28169 15991 28227 15997
rect 28534 15988 28540 16000
rect 28592 15988 28598 16040
rect 28828 16028 28856 16056
rect 31220 16028 31248 16056
rect 28828 16000 31248 16028
rect 15436 15932 15516 15960
rect 15565 15963 15623 15969
rect 15436 15920 15442 15932
rect 15565 15929 15577 15963
rect 15611 15960 15623 15963
rect 19426 15960 19432 15972
rect 15611 15932 19432 15960
rect 15611 15929 15623 15932
rect 15565 15923 15623 15929
rect 19426 15920 19432 15932
rect 19484 15920 19490 15972
rect 20346 15920 20352 15972
rect 20404 15960 20410 15972
rect 32140 15960 32168 16136
rect 32858 16124 32864 16176
rect 32916 16164 32922 16176
rect 37642 16164 37648 16176
rect 32916 16136 34192 16164
rect 32916 16124 32922 16136
rect 32306 16096 32312 16108
rect 32267 16068 32312 16096
rect 32306 16056 32312 16068
rect 32364 16056 32370 16108
rect 32490 16096 32496 16108
rect 32451 16068 32496 16096
rect 32490 16056 32496 16068
rect 32548 16056 32554 16108
rect 32585 16099 32643 16105
rect 32585 16065 32597 16099
rect 32631 16065 32643 16099
rect 32585 16059 32643 16065
rect 32600 16028 32628 16059
rect 32674 16056 32680 16108
rect 32732 16096 32738 16108
rect 32732 16068 32777 16096
rect 32732 16056 32738 16068
rect 33594 16056 33600 16108
rect 33652 16096 33658 16108
rect 33873 16099 33931 16105
rect 33873 16096 33885 16099
rect 33652 16068 33885 16096
rect 33652 16056 33658 16068
rect 33873 16065 33885 16068
rect 33919 16065 33931 16099
rect 34054 16096 34060 16108
rect 34015 16068 34060 16096
rect 33873 16059 33931 16065
rect 34054 16056 34060 16068
rect 34112 16056 34118 16108
rect 34164 16105 34192 16136
rect 35636 16136 37648 16164
rect 34149 16099 34207 16105
rect 34149 16065 34161 16099
rect 34195 16065 34207 16099
rect 34149 16059 34207 16065
rect 34241 16099 34299 16105
rect 34241 16065 34253 16099
rect 34287 16065 34299 16099
rect 34241 16059 34299 16065
rect 32950 16028 32956 16040
rect 32600 16000 32956 16028
rect 32950 15988 32956 16000
rect 33008 15988 33014 16040
rect 33686 15988 33692 16040
rect 33744 16028 33750 16040
rect 34256 16028 34284 16059
rect 33744 16000 34284 16028
rect 33744 15988 33750 16000
rect 35636 15960 35664 16136
rect 37642 16124 37648 16136
rect 37700 16124 37706 16176
rect 38381 16167 38439 16173
rect 37939 16136 38332 16164
rect 35713 16099 35771 16105
rect 35713 16065 35725 16099
rect 35759 16065 35771 16099
rect 35713 16059 35771 16065
rect 20404 15932 21128 15960
rect 32140 15932 35664 15960
rect 20404 15920 20410 15932
rect 2682 15892 2688 15904
rect 2643 15864 2688 15892
rect 2682 15852 2688 15864
rect 2740 15852 2746 15904
rect 6454 15892 6460 15904
rect 6415 15864 6460 15892
rect 6454 15852 6460 15864
rect 6512 15852 6518 15904
rect 7190 15892 7196 15904
rect 7151 15864 7196 15892
rect 7190 15852 7196 15864
rect 7248 15852 7254 15904
rect 12158 15892 12164 15904
rect 12119 15864 12164 15892
rect 12158 15852 12164 15864
rect 12216 15852 12222 15904
rect 12989 15895 13047 15901
rect 12989 15861 13001 15895
rect 13035 15892 13047 15895
rect 13078 15892 13084 15904
rect 13035 15864 13084 15892
rect 13035 15861 13047 15864
rect 12989 15855 13047 15861
rect 13078 15852 13084 15864
rect 13136 15852 13142 15904
rect 13538 15892 13544 15904
rect 13499 15864 13544 15892
rect 13538 15852 13544 15864
rect 13596 15852 13602 15904
rect 20257 15895 20315 15901
rect 20257 15861 20269 15895
rect 20303 15892 20315 15895
rect 20438 15892 20444 15904
rect 20303 15864 20444 15892
rect 20303 15861 20315 15864
rect 20257 15855 20315 15861
rect 20438 15852 20444 15864
rect 20496 15852 20502 15904
rect 20898 15892 20904 15904
rect 20859 15864 20904 15892
rect 20898 15852 20904 15864
rect 20956 15852 20962 15904
rect 21100 15901 21128 15932
rect 21085 15895 21143 15901
rect 21085 15861 21097 15895
rect 21131 15861 21143 15895
rect 21085 15855 21143 15861
rect 24489 15895 24547 15901
rect 24489 15861 24501 15895
rect 24535 15892 24547 15895
rect 25498 15892 25504 15904
rect 24535 15864 25504 15892
rect 24535 15861 24547 15864
rect 24489 15855 24547 15861
rect 25498 15852 25504 15864
rect 25556 15852 25562 15904
rect 25590 15852 25596 15904
rect 25648 15892 25654 15904
rect 30837 15895 30895 15901
rect 30837 15892 30849 15895
rect 25648 15864 30849 15892
rect 25648 15852 25654 15864
rect 30837 15861 30849 15864
rect 30883 15861 30895 15895
rect 30837 15855 30895 15861
rect 31386 15852 31392 15904
rect 31444 15892 31450 15904
rect 35728 15892 35756 16059
rect 37458 16056 37464 16108
rect 37516 16096 37522 16108
rect 37939 16105 37967 16136
rect 37737 16099 37795 16105
rect 37737 16096 37749 16099
rect 37516 16068 37749 16096
rect 37516 16056 37522 16068
rect 37737 16065 37749 16068
rect 37783 16065 37795 16099
rect 37737 16059 37795 16065
rect 37900 16099 37967 16105
rect 37900 16065 37912 16099
rect 37946 16068 37967 16099
rect 38000 16099 38058 16105
rect 37946 16065 37958 16068
rect 37900 16059 37958 16065
rect 38000 16065 38012 16099
rect 38046 16065 38058 16099
rect 38000 16059 38058 16065
rect 38105 16099 38163 16105
rect 38105 16065 38117 16099
rect 38151 16096 38163 16099
rect 38194 16096 38200 16108
rect 38151 16068 38200 16096
rect 38151 16065 38163 16068
rect 38105 16059 38163 16065
rect 37642 15988 37648 16040
rect 37700 16028 37706 16040
rect 38015 16028 38043 16059
rect 37700 16000 38043 16028
rect 37700 15988 37706 16000
rect 38120 15960 38148 16059
rect 38194 16056 38200 16068
rect 38252 16056 38258 16108
rect 38304 16096 38332 16136
rect 38381 16133 38393 16167
rect 38427 16164 38439 16167
rect 40322 16167 40380 16173
rect 40322 16164 40334 16167
rect 38427 16136 40334 16164
rect 38427 16133 38439 16136
rect 38381 16127 38439 16133
rect 40322 16133 40334 16136
rect 40368 16133 40380 16167
rect 40322 16127 40380 16133
rect 38838 16096 38844 16108
rect 38304 16068 38844 16096
rect 38838 16056 38844 16068
rect 38896 16056 38902 16108
rect 40589 16031 40647 16037
rect 40589 15997 40601 16031
rect 40635 16028 40647 16031
rect 41230 16028 41236 16040
rect 40635 16000 41236 16028
rect 40635 15997 40647 16000
rect 40589 15991 40647 15997
rect 41230 15988 41236 16000
rect 41288 15988 41294 16040
rect 36648 15932 38148 15960
rect 31444 15864 35756 15892
rect 31444 15852 31450 15864
rect 36538 15852 36544 15904
rect 36596 15892 36602 15904
rect 36648 15901 36676 15932
rect 36633 15895 36691 15901
rect 36633 15892 36645 15895
rect 36596 15864 36645 15892
rect 36596 15852 36602 15864
rect 36633 15861 36645 15864
rect 36679 15861 36691 15895
rect 36633 15855 36691 15861
rect 38654 15852 38660 15904
rect 38712 15892 38718 15904
rect 39209 15895 39267 15901
rect 39209 15892 39221 15895
rect 38712 15864 39221 15892
rect 38712 15852 38718 15864
rect 39209 15861 39221 15864
rect 39255 15861 39267 15895
rect 67634 15892 67640 15904
rect 67595 15864 67640 15892
rect 39209 15855 39267 15861
rect 67634 15852 67640 15864
rect 67692 15852 67698 15904
rect 1104 15802 68816 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 65654 15802
rect 65706 15750 65718 15802
rect 65770 15750 65782 15802
rect 65834 15750 65846 15802
rect 65898 15750 65910 15802
rect 65962 15750 68816 15802
rect 1104 15728 68816 15750
rect 2222 15688 2228 15700
rect 2183 15660 2228 15688
rect 2222 15648 2228 15660
rect 2280 15648 2286 15700
rect 6914 15648 6920 15700
rect 6972 15688 6978 15700
rect 7101 15691 7159 15697
rect 7101 15688 7113 15691
rect 6972 15660 7113 15688
rect 6972 15648 6978 15660
rect 7101 15657 7113 15660
rect 7147 15657 7159 15691
rect 7101 15651 7159 15657
rect 10873 15691 10931 15697
rect 10873 15657 10885 15691
rect 10919 15688 10931 15691
rect 11330 15688 11336 15700
rect 10919 15660 11336 15688
rect 10919 15657 10931 15660
rect 10873 15651 10931 15657
rect 11330 15648 11336 15660
rect 11388 15648 11394 15700
rect 15654 15648 15660 15700
rect 15712 15688 15718 15700
rect 15749 15691 15807 15697
rect 15749 15688 15761 15691
rect 15712 15660 15761 15688
rect 15712 15648 15718 15660
rect 15749 15657 15761 15660
rect 15795 15657 15807 15691
rect 15749 15651 15807 15657
rect 18693 15691 18751 15697
rect 18693 15657 18705 15691
rect 18739 15688 18751 15691
rect 19702 15688 19708 15700
rect 18739 15660 19708 15688
rect 18739 15657 18751 15660
rect 18693 15651 18751 15657
rect 19702 15648 19708 15660
rect 19760 15648 19766 15700
rect 19794 15648 19800 15700
rect 19852 15688 19858 15700
rect 20806 15697 20812 15700
rect 20763 15691 20812 15697
rect 20763 15688 20775 15691
rect 19852 15660 20775 15688
rect 19852 15648 19858 15660
rect 20763 15657 20775 15660
rect 20809 15657 20812 15691
rect 20763 15651 20812 15657
rect 20806 15648 20812 15651
rect 20864 15688 20870 15700
rect 21818 15688 21824 15700
rect 20864 15660 20911 15688
rect 21779 15660 21824 15688
rect 20864 15648 20870 15660
rect 21818 15648 21824 15660
rect 21876 15648 21882 15700
rect 22281 15691 22339 15697
rect 22281 15657 22293 15691
rect 22327 15688 22339 15691
rect 25590 15688 25596 15700
rect 22327 15660 25596 15688
rect 22327 15657 22339 15660
rect 22281 15651 22339 15657
rect 25590 15648 25596 15660
rect 25648 15648 25654 15700
rect 25869 15691 25927 15697
rect 25869 15657 25881 15691
rect 25915 15657 25927 15691
rect 27338 15688 27344 15700
rect 27299 15660 27344 15688
rect 25869 15651 25927 15657
rect 7006 15620 7012 15632
rect 6196 15592 7012 15620
rect 2682 15512 2688 15564
rect 2740 15552 2746 15564
rect 6196 15561 6224 15592
rect 7006 15580 7012 15592
rect 7064 15580 7070 15632
rect 10778 15580 10784 15632
rect 10836 15620 10842 15632
rect 10836 15592 15976 15620
rect 10836 15580 10842 15592
rect 6181 15555 6239 15561
rect 2740 15524 3924 15552
rect 2740 15512 2746 15524
rect 1854 15484 1860 15496
rect 1815 15456 1860 15484
rect 1854 15444 1860 15456
rect 1912 15444 1918 15496
rect 3142 15444 3148 15496
rect 3200 15484 3206 15496
rect 3786 15484 3792 15496
rect 3200 15456 3792 15484
rect 3200 15444 3206 15456
rect 3786 15444 3792 15456
rect 3844 15444 3850 15496
rect 3896 15484 3924 15524
rect 6181 15521 6193 15555
rect 6227 15521 6239 15555
rect 6181 15515 6239 15521
rect 6362 15512 6368 15564
rect 6420 15552 6426 15564
rect 6457 15555 6515 15561
rect 6457 15552 6469 15555
rect 6420 15524 6469 15552
rect 6420 15512 6426 15524
rect 6457 15521 6469 15524
rect 6503 15521 6515 15555
rect 6457 15515 6515 15521
rect 7561 15555 7619 15561
rect 7561 15521 7573 15555
rect 7607 15552 7619 15555
rect 8018 15552 8024 15564
rect 7607 15524 8024 15552
rect 7607 15521 7619 15524
rect 7561 15515 7619 15521
rect 8018 15512 8024 15524
rect 8076 15552 8082 15564
rect 9033 15555 9091 15561
rect 9033 15552 9045 15555
rect 8076 15524 9045 15552
rect 8076 15512 8082 15524
rect 9033 15521 9045 15524
rect 9079 15521 9091 15555
rect 9033 15515 9091 15521
rect 12710 15512 12716 15564
rect 12768 15552 12774 15564
rect 12768 15524 13032 15552
rect 12768 15512 12774 15524
rect 4045 15487 4103 15493
rect 4045 15484 4057 15487
rect 3896 15456 4057 15484
rect 4045 15453 4057 15456
rect 4091 15453 4103 15487
rect 4045 15447 4103 15453
rect 6917 15487 6975 15493
rect 6917 15453 6929 15487
rect 6963 15484 6975 15487
rect 7282 15484 7288 15496
rect 6963 15456 7288 15484
rect 6963 15453 6975 15456
rect 6917 15447 6975 15453
rect 7282 15444 7288 15456
rect 7340 15444 7346 15496
rect 7834 15484 7840 15496
rect 7795 15456 7840 15484
rect 7834 15444 7840 15456
rect 7892 15444 7898 15496
rect 8941 15487 8999 15493
rect 8941 15453 8953 15487
rect 8987 15453 8999 15487
rect 8941 15447 8999 15453
rect 9125 15487 9183 15493
rect 9125 15453 9137 15487
rect 9171 15484 9183 15487
rect 9674 15484 9680 15496
rect 9171 15456 9680 15484
rect 9171 15453 9183 15456
rect 9125 15447 9183 15453
rect 2041 15419 2099 15425
rect 2041 15385 2053 15419
rect 2087 15416 2099 15419
rect 5074 15416 5080 15428
rect 2087 15388 5080 15416
rect 2087 15385 2099 15388
rect 2041 15379 2099 15385
rect 5074 15376 5080 15388
rect 5132 15416 5138 15428
rect 5132 15388 5212 15416
rect 5132 15376 5138 15388
rect 5184 15357 5212 15388
rect 7742 15376 7748 15428
rect 7800 15416 7806 15428
rect 8956 15416 8984 15447
rect 7800 15388 8984 15416
rect 7800 15376 7806 15388
rect 5169 15351 5227 15357
rect 5169 15317 5181 15351
rect 5215 15317 5227 15351
rect 5169 15311 5227 15317
rect 5258 15308 5264 15360
rect 5316 15348 5322 15360
rect 6270 15348 6276 15360
rect 5316 15320 6276 15348
rect 5316 15308 5322 15320
rect 6270 15308 6276 15320
rect 6328 15348 6334 15360
rect 6914 15348 6920 15360
rect 6328 15320 6920 15348
rect 6328 15308 6334 15320
rect 6914 15308 6920 15320
rect 6972 15348 6978 15360
rect 9140 15348 9168 15447
rect 9674 15444 9680 15456
rect 9732 15444 9738 15496
rect 12158 15484 12164 15496
rect 12119 15456 12164 15484
rect 12158 15444 12164 15456
rect 12216 15444 12222 15496
rect 13004 15493 13032 15524
rect 12897 15487 12955 15493
rect 12897 15453 12909 15487
rect 12943 15453 12955 15487
rect 12897 15447 12955 15453
rect 12989 15487 13047 15493
rect 12989 15453 13001 15487
rect 13035 15453 13047 15487
rect 12989 15447 13047 15453
rect 12912 15416 12940 15447
rect 13078 15444 13084 15496
rect 13136 15484 13142 15496
rect 13136 15456 13181 15484
rect 13136 15444 13142 15456
rect 13262 15444 13268 15496
rect 13320 15484 13326 15496
rect 13320 15456 13365 15484
rect 13320 15444 13326 15456
rect 14182 15444 14188 15496
rect 14240 15484 14246 15496
rect 14366 15484 14372 15496
rect 14240 15456 14372 15484
rect 14240 15444 14246 15456
rect 14366 15444 14372 15456
rect 14424 15484 14430 15496
rect 15948 15493 15976 15592
rect 25406 15580 25412 15632
rect 25464 15620 25470 15632
rect 25685 15623 25743 15629
rect 25685 15620 25697 15623
rect 25464 15592 25697 15620
rect 25464 15580 25470 15592
rect 25685 15589 25697 15592
rect 25731 15589 25743 15623
rect 25685 15583 25743 15589
rect 19794 15552 19800 15564
rect 19720 15524 19800 15552
rect 14553 15487 14611 15493
rect 14553 15484 14565 15487
rect 14424 15456 14565 15484
rect 14424 15444 14430 15456
rect 14553 15453 14565 15456
rect 14599 15453 14611 15487
rect 14553 15447 14611 15453
rect 15933 15487 15991 15493
rect 15933 15453 15945 15487
rect 15979 15484 15991 15487
rect 16393 15487 16451 15493
rect 16393 15484 16405 15487
rect 15979 15456 16405 15484
rect 15979 15453 15991 15456
rect 15933 15447 15991 15453
rect 16393 15453 16405 15456
rect 16439 15453 16451 15487
rect 16393 15447 16451 15453
rect 16482 15444 16488 15496
rect 16540 15484 16546 15496
rect 17313 15487 17371 15493
rect 17313 15484 17325 15487
rect 16540 15456 17325 15484
rect 16540 15444 16546 15456
rect 17313 15453 17325 15456
rect 17359 15453 17371 15487
rect 17313 15447 17371 15453
rect 17580 15487 17638 15493
rect 17580 15453 17592 15487
rect 17626 15484 17638 15487
rect 18046 15484 18052 15496
rect 17626 15456 18052 15484
rect 17626 15453 17638 15456
rect 17580 15447 17638 15453
rect 18046 15444 18052 15456
rect 18104 15444 18110 15496
rect 19426 15484 19432 15496
rect 19387 15456 19432 15484
rect 19426 15444 19432 15456
rect 19484 15444 19490 15496
rect 19720 15493 19748 15524
rect 19794 15512 19800 15524
rect 19852 15512 19858 15564
rect 20714 15552 20720 15564
rect 20272 15524 20720 15552
rect 19522 15487 19580 15493
rect 19522 15453 19534 15487
rect 19568 15453 19580 15487
rect 19522 15447 19580 15453
rect 19705 15487 19763 15493
rect 19705 15453 19717 15487
rect 19751 15453 19763 15487
rect 19705 15447 19763 15453
rect 19935 15487 19993 15493
rect 19935 15453 19947 15487
rect 19981 15484 19993 15487
rect 20070 15484 20076 15496
rect 19981 15456 20076 15484
rect 19981 15453 19993 15456
rect 19935 15447 19993 15453
rect 13354 15416 13360 15428
rect 12912 15388 13360 15416
rect 13354 15376 13360 15388
rect 13412 15376 13418 15428
rect 13538 15376 13544 15428
rect 13596 15416 13602 15428
rect 14737 15419 14795 15425
rect 14737 15416 14749 15419
rect 13596 15388 14749 15416
rect 13596 15376 13602 15388
rect 14737 15385 14749 15388
rect 14783 15416 14795 15419
rect 15470 15416 15476 15428
rect 14783 15388 15476 15416
rect 14783 15385 14795 15388
rect 14737 15379 14795 15385
rect 15470 15376 15476 15388
rect 15528 15376 15534 15428
rect 17954 15376 17960 15428
rect 18012 15416 18018 15428
rect 19536 15416 19564 15447
rect 20070 15444 20076 15456
rect 20128 15484 20134 15496
rect 20272 15484 20300 15524
rect 20714 15512 20720 15524
rect 20772 15512 20778 15564
rect 24854 15512 24860 15564
rect 24912 15552 24918 15564
rect 25884 15552 25912 15651
rect 27338 15648 27344 15660
rect 27396 15648 27402 15700
rect 28626 15648 28632 15700
rect 28684 15688 28690 15700
rect 29549 15691 29607 15697
rect 29549 15688 29561 15691
rect 28684 15660 29561 15688
rect 28684 15648 28690 15660
rect 29549 15657 29561 15660
rect 29595 15657 29607 15691
rect 35437 15691 35495 15697
rect 35437 15688 35449 15691
rect 29549 15651 29607 15657
rect 29656 15660 35449 15688
rect 26881 15623 26939 15629
rect 26881 15620 26893 15623
rect 25976 15592 26893 15620
rect 25976 15561 26004 15592
rect 26881 15589 26893 15592
rect 26927 15589 26939 15623
rect 29656 15620 29684 15660
rect 35437 15657 35449 15660
rect 35483 15657 35495 15691
rect 35437 15651 35495 15657
rect 37090 15648 37096 15700
rect 37148 15688 37154 15700
rect 37734 15688 37740 15700
rect 37148 15660 37740 15688
rect 37148 15648 37154 15660
rect 37734 15648 37740 15660
rect 37792 15688 37798 15700
rect 38838 15688 38844 15700
rect 37792 15660 37872 15688
rect 38799 15660 38844 15688
rect 37792 15648 37798 15660
rect 26881 15583 26939 15589
rect 27080 15592 29684 15620
rect 24912 15524 25912 15552
rect 25961 15555 26019 15561
rect 24912 15512 24918 15524
rect 25961 15521 25973 15555
rect 26007 15521 26019 15555
rect 25961 15515 26019 15521
rect 20128 15456 20300 15484
rect 20128 15444 20134 15456
rect 20346 15444 20352 15496
rect 20404 15484 20410 15496
rect 20533 15487 20591 15493
rect 20533 15484 20545 15487
rect 20404 15456 20545 15484
rect 20404 15444 20410 15456
rect 20533 15453 20545 15456
rect 20579 15453 20591 15487
rect 22002 15484 22008 15496
rect 21963 15456 22008 15484
rect 20533 15447 20591 15453
rect 22002 15444 22008 15456
rect 22060 15444 22066 15496
rect 22094 15444 22100 15496
rect 22152 15484 22158 15496
rect 22278 15484 22284 15496
rect 22152 15456 22197 15484
rect 22239 15456 22284 15484
rect 22152 15444 22158 15456
rect 22278 15444 22284 15456
rect 22336 15444 22342 15496
rect 25041 15487 25099 15493
rect 25041 15484 25053 15487
rect 24688 15456 25053 15484
rect 18012 15388 19564 15416
rect 19797 15419 19855 15425
rect 18012 15376 18018 15388
rect 19797 15385 19809 15419
rect 19843 15416 19855 15419
rect 24688 15416 24716 15456
rect 25041 15453 25053 15456
rect 25087 15484 25099 15487
rect 25866 15484 25872 15496
rect 25087 15456 25872 15484
rect 25087 15453 25099 15456
rect 25041 15447 25099 15453
rect 25866 15444 25872 15456
rect 25924 15444 25930 15496
rect 26050 15484 26056 15496
rect 26011 15456 26056 15484
rect 26050 15444 26056 15456
rect 26108 15444 26114 15496
rect 27080 15493 27108 15592
rect 32858 15580 32864 15632
rect 32916 15580 32922 15632
rect 33686 15620 33692 15632
rect 33647 15592 33692 15620
rect 33686 15580 33692 15592
rect 33744 15580 33750 15632
rect 37642 15580 37648 15632
rect 37700 15580 37706 15632
rect 37844 15620 37872 15660
rect 38838 15648 38844 15660
rect 38896 15648 38902 15700
rect 37844 15592 37964 15620
rect 29730 15552 29736 15564
rect 28368 15524 29736 15552
rect 27065 15487 27123 15493
rect 27065 15453 27077 15487
rect 27111 15453 27123 15487
rect 27065 15447 27123 15453
rect 27154 15444 27160 15496
rect 27212 15484 27218 15496
rect 27212 15456 27257 15484
rect 27212 15444 27218 15456
rect 28166 15444 28172 15496
rect 28224 15484 28230 15496
rect 28368 15493 28396 15524
rect 29730 15512 29736 15524
rect 29788 15512 29794 15564
rect 32490 15512 32496 15564
rect 32548 15552 32554 15564
rect 32548 15524 32700 15552
rect 32548 15512 32554 15524
rect 28261 15487 28319 15493
rect 28261 15484 28273 15487
rect 28224 15456 28273 15484
rect 28224 15444 28230 15456
rect 28261 15453 28273 15456
rect 28307 15453 28319 15487
rect 28261 15447 28319 15453
rect 28353 15487 28411 15493
rect 28353 15453 28365 15487
rect 28399 15453 28411 15487
rect 28353 15447 28411 15453
rect 28629 15487 28687 15493
rect 28629 15453 28641 15487
rect 28675 15453 28687 15487
rect 28629 15447 28687 15453
rect 19843 15388 24716 15416
rect 24857 15419 24915 15425
rect 19843 15385 19855 15388
rect 19797 15379 19855 15385
rect 24857 15385 24869 15419
rect 24903 15416 24915 15419
rect 25130 15416 25136 15428
rect 24903 15388 25136 15416
rect 24903 15385 24915 15388
rect 24857 15379 24915 15385
rect 25130 15376 25136 15388
rect 25188 15376 25194 15428
rect 27246 15376 27252 15428
rect 27304 15416 27310 15428
rect 27341 15419 27399 15425
rect 27341 15416 27353 15419
rect 27304 15388 27353 15416
rect 27304 15376 27310 15388
rect 27341 15385 27353 15388
rect 27387 15385 27399 15419
rect 27341 15379 27399 15385
rect 28445 15419 28503 15425
rect 28445 15385 28457 15419
rect 28491 15385 28503 15419
rect 28644 15416 28672 15447
rect 28994 15444 29000 15496
rect 29052 15484 29058 15496
rect 30193 15487 30251 15493
rect 30193 15484 30205 15487
rect 29052 15456 30205 15484
rect 29052 15444 29058 15456
rect 30193 15453 30205 15456
rect 30239 15453 30251 15487
rect 30193 15447 30251 15453
rect 32306 15444 32312 15496
rect 32364 15484 32370 15496
rect 32585 15487 32643 15493
rect 32585 15484 32597 15487
rect 32364 15456 32597 15484
rect 32364 15444 32370 15456
rect 32585 15453 32597 15456
rect 32631 15453 32643 15487
rect 32672 15484 32700 15524
rect 32876 15493 32904 15580
rect 35802 15552 35808 15564
rect 35636 15524 35808 15552
rect 35636 15493 35664 15524
rect 35802 15512 35808 15524
rect 35860 15512 35866 15564
rect 36909 15555 36967 15561
rect 36909 15521 36921 15555
rect 36955 15552 36967 15555
rect 36955 15524 37591 15552
rect 36955 15521 36967 15524
rect 36909 15515 36967 15521
rect 32748 15487 32806 15493
rect 32748 15484 32760 15487
rect 32672 15456 32760 15484
rect 32585 15447 32643 15453
rect 32748 15453 32760 15456
rect 32794 15453 32806 15487
rect 32748 15447 32806 15453
rect 32864 15487 32922 15493
rect 32864 15453 32876 15487
rect 32910 15453 32922 15487
rect 32864 15447 32922 15453
rect 32953 15487 33011 15493
rect 32953 15453 32965 15487
rect 32999 15453 33011 15487
rect 32953 15447 33011 15453
rect 35621 15487 35679 15493
rect 35621 15453 35633 15487
rect 35667 15453 35679 15487
rect 35621 15447 35679 15453
rect 35713 15487 35771 15493
rect 35713 15453 35725 15487
rect 35759 15484 35771 15487
rect 35759 15456 35940 15484
rect 35759 15453 35771 15456
rect 35713 15447 35771 15453
rect 29454 15416 29460 15428
rect 28644 15388 29460 15416
rect 28445 15379 28503 15385
rect 12618 15348 12624 15360
rect 6972 15320 9168 15348
rect 12579 15320 12624 15348
rect 6972 15308 6978 15320
rect 12618 15308 12624 15320
rect 12676 15308 12682 15360
rect 20070 15348 20076 15360
rect 20031 15320 20076 15348
rect 20070 15308 20076 15320
rect 20128 15308 20134 15360
rect 25222 15348 25228 15360
rect 25183 15320 25228 15348
rect 25222 15308 25228 15320
rect 25280 15308 25286 15360
rect 28074 15348 28080 15360
rect 28035 15320 28080 15348
rect 28074 15308 28080 15320
rect 28132 15308 28138 15360
rect 28460 15348 28488 15379
rect 29454 15376 29460 15388
rect 29512 15376 29518 15428
rect 29546 15376 29552 15428
rect 29604 15416 29610 15428
rect 30438 15419 30496 15425
rect 30438 15416 30450 15419
rect 29604 15388 30450 15416
rect 29604 15376 29610 15388
rect 30438 15385 30450 15388
rect 30484 15385 30496 15419
rect 32600 15416 32628 15447
rect 32968 15416 32996 15447
rect 32600 15388 32812 15416
rect 32968 15388 33088 15416
rect 30438 15379 30496 15385
rect 32784 15360 32812 15388
rect 28626 15348 28632 15360
rect 28460 15320 28632 15348
rect 28626 15308 28632 15320
rect 28684 15308 28690 15360
rect 31018 15308 31024 15360
rect 31076 15348 31082 15360
rect 31573 15351 31631 15357
rect 31573 15348 31585 15351
rect 31076 15320 31585 15348
rect 31076 15308 31082 15320
rect 31573 15317 31585 15320
rect 31619 15317 31631 15351
rect 31573 15311 31631 15317
rect 32125 15351 32183 15357
rect 32125 15317 32137 15351
rect 32171 15348 32183 15351
rect 32582 15348 32588 15360
rect 32171 15320 32588 15348
rect 32171 15317 32183 15320
rect 32125 15311 32183 15317
rect 32582 15308 32588 15320
rect 32640 15308 32646 15360
rect 32766 15308 32772 15360
rect 32824 15308 32830 15360
rect 32950 15308 32956 15360
rect 33008 15348 33014 15360
rect 33060 15348 33088 15388
rect 35342 15376 35348 15428
rect 35400 15416 35406 15428
rect 35805 15419 35863 15425
rect 35805 15416 35817 15419
rect 35400 15388 35817 15416
rect 35400 15376 35406 15388
rect 35805 15385 35817 15388
rect 35851 15385 35863 15419
rect 35912 15416 35940 15456
rect 35986 15444 35992 15496
rect 36044 15484 36050 15496
rect 36541 15487 36599 15493
rect 36044 15456 36089 15484
rect 36044 15444 36050 15456
rect 36541 15453 36553 15487
rect 36587 15484 36599 15487
rect 37274 15484 37280 15496
rect 36587 15456 37280 15484
rect 36587 15453 36599 15456
rect 36541 15447 36599 15453
rect 37274 15444 37280 15456
rect 37332 15444 37338 15496
rect 37563 15493 37591 15524
rect 37663 15493 37691 15580
rect 37369 15487 37427 15493
rect 37369 15453 37381 15487
rect 37415 15484 37427 15487
rect 37548 15487 37606 15493
rect 37415 15456 37504 15484
rect 37415 15453 37427 15456
rect 37369 15447 37427 15453
rect 37476 15428 37504 15456
rect 37548 15453 37560 15487
rect 37594 15453 37606 15487
rect 37548 15447 37606 15453
rect 37648 15487 37706 15493
rect 37648 15453 37660 15487
rect 37694 15453 37706 15487
rect 37648 15447 37706 15453
rect 37737 15487 37795 15493
rect 37737 15453 37749 15487
rect 37783 15453 37795 15487
rect 37737 15447 37795 15453
rect 36725 15419 36783 15425
rect 36725 15416 36737 15419
rect 35912 15388 36737 15416
rect 35805 15379 35863 15385
rect 36725 15385 36737 15388
rect 36771 15385 36783 15419
rect 36725 15379 36783 15385
rect 33226 15348 33232 15360
rect 33008 15320 33088 15348
rect 33187 15320 33232 15348
rect 33008 15308 33014 15320
rect 33226 15308 33232 15320
rect 33284 15308 33290 15360
rect 33318 15308 33324 15360
rect 33376 15348 33382 15360
rect 35710 15348 35716 15360
rect 33376 15320 35716 15348
rect 33376 15308 33382 15320
rect 35710 15308 35716 15320
rect 35768 15308 35774 15360
rect 35820 15348 35848 15379
rect 36262 15348 36268 15360
rect 35820 15320 36268 15348
rect 36262 15308 36268 15320
rect 36320 15308 36326 15360
rect 36740 15348 36768 15379
rect 37458 15376 37464 15428
rect 37516 15376 37522 15428
rect 37752 15416 37780 15447
rect 37936 15416 37964 15592
rect 41230 15552 41236 15564
rect 41191 15524 41236 15552
rect 41230 15512 41236 15524
rect 41288 15512 41294 15564
rect 40966 15487 41024 15493
rect 40966 15484 40978 15487
rect 38028 15456 40978 15484
rect 38028 15425 38056 15456
rect 40966 15453 40978 15456
rect 41012 15453 41024 15487
rect 40966 15447 41024 15453
rect 37752 15388 37964 15416
rect 38013 15419 38071 15425
rect 38013 15385 38025 15419
rect 38059 15385 38071 15419
rect 38470 15416 38476 15428
rect 38431 15388 38476 15416
rect 38013 15379 38071 15385
rect 38470 15376 38476 15388
rect 38528 15376 38534 15428
rect 38654 15416 38660 15428
rect 38615 15388 38660 15416
rect 38654 15376 38660 15388
rect 38712 15376 38718 15428
rect 39853 15351 39911 15357
rect 39853 15348 39865 15351
rect 36740 15320 39865 15348
rect 39853 15317 39865 15320
rect 39899 15317 39911 15351
rect 39853 15311 39911 15317
rect 1104 15258 68816 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 68816 15258
rect 1104 15184 68816 15206
rect 3786 15104 3792 15156
rect 3844 15144 3850 15156
rect 8021 15147 8079 15153
rect 8021 15144 8033 15147
rect 3844 15116 8033 15144
rect 3844 15104 3850 15116
rect 8021 15113 8033 15116
rect 8067 15113 8079 15147
rect 8021 15107 8079 15113
rect 2133 15079 2191 15085
rect 2133 15045 2145 15079
rect 2179 15076 2191 15079
rect 4798 15076 4804 15088
rect 2179 15048 4804 15076
rect 2179 15045 2191 15048
rect 2133 15039 2191 15045
rect 4798 15036 4804 15048
rect 4856 15036 4862 15088
rect 5350 15076 5356 15088
rect 5311 15048 5356 15076
rect 5350 15036 5356 15048
rect 5408 15036 5414 15088
rect 6733 15079 6791 15085
rect 6733 15045 6745 15079
rect 6779 15076 6791 15079
rect 6822 15076 6828 15088
rect 6779 15048 6828 15076
rect 6779 15045 6791 15048
rect 6733 15039 6791 15045
rect 6822 15036 6828 15048
rect 6880 15036 6886 15088
rect 1949 15011 2007 15017
rect 1949 14977 1961 15011
rect 1995 15008 2007 15011
rect 4062 15008 4068 15020
rect 1995 14980 4068 15008
rect 1995 14977 2007 14980
rect 1949 14971 2007 14977
rect 4062 14968 4068 14980
rect 4120 14968 4126 15020
rect 5074 15008 5080 15020
rect 5035 14980 5080 15008
rect 5074 14968 5080 14980
rect 5132 14968 5138 15020
rect 5258 15008 5264 15020
rect 5219 14980 5264 15008
rect 5258 14968 5264 14980
rect 5316 14968 5322 15020
rect 5445 15011 5503 15017
rect 5445 14977 5457 15011
rect 5491 15008 5503 15011
rect 6546 15008 6552 15020
rect 5491 14980 6552 15008
rect 5491 14977 5503 14980
rect 5445 14971 5503 14977
rect 6546 14968 6552 14980
rect 6604 15008 6610 15020
rect 7742 15008 7748 15020
rect 6604 14980 7748 15008
rect 6604 14968 6610 14980
rect 7742 14968 7748 14980
rect 7800 14968 7806 15020
rect 8036 15008 8064 15107
rect 10134 15104 10140 15156
rect 10192 15144 10198 15156
rect 10318 15144 10324 15156
rect 10192 15116 10324 15144
rect 10192 15104 10198 15116
rect 10318 15104 10324 15116
rect 10376 15104 10382 15156
rect 12526 15104 12532 15156
rect 12584 15144 12590 15156
rect 15194 15144 15200 15156
rect 12584 15116 15200 15144
rect 12584 15104 12590 15116
rect 15194 15104 15200 15116
rect 15252 15144 15258 15156
rect 15657 15147 15715 15153
rect 15657 15144 15669 15147
rect 15252 15116 15669 15144
rect 15252 15104 15258 15116
rect 15657 15113 15669 15116
rect 15703 15113 15715 15147
rect 15657 15107 15715 15113
rect 10226 15036 10232 15088
rect 10284 15076 10290 15088
rect 11054 15076 11060 15088
rect 10284 15048 11060 15076
rect 10284 15036 10290 15048
rect 11054 15036 11060 15048
rect 11112 15036 11118 15088
rect 11701 15079 11759 15085
rect 11701 15045 11713 15079
rect 11747 15076 11759 15079
rect 12434 15076 12440 15088
rect 11747 15048 12440 15076
rect 11747 15045 11759 15048
rect 11701 15039 11759 15045
rect 12434 15036 12440 15048
rect 12492 15036 12498 15088
rect 12618 15036 12624 15088
rect 12676 15076 12682 15088
rect 12774 15079 12832 15085
rect 12774 15076 12786 15079
rect 12676 15048 12786 15076
rect 12676 15036 12682 15048
rect 12774 15045 12786 15048
rect 12820 15045 12832 15079
rect 12774 15039 12832 15045
rect 8941 15011 8999 15017
rect 8941 15008 8953 15011
rect 8036 14980 8953 15008
rect 8941 14977 8953 14980
rect 8987 15008 8999 15011
rect 9030 15008 9036 15020
rect 8987 14980 9036 15008
rect 8987 14977 8999 14980
rect 8941 14971 8999 14977
rect 9030 14968 9036 14980
rect 9088 14968 9094 15020
rect 9214 15017 9220 15020
rect 9208 14971 9220 15017
rect 9272 15008 9278 15020
rect 11882 15008 11888 15020
rect 9272 14980 9308 15008
rect 11843 14980 11888 15008
rect 9214 14968 9220 14971
rect 9272 14968 9278 14980
rect 11882 14968 11888 14980
rect 11940 14968 11946 15020
rect 14366 15008 14372 15020
rect 14327 14980 14372 15008
rect 14366 14968 14372 14980
rect 14424 14968 14430 15020
rect 15672 15008 15700 15107
rect 17954 15104 17960 15156
rect 18012 15144 18018 15156
rect 18049 15147 18107 15153
rect 18049 15144 18061 15147
rect 18012 15116 18061 15144
rect 18012 15104 18018 15116
rect 18049 15113 18061 15116
rect 18095 15113 18107 15147
rect 18049 15107 18107 15113
rect 22002 15104 22008 15156
rect 22060 15144 22066 15156
rect 28902 15144 28908 15156
rect 22060 15116 28212 15144
rect 28863 15116 28908 15144
rect 22060 15104 22066 15116
rect 17586 15036 17592 15088
rect 17644 15076 17650 15088
rect 18966 15076 18972 15088
rect 17644 15048 18972 15076
rect 17644 15036 17650 15048
rect 18966 15036 18972 15048
rect 19024 15036 19030 15088
rect 20990 15076 20996 15088
rect 20456 15048 20996 15076
rect 16482 15008 16488 15020
rect 15672 14980 16488 15008
rect 16482 14968 16488 14980
rect 16540 15008 16546 15020
rect 16669 15011 16727 15017
rect 16669 15008 16681 15011
rect 16540 14980 16681 15008
rect 16540 14968 16546 14980
rect 16669 14977 16681 14980
rect 16715 14977 16727 15011
rect 16669 14971 16727 14977
rect 16758 14968 16764 15020
rect 16816 15008 16822 15020
rect 20456 15017 20484 15048
rect 20990 15036 20996 15048
rect 21048 15036 21054 15088
rect 24854 15036 24860 15088
rect 24912 15076 24918 15088
rect 25041 15079 25099 15085
rect 25041 15076 25053 15079
rect 24912 15048 25053 15076
rect 24912 15036 24918 15048
rect 25041 15045 25053 15048
rect 25087 15045 25099 15079
rect 25041 15039 25099 15045
rect 26145 15079 26203 15085
rect 26145 15045 26157 15079
rect 26191 15076 26203 15079
rect 28086 15079 28144 15085
rect 28086 15076 28098 15079
rect 26191 15048 28098 15076
rect 26191 15045 26203 15048
rect 26145 15039 26203 15045
rect 28086 15045 28098 15048
rect 28132 15045 28144 15079
rect 28184 15076 28212 15116
rect 28902 15104 28908 15116
rect 28960 15104 28966 15156
rect 29546 15144 29552 15156
rect 29507 15116 29552 15144
rect 29546 15104 29552 15116
rect 29604 15104 29610 15156
rect 30837 15147 30895 15153
rect 30837 15113 30849 15147
rect 30883 15144 30895 15147
rect 32490 15144 32496 15156
rect 30883 15116 31754 15144
rect 32451 15116 32496 15144
rect 30883 15113 30895 15116
rect 30837 15107 30895 15113
rect 28184 15048 29132 15076
rect 28086 15039 28144 15045
rect 16925 15011 16983 15017
rect 16925 15008 16937 15011
rect 16816 14980 16937 15008
rect 16816 14968 16822 14980
rect 16925 14977 16937 14980
rect 16971 14977 16983 15011
rect 16925 14971 16983 14977
rect 20441 15011 20499 15017
rect 20441 14977 20453 15011
rect 20487 14977 20499 15011
rect 20714 15008 20720 15020
rect 20675 14980 20720 15008
rect 20441 14971 20499 14977
rect 20714 14968 20720 14980
rect 20772 14968 20778 15020
rect 22002 15008 22008 15020
rect 21963 14980 22008 15008
rect 22002 14968 22008 14980
rect 22060 14968 22066 15020
rect 22278 15008 22284 15020
rect 22239 14980 22284 15008
rect 22278 14968 22284 14980
rect 22336 14968 22342 15020
rect 24049 15011 24107 15017
rect 24049 14977 24061 15011
rect 24095 15008 24107 15011
rect 24946 15008 24952 15020
rect 24095 14980 24952 15008
rect 24095 14977 24107 14980
rect 24049 14971 24107 14977
rect 24946 14968 24952 14980
rect 25004 14968 25010 15020
rect 25314 14968 25320 15020
rect 25372 15008 25378 15020
rect 25664 15017 25722 15023
rect 25501 15011 25559 15017
rect 25664 15014 25676 15017
rect 25501 15008 25513 15011
rect 25372 14980 25513 15008
rect 25372 14968 25378 14980
rect 25501 14977 25513 14980
rect 25547 14977 25559 15011
rect 25501 14971 25559 14977
rect 25608 14986 25676 15014
rect 6822 14900 6828 14952
rect 6880 14940 6886 14952
rect 7190 14940 7196 14952
rect 6880 14912 7196 14940
rect 6880 14900 6886 14912
rect 7190 14900 7196 14912
rect 7248 14900 7254 14952
rect 12526 14940 12532 14952
rect 12487 14912 12532 14940
rect 12526 14900 12532 14912
rect 12584 14900 12590 14952
rect 22186 14940 22192 14952
rect 22147 14912 22192 14940
rect 22186 14900 22192 14912
rect 22244 14900 22250 14952
rect 24302 14940 24308 14952
rect 24263 14912 24308 14940
rect 24302 14900 24308 14912
rect 24360 14900 24366 14952
rect 25222 14900 25228 14952
rect 25280 14940 25286 14952
rect 25608 14940 25636 14986
rect 25664 14983 25676 14986
rect 25710 14983 25722 15017
rect 25664 14977 25722 14983
rect 25764 15017 25822 15023
rect 25764 14983 25776 15017
rect 25810 14983 25822 15017
rect 25764 14977 25822 14983
rect 25869 15011 25927 15017
rect 25869 14977 25881 15011
rect 25915 15008 25927 15011
rect 26234 15008 26240 15020
rect 25915 14980 26240 15008
rect 25915 14977 25927 14980
rect 25792 14940 25820 14977
rect 25869 14971 25927 14977
rect 26234 14968 26240 14980
rect 26292 14968 26298 15020
rect 28353 15011 28411 15017
rect 28353 14977 28365 15011
rect 28399 15008 28411 15011
rect 28994 15008 29000 15020
rect 28399 14980 29000 15008
rect 28399 14977 28411 14980
rect 28353 14971 28411 14977
rect 28994 14968 29000 14980
rect 29052 14968 29058 15020
rect 25280 14912 25636 14940
rect 25709 14912 25820 14940
rect 25280 14900 25286 14912
rect 5626 14872 5632 14884
rect 5587 14844 5632 14872
rect 5626 14832 5632 14844
rect 5684 14832 5690 14884
rect 5718 14832 5724 14884
rect 5776 14872 5782 14884
rect 8202 14872 8208 14884
rect 5776 14844 8208 14872
rect 5776 14832 5782 14844
rect 8202 14832 8208 14844
rect 8260 14832 8266 14884
rect 13906 14872 13912 14884
rect 13867 14844 13912 14872
rect 13906 14832 13912 14844
rect 13964 14832 13970 14884
rect 22922 14872 22928 14884
rect 22296 14844 22600 14872
rect 22883 14844 22928 14872
rect 1765 14807 1823 14813
rect 1765 14773 1777 14807
rect 1811 14804 1823 14807
rect 1946 14804 1952 14816
rect 1811 14776 1952 14804
rect 1811 14773 1823 14776
rect 1765 14767 1823 14773
rect 1946 14764 1952 14776
rect 2004 14764 2010 14816
rect 4062 14764 4068 14816
rect 4120 14804 4126 14816
rect 10502 14804 10508 14816
rect 4120 14776 10508 14804
rect 4120 14764 4126 14776
rect 10502 14764 10508 14776
rect 10560 14764 10566 14816
rect 11974 14764 11980 14816
rect 12032 14804 12038 14816
rect 22296 14813 22324 14844
rect 12069 14807 12127 14813
rect 12069 14804 12081 14807
rect 12032 14776 12081 14804
rect 12032 14764 12038 14776
rect 12069 14773 12081 14776
rect 12115 14773 12127 14807
rect 12069 14767 12127 14773
rect 22281 14807 22339 14813
rect 22281 14773 22293 14807
rect 22327 14773 22339 14807
rect 22281 14767 22339 14773
rect 22370 14764 22376 14816
rect 22428 14804 22434 14816
rect 22465 14807 22523 14813
rect 22465 14804 22477 14807
rect 22428 14776 22477 14804
rect 22428 14764 22434 14776
rect 22465 14773 22477 14776
rect 22511 14773 22523 14807
rect 22572 14804 22600 14844
rect 22922 14832 22928 14844
rect 22980 14832 22986 14884
rect 25709 14872 25737 14912
rect 25774 14872 25780 14884
rect 25709 14844 25780 14872
rect 25774 14832 25780 14844
rect 25832 14832 25838 14884
rect 25866 14832 25872 14884
rect 25924 14872 25930 14884
rect 26973 14875 27031 14881
rect 26973 14872 26985 14875
rect 25924 14844 26985 14872
rect 25924 14832 25930 14844
rect 26973 14841 26985 14844
rect 27019 14841 27031 14875
rect 29104 14872 29132 15048
rect 29270 15036 29276 15088
rect 29328 15076 29334 15088
rect 29328 15048 29960 15076
rect 29328 15036 29334 15048
rect 29638 14968 29644 15020
rect 29696 15008 29702 15020
rect 29932 15017 29960 15048
rect 31110 15036 31116 15088
rect 31168 15076 31174 15088
rect 31297 15079 31355 15085
rect 31297 15076 31309 15079
rect 31168 15048 31309 15076
rect 31168 15036 31174 15048
rect 31297 15045 31309 15048
rect 31343 15045 31355 15079
rect 31726 15076 31754 15116
rect 32490 15104 32496 15116
rect 32548 15104 32554 15156
rect 33045 15147 33103 15153
rect 33045 15113 33057 15147
rect 33091 15113 33103 15147
rect 33045 15107 33103 15113
rect 35897 15147 35955 15153
rect 35897 15113 35909 15147
rect 35943 15144 35955 15147
rect 35986 15144 35992 15156
rect 35943 15116 35992 15144
rect 35943 15113 35955 15116
rect 35897 15107 35955 15113
rect 32122 15076 32128 15088
rect 31726 15048 32128 15076
rect 31297 15039 31355 15045
rect 32122 15036 32128 15048
rect 32180 15036 32186 15088
rect 32306 15076 32312 15088
rect 32219 15048 32312 15076
rect 32306 15036 32312 15048
rect 32364 15076 32370 15088
rect 33060 15076 33088 15107
rect 35986 15104 35992 15116
rect 36044 15104 36050 15156
rect 36096 15116 37274 15144
rect 32364 15048 33088 15076
rect 32364 15036 32370 15048
rect 33226 15036 33232 15088
rect 33284 15076 33290 15088
rect 34158 15079 34216 15085
rect 34158 15076 34170 15079
rect 33284 15048 34170 15076
rect 33284 15036 33290 15048
rect 34158 15045 34170 15048
rect 34204 15045 34216 15079
rect 34158 15039 34216 15045
rect 35161 15079 35219 15085
rect 35161 15045 35173 15079
rect 35207 15076 35219 15079
rect 36096 15076 36124 15116
rect 35207 15048 36124 15076
rect 35207 15045 35219 15048
rect 35161 15039 35219 15045
rect 36262 15036 36268 15088
rect 36320 15076 36326 15088
rect 37246 15076 37274 15116
rect 37366 15104 37372 15156
rect 37424 15144 37430 15156
rect 38470 15144 38476 15156
rect 37424 15116 38476 15144
rect 37424 15104 37430 15116
rect 38470 15104 38476 15116
rect 38528 15104 38534 15156
rect 38654 15076 38660 15088
rect 36320 15048 36365 15076
rect 37246 15048 38660 15076
rect 36320 15036 36326 15048
rect 38654 15036 38660 15048
rect 38712 15036 38718 15088
rect 29825 15011 29883 15017
rect 29825 15008 29837 15011
rect 29696 14980 29837 15008
rect 29696 14968 29702 14980
rect 29825 14977 29837 14980
rect 29871 14977 29883 15011
rect 29825 14971 29883 14977
rect 29917 15011 29975 15017
rect 29917 14977 29929 15011
rect 29963 14977 29975 15011
rect 29917 14971 29975 14977
rect 30006 14968 30012 15020
rect 30064 15008 30070 15020
rect 30193 15011 30251 15017
rect 30064 14980 30109 15008
rect 30064 14968 30070 14980
rect 30193 14977 30205 15011
rect 30239 14977 30251 15011
rect 30193 14971 30251 14977
rect 30653 15011 30711 15017
rect 30653 14977 30665 15011
rect 30699 15008 30711 15011
rect 31386 15008 31392 15020
rect 30699 14980 31392 15008
rect 30699 14977 30711 14980
rect 30653 14971 30711 14977
rect 30208 14940 30236 14971
rect 31386 14968 31392 14980
rect 31444 14968 31450 15020
rect 31478 14968 31484 15020
rect 31536 15008 31542 15020
rect 35069 15011 35127 15017
rect 31536 14980 31581 15008
rect 33428 14980 34928 15008
rect 31536 14968 31542 14980
rect 30926 14940 30932 14952
rect 30208 14912 30932 14940
rect 30926 14900 30932 14912
rect 30984 14940 30990 14952
rect 33428 14940 33456 14980
rect 34422 14940 34428 14952
rect 30984 14912 33456 14940
rect 34383 14912 34428 14940
rect 30984 14900 30990 14912
rect 34422 14900 34428 14912
rect 34480 14900 34486 14952
rect 34900 14872 34928 14980
rect 35069 14977 35081 15011
rect 35115 14977 35127 15011
rect 35250 15008 35256 15020
rect 35211 14980 35256 15008
rect 35069 14971 35127 14977
rect 35084 14940 35112 14971
rect 35250 14968 35256 14980
rect 35308 14968 35314 15020
rect 35434 15008 35440 15020
rect 35395 14980 35440 15008
rect 35434 14968 35440 14980
rect 35492 14968 35498 15020
rect 35802 14968 35808 15020
rect 35860 15008 35866 15020
rect 36081 15011 36139 15017
rect 36081 15008 36093 15011
rect 35860 14980 36093 15008
rect 35860 14968 35866 14980
rect 36081 14977 36093 14980
rect 36127 14977 36139 15011
rect 36081 14971 36139 14977
rect 36173 15011 36231 15017
rect 36173 14977 36185 15011
rect 36219 15008 36231 15011
rect 36446 15008 36452 15020
rect 36219 14980 36308 15008
rect 36407 14980 36452 15008
rect 36219 14977 36231 14980
rect 36173 14971 36231 14977
rect 35820 14940 35848 14968
rect 35084 14912 35848 14940
rect 36280 14940 36308 14980
rect 36446 14968 36452 14980
rect 36504 14968 36510 15020
rect 37369 15011 37427 15017
rect 37369 14977 37381 15011
rect 37415 15008 37427 15011
rect 37550 15008 37556 15020
rect 37415 14980 37556 15008
rect 37415 14977 37427 14980
rect 37369 14971 37427 14977
rect 37550 14968 37556 14980
rect 37608 15008 37614 15020
rect 37734 15008 37740 15020
rect 37608 14980 37740 15008
rect 37608 14968 37614 14980
rect 37734 14968 37740 14980
rect 37792 14968 37798 15020
rect 36722 14940 36728 14952
rect 36280 14912 36728 14940
rect 36722 14900 36728 14912
rect 36780 14900 36786 14952
rect 29104 14844 33364 14872
rect 34900 14844 35204 14872
rect 26973 14835 27031 14841
rect 29362 14804 29368 14816
rect 22572 14776 29368 14804
rect 22465 14767 22523 14773
rect 29362 14764 29368 14776
rect 29420 14764 29426 14816
rect 33336 14804 33364 14844
rect 34885 14807 34943 14813
rect 34885 14804 34897 14807
rect 33336 14776 34897 14804
rect 34885 14773 34897 14776
rect 34931 14773 34943 14807
rect 35176 14804 35204 14844
rect 36906 14832 36912 14884
rect 36964 14872 36970 14884
rect 37829 14875 37887 14881
rect 37829 14872 37841 14875
rect 36964 14844 37841 14872
rect 36964 14832 36970 14844
rect 37829 14841 37841 14844
rect 37875 14872 37887 14875
rect 38010 14872 38016 14884
rect 37875 14844 38016 14872
rect 37875 14841 37887 14844
rect 37829 14835 37887 14841
rect 38010 14832 38016 14844
rect 38068 14832 38074 14884
rect 37458 14804 37464 14816
rect 35176 14776 37464 14804
rect 34885 14767 34943 14773
rect 37458 14764 37464 14776
rect 37516 14764 37522 14816
rect 1104 14714 68816 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 65654 14714
rect 65706 14662 65718 14714
rect 65770 14662 65782 14714
rect 65834 14662 65846 14714
rect 65898 14662 65910 14714
rect 65962 14662 68816 14714
rect 1104 14640 68816 14662
rect 7285 14603 7343 14609
rect 7285 14569 7297 14603
rect 7331 14600 7343 14603
rect 9214 14600 9220 14612
rect 7331 14572 9220 14600
rect 7331 14569 7343 14572
rect 7285 14563 7343 14569
rect 9214 14560 9220 14572
rect 9272 14560 9278 14612
rect 9766 14560 9772 14612
rect 9824 14600 9830 14612
rect 9861 14603 9919 14609
rect 9861 14600 9873 14603
rect 9824 14572 9873 14600
rect 9824 14560 9830 14572
rect 9861 14569 9873 14572
rect 9907 14600 9919 14603
rect 10778 14600 10784 14612
rect 9907 14572 10784 14600
rect 9907 14569 9919 14572
rect 9861 14563 9919 14569
rect 10778 14560 10784 14572
rect 10836 14560 10842 14612
rect 11882 14560 11888 14612
rect 11940 14600 11946 14612
rect 11977 14603 12035 14609
rect 11977 14600 11989 14603
rect 11940 14572 11989 14600
rect 11940 14560 11946 14572
rect 11977 14569 11989 14572
rect 12023 14600 12035 14603
rect 17218 14600 17224 14612
rect 12023 14572 12434 14600
rect 17179 14572 17224 14600
rect 12023 14569 12035 14572
rect 11977 14563 12035 14569
rect 2130 14492 2136 14544
rect 2188 14492 2194 14544
rect 2222 14492 2228 14544
rect 2280 14532 2286 14544
rect 2869 14535 2927 14541
rect 2869 14532 2881 14535
rect 2280 14504 2881 14532
rect 2280 14492 2286 14504
rect 2869 14501 2881 14504
rect 2915 14532 2927 14535
rect 7466 14532 7472 14544
rect 2915 14504 7472 14532
rect 2915 14501 2927 14504
rect 2869 14495 2927 14501
rect 7466 14492 7472 14504
rect 7524 14492 7530 14544
rect 9309 14535 9367 14541
rect 9309 14532 9321 14535
rect 7944 14504 9321 14532
rect 2148 14464 2176 14492
rect 4065 14467 4123 14473
rect 4065 14464 4077 14467
rect 2056 14436 4077 14464
rect 1762 14396 1768 14408
rect 1723 14368 1768 14396
rect 1762 14356 1768 14368
rect 1820 14356 1826 14408
rect 1946 14396 1952 14408
rect 1907 14368 1952 14396
rect 1946 14356 1952 14368
rect 2004 14356 2010 14408
rect 2056 14405 2084 14436
rect 4065 14433 4077 14436
rect 4111 14433 4123 14467
rect 6454 14464 6460 14476
rect 4065 14427 4123 14433
rect 4540 14436 6460 14464
rect 2041 14399 2099 14405
rect 2041 14365 2053 14399
rect 2087 14365 2099 14399
rect 2041 14359 2099 14365
rect 2133 14399 2191 14405
rect 2133 14365 2145 14399
rect 2179 14396 2191 14399
rect 2222 14396 2228 14408
rect 2179 14368 2228 14396
rect 2179 14365 2191 14368
rect 2133 14359 2191 14365
rect 2222 14356 2228 14368
rect 2280 14356 2286 14408
rect 3786 14396 3792 14408
rect 3699 14368 3792 14396
rect 3786 14356 3792 14368
rect 3844 14396 3850 14408
rect 4540 14396 4568 14436
rect 3844 14368 4568 14396
rect 3844 14356 3850 14368
rect 4890 14356 4896 14408
rect 4948 14396 4954 14408
rect 5077 14399 5135 14405
rect 5077 14396 5089 14399
rect 4948 14368 5089 14396
rect 4948 14356 4954 14368
rect 5077 14365 5089 14368
rect 5123 14365 5135 14399
rect 5258 14396 5264 14408
rect 5219 14368 5264 14396
rect 5077 14359 5135 14365
rect 5258 14356 5264 14368
rect 5316 14356 5322 14408
rect 5368 14405 5396 14436
rect 6454 14424 6460 14436
rect 6512 14424 6518 14476
rect 7834 14464 7840 14476
rect 6932 14436 7840 14464
rect 5353 14399 5411 14405
rect 5353 14365 5365 14399
rect 5399 14365 5411 14399
rect 5353 14359 5411 14365
rect 5445 14399 5503 14405
rect 5445 14365 5457 14399
rect 5491 14396 5503 14399
rect 5718 14396 5724 14408
rect 5491 14368 5724 14396
rect 5491 14365 5503 14368
rect 5445 14359 5503 14365
rect 5718 14356 5724 14368
rect 5776 14356 5782 14408
rect 6641 14399 6699 14405
rect 6641 14365 6653 14399
rect 6687 14365 6699 14399
rect 6822 14396 6828 14408
rect 6783 14368 6828 14396
rect 6641 14359 6699 14365
rect 6656 14328 6684 14359
rect 6822 14356 6828 14368
rect 6880 14356 6886 14408
rect 6932 14405 6960 14436
rect 7834 14424 7840 14436
rect 7892 14424 7898 14476
rect 6917 14399 6975 14405
rect 6917 14365 6929 14399
rect 6963 14365 6975 14399
rect 6917 14359 6975 14365
rect 7009 14399 7067 14405
rect 7009 14365 7021 14399
rect 7055 14396 7067 14399
rect 7466 14396 7472 14408
rect 7055 14368 7472 14396
rect 7055 14365 7067 14368
rect 7009 14359 7067 14365
rect 7466 14356 7472 14368
rect 7524 14356 7530 14408
rect 7650 14356 7656 14408
rect 7708 14396 7714 14408
rect 7944 14405 7972 14504
rect 9309 14501 9321 14504
rect 9355 14501 9367 14535
rect 9309 14495 9367 14501
rect 9030 14424 9036 14476
rect 9088 14464 9094 14476
rect 10597 14467 10655 14473
rect 10597 14464 10609 14467
rect 9088 14436 10609 14464
rect 9088 14424 9094 14436
rect 10597 14433 10609 14436
rect 10643 14433 10655 14467
rect 12406 14464 12434 14572
rect 17218 14560 17224 14572
rect 17276 14560 17282 14612
rect 20162 14560 20168 14612
rect 20220 14600 20226 14612
rect 22281 14603 22339 14609
rect 22281 14600 22293 14603
rect 20220 14572 22293 14600
rect 20220 14560 20226 14572
rect 22281 14569 22293 14572
rect 22327 14569 22339 14603
rect 22281 14563 22339 14569
rect 24946 14560 24952 14612
rect 25004 14600 25010 14612
rect 25041 14603 25099 14609
rect 25041 14600 25053 14603
rect 25004 14572 25053 14600
rect 25004 14560 25010 14572
rect 25041 14569 25053 14572
rect 25087 14569 25099 14603
rect 25041 14563 25099 14569
rect 26068 14572 28856 14600
rect 22097 14535 22155 14541
rect 22097 14501 22109 14535
rect 22143 14532 22155 14535
rect 22462 14532 22468 14544
rect 22143 14504 22468 14532
rect 22143 14501 22155 14504
rect 22097 14495 22155 14501
rect 22462 14492 22468 14504
rect 22520 14492 22526 14544
rect 25314 14492 25320 14544
rect 25372 14532 25378 14544
rect 25372 14504 25912 14532
rect 25372 14492 25378 14504
rect 15378 14464 15384 14476
rect 12406 14436 14964 14464
rect 10597 14427 10655 14433
rect 7745 14399 7803 14405
rect 7745 14396 7757 14399
rect 7708 14368 7757 14396
rect 7708 14356 7714 14368
rect 7745 14365 7757 14368
rect 7791 14365 7803 14399
rect 7745 14359 7803 14365
rect 7929 14399 7987 14405
rect 7929 14365 7941 14399
rect 7975 14365 7987 14399
rect 7929 14359 7987 14365
rect 8021 14399 8079 14405
rect 8021 14365 8033 14399
rect 8067 14365 8079 14399
rect 8021 14359 8079 14365
rect 8113 14399 8171 14405
rect 8113 14365 8125 14399
rect 8159 14396 8171 14399
rect 8202 14396 8208 14408
rect 8159 14368 8208 14396
rect 8159 14365 8171 14368
rect 8113 14359 8171 14365
rect 6656 14300 7052 14328
rect 7024 14272 7052 14300
rect 7190 14288 7196 14340
rect 7248 14328 7254 14340
rect 7668 14328 7696 14356
rect 7248 14300 7696 14328
rect 7248 14288 7254 14300
rect 8036 14272 8064 14359
rect 8202 14356 8208 14368
rect 8260 14356 8266 14408
rect 9214 14356 9220 14408
rect 9272 14396 9278 14408
rect 14090 14396 14096 14408
rect 9272 14368 14096 14396
rect 9272 14356 9278 14368
rect 14090 14356 14096 14368
rect 14148 14356 14154 14408
rect 14458 14356 14464 14408
rect 14516 14396 14522 14408
rect 14829 14399 14887 14405
rect 14829 14396 14841 14399
rect 14516 14368 14841 14396
rect 14516 14356 14522 14368
rect 14829 14365 14841 14368
rect 14875 14365 14887 14399
rect 14829 14359 14887 14365
rect 8941 14331 8999 14337
rect 8941 14328 8953 14331
rect 8128 14300 8953 14328
rect 8128 14272 8156 14300
rect 8941 14297 8953 14300
rect 8987 14297 8999 14331
rect 9122 14328 9128 14340
rect 9083 14300 9128 14328
rect 8941 14291 8999 14297
rect 9122 14288 9128 14300
rect 9180 14288 9186 14340
rect 10864 14331 10922 14337
rect 10864 14297 10876 14331
rect 10910 14328 10922 14331
rect 11238 14328 11244 14340
rect 10910 14300 11244 14328
rect 10910 14297 10922 14300
rect 10864 14291 10922 14297
rect 11238 14288 11244 14300
rect 11296 14288 11302 14340
rect 11330 14288 11336 14340
rect 11388 14328 11394 14340
rect 12250 14328 12256 14340
rect 11388 14300 12256 14328
rect 11388 14288 11394 14300
rect 12250 14288 12256 14300
rect 12308 14328 12314 14340
rect 14185 14331 14243 14337
rect 14185 14328 14197 14331
rect 12308 14300 14197 14328
rect 12308 14288 12314 14300
rect 14185 14297 14197 14300
rect 14231 14328 14243 14331
rect 14366 14328 14372 14340
rect 14231 14300 14372 14328
rect 14231 14297 14243 14300
rect 14185 14291 14243 14297
rect 14366 14288 14372 14300
rect 14424 14288 14430 14340
rect 14936 14328 14964 14436
rect 15028 14436 15384 14464
rect 15028 14405 15056 14436
rect 15378 14424 15384 14436
rect 15436 14424 15442 14476
rect 16114 14424 16120 14476
rect 16172 14424 16178 14476
rect 22370 14464 22376 14476
rect 22331 14436 22376 14464
rect 22370 14424 22376 14436
rect 22428 14424 22434 14476
rect 25774 14464 25780 14476
rect 25424 14436 25780 14464
rect 15013 14399 15071 14405
rect 15013 14365 15025 14399
rect 15059 14365 15071 14399
rect 15013 14359 15071 14365
rect 15105 14399 15163 14405
rect 15105 14365 15117 14399
rect 15151 14365 15163 14399
rect 15105 14359 15163 14365
rect 15197 14399 15255 14405
rect 15197 14365 15209 14399
rect 15243 14396 15255 14399
rect 15286 14396 15292 14408
rect 15243 14368 15292 14396
rect 15243 14365 15255 14368
rect 15197 14359 15255 14365
rect 15120 14328 15148 14359
rect 15286 14356 15292 14368
rect 15344 14356 15350 14408
rect 15841 14399 15899 14405
rect 15841 14396 15853 14399
rect 15396 14368 15853 14396
rect 14936 14300 15148 14328
rect 2409 14263 2467 14269
rect 2409 14229 2421 14263
rect 2455 14260 2467 14263
rect 2774 14260 2780 14272
rect 2455 14232 2780 14260
rect 2455 14229 2467 14232
rect 2409 14223 2467 14229
rect 2774 14220 2780 14232
rect 2832 14220 2838 14272
rect 5718 14260 5724 14272
rect 5679 14232 5724 14260
rect 5718 14220 5724 14232
rect 5776 14220 5782 14272
rect 7006 14220 7012 14272
rect 7064 14220 7070 14272
rect 8018 14220 8024 14272
rect 8076 14220 8082 14272
rect 8110 14220 8116 14272
rect 8168 14220 8174 14272
rect 8386 14260 8392 14272
rect 8347 14232 8392 14260
rect 8386 14220 8392 14232
rect 8444 14220 8450 14272
rect 12618 14220 12624 14272
rect 12676 14260 12682 14272
rect 12805 14263 12863 14269
rect 12805 14260 12817 14263
rect 12676 14232 12817 14260
rect 12676 14220 12682 14232
rect 12805 14229 12817 14232
rect 12851 14229 12863 14263
rect 13354 14260 13360 14272
rect 13315 14232 13360 14260
rect 12805 14223 12863 14229
rect 13354 14220 13360 14232
rect 13412 14220 13418 14272
rect 15396 14269 15424 14368
rect 15841 14365 15853 14368
rect 15887 14365 15899 14399
rect 15841 14359 15899 14365
rect 15930 14356 15936 14408
rect 15988 14396 15994 14408
rect 16132 14396 16160 14424
rect 16306 14399 16364 14405
rect 16306 14396 16318 14399
rect 15988 14368 16033 14396
rect 16132 14368 16318 14396
rect 15988 14356 15994 14368
rect 16306 14365 16318 14368
rect 16352 14365 16364 14399
rect 17126 14396 17132 14408
rect 17087 14368 17132 14396
rect 16306 14359 16364 14365
rect 17126 14356 17132 14368
rect 17184 14356 17190 14408
rect 17313 14399 17371 14405
rect 17313 14365 17325 14399
rect 17359 14396 17371 14399
rect 20162 14396 20168 14408
rect 17359 14368 20168 14396
rect 17359 14365 17371 14368
rect 17313 14359 17371 14365
rect 20162 14356 20168 14368
rect 20220 14356 20226 14408
rect 20714 14396 20720 14408
rect 20675 14368 20720 14396
rect 20714 14356 20720 14368
rect 20772 14356 20778 14408
rect 22465 14399 22523 14405
rect 22465 14365 22477 14399
rect 22511 14396 22523 14399
rect 23934 14396 23940 14408
rect 22511 14368 23940 14396
rect 22511 14365 22523 14368
rect 22465 14359 22523 14365
rect 23934 14356 23940 14368
rect 23992 14356 23998 14408
rect 25314 14396 25320 14408
rect 25275 14368 25320 14396
rect 25314 14356 25320 14368
rect 25372 14356 25378 14408
rect 25424 14405 25452 14436
rect 25774 14424 25780 14436
rect 25832 14424 25838 14476
rect 25409 14399 25467 14405
rect 25409 14365 25421 14399
rect 25455 14365 25467 14399
rect 25409 14359 25467 14365
rect 25498 14356 25504 14408
rect 25556 14396 25562 14408
rect 25685 14399 25743 14405
rect 25556 14368 25601 14396
rect 25556 14356 25562 14368
rect 25685 14365 25697 14399
rect 25731 14396 25743 14399
rect 25884 14396 25912 14504
rect 25731 14368 25912 14396
rect 25731 14365 25743 14368
rect 25685 14359 25743 14365
rect 15746 14288 15752 14340
rect 15804 14328 15810 14340
rect 16117 14331 16175 14337
rect 16117 14328 16129 14331
rect 15804 14300 16129 14328
rect 15804 14288 15810 14300
rect 16117 14297 16129 14300
rect 16163 14297 16175 14331
rect 16117 14291 16175 14297
rect 16209 14331 16267 14337
rect 16209 14297 16221 14331
rect 16255 14328 16267 14331
rect 26068 14328 26096 14572
rect 26789 14535 26847 14541
rect 26789 14501 26801 14535
rect 26835 14532 26847 14535
rect 27246 14532 27252 14544
rect 26835 14504 27252 14532
rect 26835 14501 26847 14504
rect 26789 14495 26847 14501
rect 27246 14492 27252 14504
rect 27304 14492 27310 14544
rect 28166 14532 28172 14544
rect 28092 14504 28172 14532
rect 27982 14356 27988 14408
rect 28040 14396 28046 14408
rect 28092 14405 28120 14504
rect 28166 14492 28172 14504
rect 28224 14492 28230 14544
rect 28828 14532 28856 14572
rect 28902 14560 28908 14612
rect 28960 14600 28966 14612
rect 28960 14572 34192 14600
rect 28960 14560 28966 14572
rect 29730 14532 29736 14544
rect 28828 14504 29736 14532
rect 29730 14492 29736 14504
rect 29788 14492 29794 14544
rect 29917 14535 29975 14541
rect 29917 14501 29929 14535
rect 29963 14532 29975 14535
rect 30006 14532 30012 14544
rect 29963 14504 30012 14532
rect 29963 14501 29975 14504
rect 29917 14495 29975 14501
rect 30006 14492 30012 14504
rect 30064 14492 30070 14544
rect 30469 14535 30527 14541
rect 30469 14501 30481 14535
rect 30515 14532 30527 14535
rect 30558 14532 30564 14544
rect 30515 14504 30564 14532
rect 30515 14501 30527 14504
rect 30469 14495 30527 14501
rect 30558 14492 30564 14504
rect 30616 14492 30622 14544
rect 30926 14532 30932 14544
rect 30887 14504 30932 14532
rect 30926 14492 30932 14504
rect 30984 14492 30990 14544
rect 32306 14532 32312 14544
rect 31726 14504 32312 14532
rect 31726 14464 31754 14504
rect 32306 14492 32312 14504
rect 32364 14492 32370 14544
rect 28184 14436 31754 14464
rect 28184 14405 28212 14436
rect 28077 14399 28135 14405
rect 28077 14396 28089 14399
rect 28040 14368 28089 14396
rect 28040 14356 28046 14368
rect 28077 14365 28089 14368
rect 28123 14365 28135 14399
rect 28077 14359 28135 14365
rect 28169 14399 28227 14405
rect 28169 14365 28181 14399
rect 28215 14365 28227 14399
rect 28169 14359 28227 14365
rect 28350 14356 28356 14408
rect 28408 14396 28414 14408
rect 28445 14399 28503 14405
rect 28445 14396 28457 14399
rect 28408 14368 28457 14396
rect 28408 14356 28414 14368
rect 28445 14365 28457 14368
rect 28491 14365 28503 14399
rect 28445 14359 28503 14365
rect 30558 14356 30564 14408
rect 30616 14396 30622 14408
rect 31570 14396 31576 14408
rect 30616 14368 31576 14396
rect 30616 14356 30622 14368
rect 31570 14356 31576 14368
rect 31628 14396 31634 14408
rect 31662 14396 31668 14408
rect 31628 14368 31668 14396
rect 31628 14356 31634 14368
rect 31662 14356 31668 14368
rect 31720 14356 31726 14408
rect 31941 14399 31999 14405
rect 31941 14365 31953 14399
rect 31987 14396 31999 14399
rect 33134 14396 33140 14408
rect 31987 14368 33140 14396
rect 31987 14365 31999 14368
rect 31941 14359 31999 14365
rect 16255 14300 26096 14328
rect 16255 14297 16267 14300
rect 16209 14291 16267 14297
rect 15381 14263 15439 14269
rect 15381 14229 15393 14263
rect 15427 14229 15439 14263
rect 16132 14260 16160 14291
rect 26234 14288 26240 14340
rect 26292 14328 26298 14340
rect 27706 14328 27712 14340
rect 26292 14300 27712 14328
rect 26292 14288 26298 14300
rect 27706 14288 27712 14300
rect 27764 14288 27770 14340
rect 28261 14331 28319 14337
rect 28261 14297 28273 14331
rect 28307 14328 28319 14331
rect 28626 14328 28632 14340
rect 28307 14300 28632 14328
rect 28307 14297 28319 14300
rect 28261 14291 28319 14297
rect 28626 14288 28632 14300
rect 28684 14288 28690 14340
rect 29086 14288 29092 14340
rect 29144 14328 29150 14340
rect 29549 14331 29607 14337
rect 29549 14328 29561 14331
rect 29144 14300 29561 14328
rect 29144 14288 29150 14300
rect 29549 14297 29561 14300
rect 29595 14297 29607 14331
rect 29730 14328 29736 14340
rect 29691 14300 29736 14328
rect 29549 14291 29607 14297
rect 29730 14288 29736 14300
rect 29788 14328 29794 14340
rect 31018 14328 31024 14340
rect 29788 14300 31024 14328
rect 29788 14288 29794 14300
rect 31018 14288 31024 14300
rect 31076 14288 31082 14340
rect 31113 14331 31171 14337
rect 31113 14297 31125 14331
rect 31159 14297 31171 14331
rect 31113 14291 31171 14297
rect 16390 14260 16396 14272
rect 16132 14232 16396 14260
rect 15381 14223 15439 14229
rect 16390 14220 16396 14232
rect 16448 14220 16454 14272
rect 16485 14263 16543 14269
rect 16485 14229 16497 14263
rect 16531 14260 16543 14263
rect 16666 14260 16672 14272
rect 16531 14232 16672 14260
rect 16531 14229 16543 14232
rect 16485 14223 16543 14229
rect 16666 14220 16672 14232
rect 16724 14220 16730 14272
rect 17126 14220 17132 14272
rect 17184 14260 17190 14272
rect 17497 14263 17555 14269
rect 17497 14260 17509 14263
rect 17184 14232 17509 14260
rect 17184 14220 17190 14232
rect 17497 14229 17509 14232
rect 17543 14229 17555 14263
rect 17497 14223 17555 14229
rect 18782 14220 18788 14272
rect 18840 14260 18846 14272
rect 20257 14263 20315 14269
rect 20257 14260 20269 14263
rect 18840 14232 20269 14260
rect 18840 14220 18846 14232
rect 20257 14229 20269 14232
rect 20303 14260 20315 14263
rect 20714 14260 20720 14272
rect 20303 14232 20720 14260
rect 20303 14229 20315 14232
rect 20257 14223 20315 14229
rect 20714 14220 20720 14232
rect 20772 14220 20778 14272
rect 20901 14263 20959 14269
rect 20901 14229 20913 14263
rect 20947 14260 20959 14263
rect 22922 14260 22928 14272
rect 20947 14232 22928 14260
rect 20947 14229 20959 14232
rect 20901 14223 20959 14229
rect 22922 14220 22928 14232
rect 22980 14220 22986 14272
rect 24581 14263 24639 14269
rect 24581 14229 24593 14263
rect 24627 14260 24639 14263
rect 24946 14260 24952 14272
rect 24627 14232 24952 14260
rect 24627 14229 24639 14232
rect 24581 14223 24639 14229
rect 24946 14220 24952 14232
rect 25004 14220 25010 14272
rect 27338 14220 27344 14272
rect 27396 14260 27402 14272
rect 27893 14263 27951 14269
rect 27893 14260 27905 14263
rect 27396 14232 27905 14260
rect 27396 14220 27402 14232
rect 27893 14229 27905 14232
rect 27939 14229 27951 14263
rect 27893 14223 27951 14229
rect 28997 14263 29055 14269
rect 28997 14229 29009 14263
rect 29043 14260 29055 14263
rect 29638 14260 29644 14272
rect 29043 14232 29644 14260
rect 29043 14229 29055 14232
rect 28997 14223 29055 14229
rect 29638 14220 29644 14232
rect 29696 14220 29702 14272
rect 31128 14260 31156 14291
rect 31478 14260 31484 14272
rect 31128 14232 31484 14260
rect 31478 14220 31484 14232
rect 31536 14260 31542 14272
rect 31956 14260 31984 14359
rect 33134 14356 33140 14368
rect 33192 14356 33198 14408
rect 34164 14337 34192 14572
rect 37642 14492 37648 14544
rect 37700 14532 37706 14544
rect 37918 14532 37924 14544
rect 37700 14504 37924 14532
rect 37700 14492 37706 14504
rect 37918 14492 37924 14504
rect 37976 14492 37982 14544
rect 34238 14356 34244 14408
rect 34296 14396 34302 14408
rect 37274 14396 37280 14408
rect 34296 14368 37280 14396
rect 34296 14356 34302 14368
rect 37274 14356 37280 14368
rect 37332 14356 37338 14408
rect 37458 14356 37464 14408
rect 37516 14396 37522 14408
rect 37939 14405 37967 14492
rect 37645 14399 37703 14405
rect 37924 14399 37982 14405
rect 37645 14396 37657 14399
rect 37516 14368 37657 14396
rect 37516 14356 37522 14368
rect 37645 14365 37657 14368
rect 37691 14365 37703 14399
rect 37645 14359 37703 14365
rect 37824 14393 37882 14399
rect 37824 14359 37836 14393
rect 37870 14359 37882 14393
rect 37924 14365 37936 14399
rect 37970 14365 37982 14399
rect 37924 14359 37982 14365
rect 37824 14353 37882 14359
rect 38010 14356 38016 14408
rect 38068 14405 38074 14408
rect 38068 14399 38091 14405
rect 38079 14365 38091 14399
rect 38930 14396 38936 14408
rect 38891 14368 38936 14396
rect 38068 14359 38091 14365
rect 38068 14356 38074 14359
rect 38930 14356 38936 14368
rect 38988 14356 38994 14408
rect 68094 14396 68100 14408
rect 68055 14368 68100 14396
rect 68094 14356 68100 14368
rect 68152 14356 68158 14408
rect 34149 14331 34207 14337
rect 34149 14297 34161 14331
rect 34195 14328 34207 14331
rect 35894 14328 35900 14340
rect 34195 14300 35900 14328
rect 34195 14297 34207 14300
rect 34149 14291 34207 14297
rect 35894 14288 35900 14300
rect 35952 14328 35958 14340
rect 36814 14328 36820 14340
rect 35952 14300 36820 14328
rect 35952 14288 35958 14300
rect 36814 14288 36820 14300
rect 36872 14288 36878 14340
rect 32950 14260 32956 14272
rect 31536 14232 31984 14260
rect 32911 14232 32956 14260
rect 31536 14220 31542 14232
rect 32950 14220 32956 14232
rect 33008 14220 33014 14272
rect 34422 14220 34428 14272
rect 34480 14260 34486 14272
rect 35529 14263 35587 14269
rect 35529 14260 35541 14263
rect 34480 14232 35541 14260
rect 34480 14220 34486 14232
rect 35529 14229 35541 14232
rect 35575 14260 35587 14263
rect 36630 14260 36636 14272
rect 35575 14232 36636 14260
rect 35575 14229 35587 14232
rect 35529 14223 35587 14229
rect 36630 14220 36636 14232
rect 36688 14220 36694 14272
rect 37734 14220 37740 14272
rect 37792 14260 37798 14272
rect 37839 14260 37867 14353
rect 38749 14331 38807 14337
rect 38749 14297 38761 14331
rect 38795 14328 38807 14331
rect 38838 14328 38844 14340
rect 38795 14300 38844 14328
rect 38795 14297 38807 14300
rect 38749 14291 38807 14297
rect 38838 14288 38844 14300
rect 38896 14288 38902 14340
rect 38286 14260 38292 14272
rect 37792 14232 37867 14260
rect 38247 14232 38292 14260
rect 37792 14220 37798 14232
rect 38286 14220 38292 14232
rect 38344 14220 38350 14272
rect 39114 14260 39120 14272
rect 39075 14232 39120 14260
rect 39114 14220 39120 14232
rect 39172 14220 39178 14272
rect 1104 14170 68816 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 68816 14170
rect 1104 14096 68816 14118
rect 4062 14056 4068 14068
rect 4023 14028 4068 14056
rect 4062 14016 4068 14028
rect 4120 14016 4126 14068
rect 6638 14016 6644 14068
rect 6696 14056 6702 14068
rect 6733 14059 6791 14065
rect 6733 14056 6745 14059
rect 6696 14028 6745 14056
rect 6696 14016 6702 14028
rect 6733 14025 6745 14028
rect 6779 14056 6791 14059
rect 7282 14056 7288 14068
rect 6779 14028 7288 14056
rect 6779 14025 6791 14028
rect 6733 14019 6791 14025
rect 7282 14016 7288 14028
rect 7340 14056 7346 14068
rect 8110 14056 8116 14068
rect 7340 14028 8116 14056
rect 7340 14016 7346 14028
rect 8110 14016 8116 14028
rect 8168 14016 8174 14068
rect 9122 14016 9128 14068
rect 9180 14056 9186 14068
rect 10781 14059 10839 14065
rect 10781 14056 10793 14059
rect 9180 14028 10793 14056
rect 9180 14016 9186 14028
rect 10781 14025 10793 14028
rect 10827 14056 10839 14059
rect 11146 14056 11152 14068
rect 10827 14028 11152 14056
rect 10827 14025 10839 14028
rect 10781 14019 10839 14025
rect 11146 14016 11152 14028
rect 11204 14016 11210 14068
rect 11238 14016 11244 14068
rect 11296 14056 11302 14068
rect 11517 14059 11575 14065
rect 11517 14056 11529 14059
rect 11296 14028 11529 14056
rect 11296 14016 11302 14028
rect 11517 14025 11529 14028
rect 11563 14025 11575 14059
rect 11517 14019 11575 14025
rect 13909 14059 13967 14065
rect 13909 14025 13921 14059
rect 13955 14056 13967 14059
rect 14182 14056 14188 14068
rect 13955 14028 14188 14056
rect 13955 14025 13967 14028
rect 13909 14019 13967 14025
rect 14182 14016 14188 14028
rect 14240 14016 14246 14068
rect 16868 14028 20024 14056
rect 3142 13988 3148 14000
rect 2700 13960 3148 13988
rect 2700 13929 2728 13960
rect 3142 13948 3148 13960
rect 3200 13948 3206 14000
rect 4614 13988 4620 14000
rect 4527 13960 4620 13988
rect 2685 13923 2743 13929
rect 2685 13889 2697 13923
rect 2731 13889 2743 13923
rect 2685 13883 2743 13889
rect 2774 13880 2780 13932
rect 2832 13920 2838 13932
rect 4540 13929 4568 13960
rect 4614 13948 4620 13960
rect 4672 13988 4678 14000
rect 7193 13991 7251 13997
rect 7193 13988 7205 13991
rect 4672 13960 7205 13988
rect 4672 13948 4678 13960
rect 7193 13957 7205 13960
rect 7239 13957 7251 13991
rect 7193 13951 7251 13957
rect 8386 13948 8392 14000
rect 8444 13988 8450 14000
rect 9646 13991 9704 13997
rect 9646 13988 9658 13991
rect 8444 13960 9658 13988
rect 8444 13948 8450 13960
rect 9646 13957 9658 13960
rect 9692 13957 9704 13991
rect 13262 13988 13268 14000
rect 9646 13951 9704 13957
rect 12544 13960 13268 13988
rect 2941 13923 2999 13929
rect 2941 13920 2953 13923
rect 2832 13892 2953 13920
rect 2832 13880 2838 13892
rect 2941 13889 2953 13892
rect 2987 13889 2999 13923
rect 2941 13883 2999 13889
rect 4525 13923 4583 13929
rect 4525 13889 4537 13923
rect 4571 13889 4583 13923
rect 4798 13920 4804 13932
rect 4759 13892 4804 13920
rect 4525 13883 4583 13889
rect 4798 13880 4804 13892
rect 4856 13880 4862 13932
rect 6457 13923 6515 13929
rect 6457 13889 6469 13923
rect 6503 13889 6515 13923
rect 6457 13883 6515 13889
rect 6549 13923 6607 13929
rect 6549 13889 6561 13923
rect 6595 13920 6607 13923
rect 6822 13920 6828 13932
rect 6595 13892 6828 13920
rect 6595 13889 6607 13892
rect 6549 13883 6607 13889
rect 1762 13812 1768 13864
rect 1820 13852 1826 13864
rect 1949 13855 2007 13861
rect 1949 13852 1961 13855
rect 1820 13824 1961 13852
rect 1820 13812 1826 13824
rect 1949 13821 1961 13824
rect 1995 13821 2007 13855
rect 1949 13815 2007 13821
rect 2225 13855 2283 13861
rect 2225 13821 2237 13855
rect 2271 13852 2283 13855
rect 2271 13824 2728 13852
rect 2271 13821 2283 13824
rect 2225 13815 2283 13821
rect 2700 13716 2728 13824
rect 6472 13784 6500 13883
rect 6822 13880 6828 13892
rect 6880 13880 6886 13932
rect 7377 13923 7435 13929
rect 7377 13889 7389 13923
rect 7423 13920 7435 13923
rect 7742 13920 7748 13932
rect 7423 13892 7748 13920
rect 7423 13889 7435 13892
rect 7377 13883 7435 13889
rect 7742 13880 7748 13892
rect 7800 13920 7806 13932
rect 8665 13923 8723 13929
rect 8665 13920 8677 13923
rect 7800 13892 8677 13920
rect 7800 13880 7806 13892
rect 8665 13889 8677 13892
rect 8711 13889 8723 13923
rect 8665 13883 8723 13889
rect 9030 13880 9036 13932
rect 9088 13920 9094 13932
rect 9401 13923 9459 13929
rect 9401 13920 9413 13923
rect 9088 13892 9413 13920
rect 9088 13880 9094 13892
rect 9401 13889 9413 13892
rect 9447 13889 9459 13923
rect 11790 13920 11796 13932
rect 9401 13883 9459 13889
rect 9508 13892 11652 13920
rect 11751 13892 11796 13920
rect 7561 13855 7619 13861
rect 7561 13821 7573 13855
rect 7607 13821 7619 13855
rect 7561 13815 7619 13821
rect 8941 13855 8999 13861
rect 8941 13821 8953 13855
rect 8987 13852 8999 13855
rect 9508 13852 9536 13892
rect 8987 13824 9536 13852
rect 8987 13821 8999 13824
rect 8941 13815 8999 13821
rect 7576 13784 7604 13815
rect 8294 13784 8300 13796
rect 6472 13756 8300 13784
rect 3050 13716 3056 13728
rect 2700 13688 3056 13716
rect 3050 13676 3056 13688
rect 3108 13676 3114 13728
rect 5902 13676 5908 13728
rect 5960 13716 5966 13728
rect 6472 13716 6500 13756
rect 8294 13744 8300 13756
rect 8352 13784 8358 13796
rect 9030 13784 9036 13796
rect 8352 13756 9036 13784
rect 8352 13744 8358 13756
rect 9030 13744 9036 13756
rect 9088 13744 9094 13796
rect 11624 13784 11652 13892
rect 11790 13880 11796 13892
rect 11848 13880 11854 13932
rect 11885 13923 11943 13929
rect 11885 13889 11897 13923
rect 11931 13889 11943 13923
rect 11885 13883 11943 13889
rect 11900 13852 11928 13883
rect 11974 13880 11980 13932
rect 12032 13920 12038 13932
rect 12161 13923 12219 13929
rect 12032 13892 12077 13920
rect 12032 13880 12038 13892
rect 12161 13889 12173 13923
rect 12207 13920 12219 13923
rect 12544 13920 12572 13960
rect 13262 13948 13268 13960
rect 13320 13948 13326 14000
rect 14829 13991 14887 13997
rect 14829 13957 14841 13991
rect 14875 13988 14887 13991
rect 15933 13991 15991 13997
rect 14875 13960 15884 13988
rect 14875 13957 14887 13960
rect 14829 13951 14887 13957
rect 12207 13892 12572 13920
rect 12207 13889 12219 13892
rect 12161 13883 12219 13889
rect 12618 13880 12624 13932
rect 12676 13920 12682 13932
rect 13081 13923 13139 13929
rect 13081 13920 13093 13923
rect 12676 13892 13093 13920
rect 12676 13880 12682 13892
rect 13081 13889 13093 13892
rect 13127 13889 13139 13923
rect 14090 13920 14096 13932
rect 14051 13892 14096 13920
rect 13081 13883 13139 13889
rect 14090 13880 14096 13892
rect 14148 13920 14154 13932
rect 14645 13923 14703 13929
rect 14645 13920 14657 13923
rect 14148 13892 14657 13920
rect 14148 13880 14154 13892
rect 14645 13889 14657 13892
rect 14691 13889 14703 13923
rect 15562 13920 15568 13932
rect 15523 13892 15568 13920
rect 14645 13883 14703 13889
rect 15562 13880 15568 13892
rect 15620 13880 15626 13932
rect 15749 13923 15807 13929
rect 15749 13889 15761 13923
rect 15795 13889 15807 13923
rect 15856 13920 15884 13960
rect 15933 13957 15945 13991
rect 15979 13988 15991 13991
rect 16114 13988 16120 14000
rect 15979 13960 16120 13988
rect 15979 13957 15991 13960
rect 15933 13951 15991 13957
rect 16114 13948 16120 13960
rect 16172 13948 16178 14000
rect 16666 13920 16672 13932
rect 15856 13892 16528 13920
rect 16627 13892 16672 13920
rect 15749 13883 15807 13889
rect 12710 13852 12716 13864
rect 11900 13824 12716 13852
rect 12710 13812 12716 13824
rect 12768 13812 12774 13864
rect 13630 13852 13636 13864
rect 13280 13824 13636 13852
rect 11882 13784 11888 13796
rect 11624 13756 11888 13784
rect 11882 13744 11888 13756
rect 11940 13744 11946 13796
rect 13280 13793 13308 13824
rect 13630 13812 13636 13824
rect 13688 13812 13694 13864
rect 15194 13812 15200 13864
rect 15252 13852 15258 13864
rect 15764 13852 15792 13883
rect 15252 13824 15792 13852
rect 15252 13812 15258 13824
rect 13265 13787 13323 13793
rect 13265 13753 13277 13787
rect 13311 13753 13323 13787
rect 16500 13784 16528 13892
rect 16666 13880 16672 13892
rect 16724 13880 16730 13932
rect 16868 13929 16896 14028
rect 19996 13988 20024 14028
rect 20162 14016 20168 14068
rect 20220 14056 20226 14068
rect 24029 14059 24087 14065
rect 24029 14056 24041 14059
rect 20220 14028 24041 14056
rect 20220 14016 20226 14028
rect 24029 14025 24041 14028
rect 24075 14025 24087 14059
rect 32490 14056 32496 14068
rect 24029 14019 24087 14025
rect 27908 14028 32496 14056
rect 23382 13988 23388 14000
rect 18064 13960 19932 13988
rect 19996 13960 23388 13988
rect 18064 13929 18092 13960
rect 16853 13923 16911 13929
rect 16853 13889 16865 13923
rect 16899 13889 16911 13923
rect 16853 13883 16911 13889
rect 18049 13923 18107 13929
rect 18049 13889 18061 13923
rect 18095 13889 18107 13923
rect 18049 13883 18107 13889
rect 18138 13880 18144 13932
rect 18196 13920 18202 13932
rect 19904 13929 19932 13960
rect 23382 13948 23388 13960
rect 23440 13948 23446 14000
rect 25314 13948 25320 14000
rect 25372 13988 25378 14000
rect 25961 13991 26019 13997
rect 25961 13988 25973 13991
rect 25372 13960 25973 13988
rect 25372 13948 25378 13960
rect 25961 13957 25973 13960
rect 26007 13988 26019 13991
rect 27908 13988 27936 14028
rect 32490 14016 32496 14028
rect 32548 14016 32554 14068
rect 32766 14016 32772 14068
rect 32824 14056 32830 14068
rect 33689 14059 33747 14065
rect 32824 14028 33088 14056
rect 32824 14016 32830 14028
rect 26007 13960 27936 13988
rect 28077 13991 28135 13997
rect 26007 13957 26019 13960
rect 25961 13951 26019 13957
rect 28077 13957 28089 13991
rect 28123 13988 28135 13991
rect 30558 13988 30564 14000
rect 28123 13960 30564 13988
rect 28123 13957 28135 13960
rect 28077 13951 28135 13957
rect 30558 13948 30564 13960
rect 30616 13948 30622 14000
rect 31205 13991 31263 13997
rect 31205 13957 31217 13991
rect 31251 13988 31263 13991
rect 31251 13960 31524 13988
rect 31251 13957 31263 13960
rect 31205 13951 31263 13957
rect 18305 13923 18363 13929
rect 18305 13920 18317 13923
rect 18196 13892 18317 13920
rect 18196 13880 18202 13892
rect 18305 13889 18317 13892
rect 18351 13889 18363 13923
rect 18305 13883 18363 13889
rect 19889 13923 19947 13929
rect 19889 13889 19901 13923
rect 19935 13920 19947 13923
rect 19978 13920 19984 13932
rect 19935 13892 19984 13920
rect 19935 13889 19947 13892
rect 19889 13883 19947 13889
rect 19978 13880 19984 13892
rect 20036 13880 20042 13932
rect 20162 13929 20168 13932
rect 20156 13883 20168 13929
rect 20220 13920 20226 13932
rect 22278 13920 22284 13932
rect 20220 13892 20256 13920
rect 22239 13892 22284 13920
rect 20162 13880 20168 13883
rect 20220 13880 20226 13892
rect 22278 13880 22284 13892
rect 22336 13920 22342 13932
rect 22646 13920 22652 13932
rect 22336 13892 22652 13920
rect 22336 13880 22342 13892
rect 22646 13880 22652 13892
rect 22704 13920 22710 13932
rect 22925 13923 22983 13929
rect 22925 13920 22937 13923
rect 22704 13892 22937 13920
rect 22704 13880 22710 13892
rect 22925 13889 22937 13892
rect 22971 13889 22983 13923
rect 23566 13920 23572 13932
rect 23527 13892 23572 13920
rect 22925 13883 22983 13889
rect 23566 13880 23572 13892
rect 23624 13880 23630 13932
rect 23845 13923 23903 13929
rect 23845 13889 23857 13923
rect 23891 13920 23903 13923
rect 24486 13920 24492 13932
rect 23891 13892 24492 13920
rect 23891 13889 23903 13892
rect 23845 13883 23903 13889
rect 24486 13880 24492 13892
rect 24544 13880 24550 13932
rect 24946 13880 24952 13932
rect 25004 13920 25010 13932
rect 25041 13923 25099 13929
rect 25041 13920 25053 13923
rect 25004 13892 25053 13920
rect 25004 13880 25010 13892
rect 25041 13889 25053 13892
rect 25087 13889 25099 13923
rect 25041 13883 25099 13889
rect 25133 13923 25191 13929
rect 25133 13889 25145 13923
rect 25179 13889 25191 13923
rect 25133 13883 25191 13889
rect 16574 13812 16580 13864
rect 16632 13852 16638 13864
rect 22465 13855 22523 13861
rect 16632 13824 17080 13852
rect 16632 13812 16638 13824
rect 17052 13793 17080 13824
rect 22465 13821 22477 13855
rect 22511 13852 22523 13855
rect 23658 13852 23664 13864
rect 22511 13824 23520 13852
rect 23619 13824 23664 13852
rect 22511 13821 22523 13824
rect 22465 13815 22523 13821
rect 17037 13787 17095 13793
rect 16500 13756 16988 13784
rect 13265 13747 13323 13753
rect 5960 13688 6500 13716
rect 5960 13676 5966 13688
rect 7834 13676 7840 13728
rect 7892 13716 7898 13728
rect 11790 13716 11796 13728
rect 7892 13688 11796 13716
rect 7892 13676 7898 13688
rect 11790 13676 11796 13688
rect 11848 13676 11854 13728
rect 16666 13716 16672 13728
rect 16627 13688 16672 13716
rect 16666 13676 16672 13688
rect 16724 13676 16730 13728
rect 16960 13716 16988 13756
rect 17037 13753 17049 13787
rect 17083 13753 17095 13787
rect 23492 13784 23520 13824
rect 23658 13812 23664 13824
rect 23716 13812 23722 13864
rect 24964 13852 24992 13880
rect 23768 13824 24992 13852
rect 25148 13852 25176 13883
rect 25222 13880 25228 13932
rect 25280 13920 25286 13932
rect 25409 13923 25467 13929
rect 25280 13892 25325 13920
rect 25280 13880 25286 13892
rect 25409 13889 25421 13923
rect 25455 13889 25467 13923
rect 27062 13920 27068 13932
rect 27023 13892 27068 13920
rect 25409 13883 25467 13889
rect 25148 13824 25268 13852
rect 23768 13784 23796 13824
rect 25240 13784 25268 13824
rect 25314 13812 25320 13864
rect 25372 13852 25378 13864
rect 25424 13852 25452 13883
rect 27062 13880 27068 13892
rect 27120 13880 27126 13932
rect 27982 13920 27988 13932
rect 27943 13892 27988 13920
rect 27982 13880 27988 13892
rect 28040 13880 28046 13932
rect 28169 13923 28227 13929
rect 28169 13889 28181 13923
rect 28215 13889 28227 13923
rect 28169 13883 28227 13889
rect 25372 13824 25452 13852
rect 25372 13812 25378 13824
rect 27890 13812 27896 13864
rect 27948 13852 27954 13864
rect 28184 13852 28212 13883
rect 28258 13880 28264 13932
rect 28316 13920 28322 13932
rect 28353 13923 28411 13929
rect 28353 13920 28365 13923
rect 28316 13892 28365 13920
rect 28316 13880 28322 13892
rect 28353 13889 28365 13892
rect 28399 13889 28411 13923
rect 30576 13920 30604 13948
rect 31389 13923 31447 13929
rect 31389 13920 31401 13923
rect 30576 13892 31401 13920
rect 28353 13883 28411 13889
rect 31389 13889 31401 13892
rect 31435 13889 31447 13923
rect 31496 13920 31524 13960
rect 32122 13920 32128 13932
rect 31496 13892 32128 13920
rect 31389 13883 31447 13889
rect 32122 13880 32128 13892
rect 32180 13880 32186 13932
rect 33060 13929 33088 14028
rect 33689 14025 33701 14059
rect 33735 14056 33747 14059
rect 34514 14056 34520 14068
rect 33735 14028 34520 14056
rect 33735 14025 33747 14028
rect 33689 14019 33747 14025
rect 34514 14016 34520 14028
rect 34572 14016 34578 14068
rect 35253 14059 35311 14065
rect 35253 14056 35265 14059
rect 34624 14028 35265 14056
rect 33134 13948 33140 14000
rect 33192 13988 33198 14000
rect 33781 13991 33839 13997
rect 33781 13988 33793 13991
rect 33192 13960 33793 13988
rect 33192 13948 33198 13960
rect 33781 13957 33793 13960
rect 33827 13988 33839 13991
rect 34238 13988 34244 14000
rect 33827 13960 34244 13988
rect 33827 13957 33839 13960
rect 33781 13951 33839 13957
rect 34238 13948 34244 13960
rect 34296 13948 34302 14000
rect 34624 13997 34652 14028
rect 35253 14025 35265 14028
rect 35299 14056 35311 14059
rect 36446 14056 36452 14068
rect 35299 14028 36452 14056
rect 35299 14025 35311 14028
rect 35253 14019 35311 14025
rect 36446 14016 36452 14028
rect 36504 14016 36510 14068
rect 37734 14056 37740 14068
rect 37695 14028 37740 14056
rect 37734 14016 37740 14028
rect 37792 14016 37798 14068
rect 38933 14059 38991 14065
rect 38933 14056 38945 14059
rect 37844 14028 38945 14056
rect 34609 13991 34667 13997
rect 34609 13957 34621 13991
rect 34655 13957 34667 13991
rect 34609 13951 34667 13957
rect 36722 13948 36728 14000
rect 36780 13988 36786 14000
rect 37553 13991 37611 13997
rect 37553 13988 37565 13991
rect 36780 13960 37565 13988
rect 36780 13948 36786 13960
rect 37553 13957 37565 13960
rect 37599 13988 37611 13991
rect 37844 13988 37872 14028
rect 38933 14025 38945 14028
rect 38979 14025 38991 14059
rect 38933 14019 38991 14025
rect 37599 13960 37872 13988
rect 37599 13957 37611 13960
rect 37553 13951 37611 13957
rect 38286 13948 38292 14000
rect 38344 13988 38350 14000
rect 40046 13991 40104 13997
rect 40046 13988 40058 13991
rect 38344 13960 40058 13988
rect 38344 13948 38350 13960
rect 40046 13957 40058 13960
rect 40092 13957 40104 13991
rect 40046 13951 40104 13957
rect 32631 13923 32689 13929
rect 32631 13920 32643 13923
rect 32232 13892 32643 13920
rect 28626 13852 28632 13864
rect 27948 13824 28632 13852
rect 27948 13812 27954 13824
rect 28626 13812 28632 13824
rect 28684 13852 28690 13864
rect 28813 13855 28871 13861
rect 28813 13852 28825 13855
rect 28684 13824 28825 13852
rect 28684 13812 28690 13824
rect 28813 13821 28825 13824
rect 28859 13821 28871 13855
rect 28813 13815 28871 13821
rect 29089 13855 29147 13861
rect 29089 13821 29101 13855
rect 29135 13852 29147 13855
rect 29178 13852 29184 13864
rect 29135 13824 29184 13852
rect 29135 13821 29147 13824
rect 29089 13815 29147 13821
rect 29178 13812 29184 13824
rect 29236 13812 29242 13864
rect 29638 13812 29644 13864
rect 29696 13852 29702 13864
rect 30653 13855 30711 13861
rect 30653 13852 30665 13855
rect 29696 13824 30665 13852
rect 29696 13812 29702 13824
rect 30653 13821 30665 13824
rect 30699 13852 30711 13855
rect 32232 13852 32260 13892
rect 32631 13889 32643 13892
rect 32677 13889 32689 13923
rect 32631 13883 32689 13889
rect 32766 13923 32824 13929
rect 32766 13889 32778 13923
rect 32812 13889 32824 13923
rect 32766 13883 32824 13889
rect 32882 13923 32940 13929
rect 32882 13889 32894 13923
rect 32928 13920 32940 13923
rect 33045 13923 33103 13929
rect 32928 13892 32996 13920
rect 32928 13889 32940 13892
rect 32882 13883 32940 13889
rect 30699 13824 32260 13852
rect 32781 13852 32809 13883
rect 32781 13824 32904 13852
rect 30699 13821 30711 13824
rect 30653 13815 30711 13821
rect 32876 13796 32904 13824
rect 25498 13784 25504 13796
rect 23492 13756 23796 13784
rect 23860 13756 24900 13784
rect 25240 13756 25504 13784
rect 17037 13747 17095 13753
rect 17494 13716 17500 13728
rect 16960 13688 17500 13716
rect 17494 13676 17500 13688
rect 17552 13676 17558 13728
rect 19426 13716 19432 13728
rect 19339 13688 19432 13716
rect 19426 13676 19432 13688
rect 19484 13716 19490 13728
rect 20254 13716 20260 13728
rect 19484 13688 20260 13716
rect 19484 13676 19490 13688
rect 20254 13676 20260 13688
rect 20312 13676 20318 13728
rect 21266 13716 21272 13728
rect 21227 13688 21272 13716
rect 21266 13676 21272 13688
rect 21324 13676 21330 13728
rect 23860 13725 23888 13756
rect 23845 13719 23903 13725
rect 23845 13685 23857 13719
rect 23891 13685 23903 13719
rect 24762 13716 24768 13728
rect 24723 13688 24768 13716
rect 23845 13679 23903 13685
rect 24762 13676 24768 13688
rect 24820 13676 24826 13728
rect 24872 13716 24900 13756
rect 25498 13744 25504 13756
rect 25556 13744 25562 13796
rect 25774 13744 25780 13796
rect 25832 13784 25838 13796
rect 27801 13787 27859 13793
rect 27801 13784 27813 13787
rect 25832 13756 27813 13784
rect 25832 13744 25838 13756
rect 27801 13753 27813 13756
rect 27847 13753 27859 13787
rect 27801 13747 27859 13753
rect 31573 13787 31631 13793
rect 31573 13753 31585 13787
rect 31619 13784 31631 13787
rect 31619 13756 32740 13784
rect 31619 13753 31631 13756
rect 31573 13747 31631 13753
rect 28074 13716 28080 13728
rect 24872 13688 28080 13716
rect 28074 13676 28080 13688
rect 28132 13676 28138 13728
rect 28994 13676 29000 13728
rect 29052 13716 29058 13728
rect 29822 13716 29828 13728
rect 29052 13688 29828 13716
rect 29052 13676 29058 13688
rect 29822 13676 29828 13688
rect 29880 13676 29886 13728
rect 32398 13716 32404 13728
rect 32359 13688 32404 13716
rect 32398 13676 32404 13688
rect 32456 13676 32462 13728
rect 32712 13716 32740 13756
rect 32858 13744 32864 13796
rect 32916 13744 32922 13796
rect 32968 13716 32996 13892
rect 33045 13889 33057 13923
rect 33091 13889 33103 13923
rect 33045 13883 33103 13889
rect 34793 13923 34851 13929
rect 34793 13889 34805 13923
rect 34839 13920 34851 13923
rect 35894 13920 35900 13932
rect 34839 13892 35900 13920
rect 34839 13889 34851 13892
rect 34793 13883 34851 13889
rect 35894 13880 35900 13892
rect 35952 13880 35958 13932
rect 35986 13880 35992 13932
rect 36044 13920 36050 13932
rect 36366 13923 36424 13929
rect 36366 13920 36378 13923
rect 36044 13892 36378 13920
rect 36044 13880 36050 13892
rect 36366 13889 36378 13892
rect 36412 13889 36424 13923
rect 36630 13920 36636 13932
rect 36591 13892 36636 13920
rect 36366 13883 36424 13889
rect 36630 13880 36636 13892
rect 36688 13880 36694 13932
rect 37366 13920 37372 13932
rect 37327 13892 37372 13920
rect 37366 13880 37372 13892
rect 37424 13880 37430 13932
rect 40313 13923 40371 13929
rect 40313 13889 40325 13923
rect 40359 13920 40371 13923
rect 41230 13920 41236 13932
rect 40359 13892 41236 13920
rect 40359 13889 40371 13892
rect 40313 13883 40371 13889
rect 41230 13880 41236 13892
rect 41288 13880 41294 13932
rect 34425 13855 34483 13861
rect 34425 13821 34437 13855
rect 34471 13852 34483 13855
rect 35526 13852 35532 13864
rect 34471 13824 35532 13852
rect 34471 13821 34483 13824
rect 34425 13815 34483 13821
rect 35526 13812 35532 13824
rect 35584 13812 35590 13864
rect 32712 13688 32996 13716
rect 33042 13676 33048 13728
rect 33100 13716 33106 13728
rect 37826 13716 37832 13728
rect 33100 13688 37832 13716
rect 33100 13676 33106 13688
rect 37826 13676 37832 13688
rect 37884 13676 37890 13728
rect 38010 13676 38016 13728
rect 38068 13716 38074 13728
rect 39114 13716 39120 13728
rect 38068 13688 39120 13716
rect 38068 13676 38074 13688
rect 39114 13676 39120 13688
rect 39172 13676 39178 13728
rect 1104 13626 68816 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 65654 13626
rect 65706 13574 65718 13626
rect 65770 13574 65782 13626
rect 65834 13574 65846 13626
rect 65898 13574 65910 13626
rect 65962 13574 68816 13626
rect 1104 13552 68816 13574
rect 2866 13472 2872 13524
rect 2924 13512 2930 13524
rect 2961 13515 3019 13521
rect 2961 13512 2973 13515
rect 2924 13484 2973 13512
rect 2924 13472 2930 13484
rect 2961 13481 2973 13484
rect 3007 13512 3019 13515
rect 3050 13512 3056 13524
rect 3007 13484 3056 13512
rect 3007 13481 3019 13484
rect 2961 13475 3019 13481
rect 3050 13472 3056 13484
rect 3108 13472 3114 13524
rect 4617 13515 4675 13521
rect 4617 13481 4629 13515
rect 4663 13512 4675 13515
rect 5258 13512 5264 13524
rect 4663 13484 5264 13512
rect 4663 13481 4675 13484
rect 4617 13475 4675 13481
rect 5258 13472 5264 13484
rect 5316 13472 5322 13524
rect 8202 13472 8208 13524
rect 8260 13512 8266 13524
rect 9309 13515 9367 13521
rect 9309 13512 9321 13515
rect 8260 13484 9321 13512
rect 8260 13472 8266 13484
rect 9309 13481 9321 13484
rect 9355 13481 9367 13515
rect 9309 13475 9367 13481
rect 11790 13472 11796 13524
rect 11848 13512 11854 13524
rect 12529 13515 12587 13521
rect 12529 13512 12541 13515
rect 11848 13484 12541 13512
rect 11848 13472 11854 13484
rect 12529 13481 12541 13484
rect 12575 13481 12587 13515
rect 12529 13475 12587 13481
rect 13541 13515 13599 13521
rect 13541 13481 13553 13515
rect 13587 13512 13599 13515
rect 14734 13512 14740 13524
rect 13587 13484 14740 13512
rect 13587 13481 13599 13484
rect 13541 13475 13599 13481
rect 14734 13472 14740 13484
rect 14792 13472 14798 13524
rect 17313 13515 17371 13521
rect 17313 13481 17325 13515
rect 17359 13512 17371 13515
rect 17494 13512 17500 13524
rect 17359 13484 17500 13512
rect 17359 13481 17371 13484
rect 17313 13475 17371 13481
rect 17494 13472 17500 13484
rect 17552 13512 17558 13524
rect 17552 13484 18644 13512
rect 17552 13472 17558 13484
rect 6457 13447 6515 13453
rect 6457 13413 6469 13447
rect 6503 13444 6515 13447
rect 13449 13447 13507 13453
rect 6503 13416 11836 13444
rect 6503 13413 6515 13416
rect 6457 13407 6515 13413
rect 3142 13336 3148 13388
rect 3200 13376 3206 13388
rect 5077 13379 5135 13385
rect 5077 13376 5089 13379
rect 3200 13348 5089 13376
rect 3200 13336 3206 13348
rect 5077 13345 5089 13348
rect 5123 13345 5135 13379
rect 5077 13339 5135 13345
rect 4249 13311 4307 13317
rect 4249 13277 4261 13311
rect 4295 13308 4307 13311
rect 4614 13308 4620 13320
rect 4295 13280 4620 13308
rect 4295 13277 4307 13280
rect 4249 13271 4307 13277
rect 4614 13268 4620 13280
rect 4672 13268 4678 13320
rect 5344 13311 5402 13317
rect 5344 13277 5356 13311
rect 5390 13308 5402 13311
rect 5718 13308 5724 13320
rect 5390 13280 5724 13308
rect 5390 13277 5402 13280
rect 5344 13271 5402 13277
rect 5718 13268 5724 13280
rect 5776 13268 5782 13320
rect 2222 13240 2228 13252
rect 2183 13212 2228 13240
rect 2222 13200 2228 13212
rect 2280 13200 2286 13252
rect 2314 13200 2320 13252
rect 2372 13240 2378 13252
rect 2409 13243 2467 13249
rect 2409 13240 2421 13243
rect 2372 13212 2421 13240
rect 2372 13200 2378 13212
rect 2409 13209 2421 13212
rect 2455 13209 2467 13243
rect 2409 13203 2467 13209
rect 4433 13243 4491 13249
rect 4433 13209 4445 13243
rect 4479 13240 4491 13243
rect 6472 13240 6500 13407
rect 7098 13376 7104 13388
rect 7059 13348 7104 13376
rect 7098 13336 7104 13348
rect 7156 13376 7162 13388
rect 7834 13376 7840 13388
rect 7156 13348 7840 13376
rect 7156 13336 7162 13348
rect 7834 13336 7840 13348
rect 7892 13336 7898 13388
rect 9674 13336 9680 13388
rect 9732 13376 9738 13388
rect 10229 13379 10287 13385
rect 10229 13376 10241 13379
rect 9732 13348 10241 13376
rect 9732 13336 9738 13348
rect 10229 13345 10241 13348
rect 10275 13345 10287 13379
rect 10229 13339 10287 13345
rect 6546 13268 6552 13320
rect 6604 13308 6610 13320
rect 7929 13311 7987 13317
rect 7929 13308 7941 13311
rect 6604 13280 7941 13308
rect 6604 13268 6610 13280
rect 7929 13277 7941 13280
rect 7975 13277 7987 13311
rect 9953 13311 10011 13317
rect 7929 13271 7987 13277
rect 8036 13280 9536 13308
rect 7285 13243 7343 13249
rect 7285 13240 7297 13243
rect 4479 13212 6500 13240
rect 6564 13212 7297 13240
rect 4479 13209 4491 13212
rect 4433 13203 4491 13209
rect 2041 13175 2099 13181
rect 2041 13141 2053 13175
rect 2087 13172 2099 13175
rect 2130 13172 2136 13184
rect 2087 13144 2136 13172
rect 2087 13141 2099 13144
rect 2041 13135 2099 13141
rect 2130 13132 2136 13144
rect 2188 13132 2194 13184
rect 5258 13132 5264 13184
rect 5316 13172 5322 13184
rect 6564 13172 6592 13212
rect 7285 13209 7297 13212
rect 7331 13240 7343 13243
rect 8036 13240 8064 13280
rect 7331 13212 8064 13240
rect 8113 13243 8171 13249
rect 7331 13209 7343 13212
rect 7285 13203 7343 13209
rect 8113 13209 8125 13243
rect 8159 13240 8171 13243
rect 8570 13240 8576 13252
rect 8159 13212 8576 13240
rect 8159 13209 8171 13212
rect 8113 13203 8171 13209
rect 8570 13200 8576 13212
rect 8628 13200 8634 13252
rect 8662 13200 8668 13252
rect 8720 13240 8726 13252
rect 9398 13240 9404 13252
rect 8720 13212 9404 13240
rect 8720 13200 8726 13212
rect 9398 13200 9404 13212
rect 9456 13200 9462 13252
rect 8294 13172 8300 13184
rect 5316 13144 6592 13172
rect 8255 13144 8300 13172
rect 5316 13132 5322 13144
rect 8294 13132 8300 13144
rect 8352 13132 8358 13184
rect 9508 13172 9536 13280
rect 9953 13277 9965 13311
rect 9999 13277 10011 13311
rect 9953 13271 10011 13277
rect 9968 13240 9996 13271
rect 11146 13268 11152 13320
rect 11204 13308 11210 13320
rect 11808 13317 11836 13416
rect 13449 13413 13461 13447
rect 13495 13444 13507 13447
rect 14461 13447 14519 13453
rect 14461 13444 14473 13447
rect 13495 13416 14473 13444
rect 13495 13413 13507 13416
rect 13449 13407 13507 13413
rect 14461 13413 14473 13416
rect 14507 13444 14519 13447
rect 15102 13444 15108 13456
rect 14507 13416 15108 13444
rect 14507 13413 14519 13416
rect 14461 13407 14519 13413
rect 15102 13404 15108 13416
rect 15160 13444 15166 13456
rect 16577 13447 16635 13453
rect 16577 13444 16589 13447
rect 15160 13416 16589 13444
rect 15160 13404 15166 13416
rect 16577 13413 16589 13416
rect 16623 13413 16635 13447
rect 16758 13444 16764 13456
rect 16719 13416 16764 13444
rect 16577 13407 16635 13413
rect 16758 13404 16764 13416
rect 16816 13404 16822 13456
rect 15286 13376 15292 13388
rect 15247 13348 15292 13376
rect 15286 13336 15292 13348
rect 15344 13336 15350 13388
rect 18616 13385 18644 13484
rect 19334 13472 19340 13524
rect 19392 13512 19398 13524
rect 19429 13515 19487 13521
rect 19429 13512 19441 13515
rect 19392 13484 19441 13512
rect 19392 13472 19398 13484
rect 19429 13481 19441 13484
rect 19475 13481 19487 13515
rect 19429 13475 19487 13481
rect 21269 13515 21327 13521
rect 21269 13481 21281 13515
rect 21315 13512 21327 13515
rect 26142 13512 26148 13524
rect 21315 13484 26148 13512
rect 21315 13481 21327 13484
rect 21269 13475 21327 13481
rect 26142 13472 26148 13484
rect 26200 13472 26206 13524
rect 35986 13512 35992 13524
rect 29840 13484 35848 13512
rect 35947 13484 35992 13512
rect 18601 13379 18659 13385
rect 18601 13345 18613 13379
rect 18647 13345 18659 13379
rect 18601 13339 18659 13345
rect 19334 13336 19340 13388
rect 19392 13376 19398 13388
rect 19886 13376 19892 13388
rect 19392 13348 19892 13376
rect 19392 13336 19398 13348
rect 19886 13336 19892 13348
rect 19944 13336 19950 13388
rect 23477 13379 23535 13385
rect 23477 13345 23489 13379
rect 23523 13376 23535 13379
rect 23842 13376 23848 13388
rect 23523 13348 23848 13376
rect 23523 13345 23535 13348
rect 23477 13339 23535 13345
rect 23842 13336 23848 13348
rect 23900 13376 23906 13388
rect 24302 13376 24308 13388
rect 23900 13348 24308 13376
rect 23900 13336 23906 13348
rect 24302 13336 24308 13348
rect 24360 13336 24366 13388
rect 24946 13336 24952 13388
rect 25004 13376 25010 13388
rect 25593 13379 25651 13385
rect 25593 13376 25605 13379
rect 25004 13348 25605 13376
rect 25004 13336 25010 13348
rect 25593 13345 25605 13348
rect 25639 13345 25651 13379
rect 25593 13339 25651 13345
rect 28644 13348 29132 13376
rect 11517 13311 11575 13317
rect 11517 13308 11529 13311
rect 11204 13280 11529 13308
rect 11204 13268 11210 13280
rect 11517 13277 11529 13280
rect 11563 13277 11575 13311
rect 11517 13271 11575 13277
rect 11793 13311 11851 13317
rect 11793 13277 11805 13311
rect 11839 13277 11851 13311
rect 11793 13271 11851 13277
rect 11882 13268 11888 13320
rect 11940 13308 11946 13320
rect 11940 13280 11985 13308
rect 11940 13268 11946 13280
rect 14550 13268 14556 13320
rect 14608 13268 14614 13320
rect 15194 13268 15200 13320
rect 15252 13308 15258 13320
rect 15381 13311 15439 13317
rect 15381 13308 15393 13311
rect 15252 13280 15393 13308
rect 15252 13268 15258 13280
rect 15381 13277 15393 13280
rect 15427 13277 15439 13311
rect 15381 13271 15439 13277
rect 15565 13311 15623 13317
rect 15565 13277 15577 13311
rect 15611 13277 15623 13311
rect 15565 13271 15623 13277
rect 18325 13311 18383 13317
rect 18325 13277 18337 13311
rect 18371 13277 18383 13311
rect 18325 13271 18383 13277
rect 19521 13311 19579 13317
rect 19521 13277 19533 13311
rect 19567 13277 19579 13311
rect 19521 13271 19579 13277
rect 19613 13311 19671 13317
rect 19613 13277 19625 13311
rect 19659 13308 19671 13311
rect 20070 13308 20076 13320
rect 19659 13280 20076 13308
rect 19659 13277 19671 13280
rect 19613 13271 19671 13277
rect 11698 13240 11704 13252
rect 9968 13212 11704 13240
rect 11698 13200 11704 13212
rect 11756 13200 11762 13252
rect 13081 13243 13139 13249
rect 11808 13212 12434 13240
rect 11808 13172 11836 13212
rect 12066 13172 12072 13184
rect 9508 13144 11836 13172
rect 12027 13144 12072 13172
rect 12066 13132 12072 13144
rect 12124 13132 12130 13184
rect 12406 13172 12434 13212
rect 13081 13209 13093 13243
rect 13127 13240 13139 13243
rect 13170 13240 13176 13252
rect 13127 13212 13176 13240
rect 13127 13209 13139 13212
rect 13081 13203 13139 13209
rect 13170 13200 13176 13212
rect 13228 13200 13234 13252
rect 13814 13240 13820 13252
rect 13464 13212 13820 13240
rect 13464 13172 13492 13212
rect 13814 13200 13820 13212
rect 13872 13200 13878 13252
rect 14093 13243 14151 13249
rect 14093 13209 14105 13243
rect 14139 13240 14151 13243
rect 14568 13240 14596 13268
rect 15580 13240 15608 13271
rect 16298 13240 16304 13252
rect 14139 13212 15608 13240
rect 16259 13212 16304 13240
rect 14139 13209 14151 13212
rect 14093 13203 14151 13209
rect 16298 13200 16304 13212
rect 16356 13200 16362 13252
rect 18340 13240 18368 13271
rect 18690 13240 18696 13252
rect 18340 13212 18696 13240
rect 18690 13200 18696 13212
rect 18748 13200 18754 13252
rect 19536 13240 19564 13271
rect 20070 13268 20076 13280
rect 20128 13268 20134 13320
rect 20714 13268 20720 13320
rect 20772 13308 20778 13320
rect 21085 13311 21143 13317
rect 21085 13308 21097 13311
rect 20772 13280 21097 13308
rect 20772 13268 20778 13280
rect 21085 13277 21097 13280
rect 21131 13277 21143 13311
rect 21085 13271 21143 13277
rect 23221 13311 23279 13317
rect 23221 13277 23233 13311
rect 23267 13308 23279 13311
rect 24762 13308 24768 13320
rect 23267 13280 24768 13308
rect 23267 13277 23279 13280
rect 23221 13271 23279 13277
rect 24762 13268 24768 13280
rect 24820 13268 24826 13320
rect 25314 13308 25320 13320
rect 25275 13280 25320 13308
rect 25314 13268 25320 13280
rect 25372 13268 25378 13320
rect 26234 13308 26240 13320
rect 26195 13280 26240 13308
rect 26234 13268 26240 13280
rect 26292 13268 26298 13320
rect 28644 13317 28672 13348
rect 29104 13320 29132 13348
rect 28629 13311 28687 13317
rect 28629 13277 28641 13311
rect 28675 13277 28687 13311
rect 28629 13271 28687 13277
rect 28718 13268 28724 13320
rect 28776 13308 28782 13320
rect 28994 13308 29000 13320
rect 28776 13280 28821 13308
rect 28955 13280 29000 13308
rect 28776 13268 28782 13280
rect 28994 13268 29000 13280
rect 29052 13268 29058 13320
rect 29086 13268 29092 13320
rect 29144 13308 29150 13320
rect 29840 13317 29868 13484
rect 30558 13444 30564 13456
rect 30519 13416 30564 13444
rect 30558 13404 30564 13416
rect 30616 13404 30622 13456
rect 34698 13404 34704 13456
rect 34756 13444 34762 13456
rect 34793 13447 34851 13453
rect 34793 13444 34805 13447
rect 34756 13416 34805 13444
rect 34756 13404 34762 13416
rect 34793 13413 34805 13416
rect 34839 13413 34851 13447
rect 35820 13444 35848 13484
rect 35986 13472 35992 13484
rect 36044 13472 36050 13524
rect 37369 13515 37427 13521
rect 37369 13481 37381 13515
rect 37415 13512 37427 13515
rect 37550 13512 37556 13524
rect 37415 13484 37556 13512
rect 37415 13481 37427 13484
rect 37369 13475 37427 13481
rect 37550 13472 37556 13484
rect 37608 13512 37614 13524
rect 38286 13512 38292 13524
rect 37608 13484 38292 13512
rect 37608 13472 37614 13484
rect 38286 13472 38292 13484
rect 38344 13472 38350 13524
rect 38746 13444 38752 13456
rect 35820 13416 38752 13444
rect 34793 13407 34851 13413
rect 32306 13336 32312 13388
rect 32364 13376 32370 13388
rect 32766 13376 32772 13388
rect 32364 13348 32772 13376
rect 32364 13336 32370 13348
rect 32766 13336 32772 13348
rect 32824 13336 32830 13388
rect 34149 13379 34207 13385
rect 34149 13345 34161 13379
rect 34195 13376 34207 13379
rect 34422 13376 34428 13388
rect 34195 13348 34428 13376
rect 34195 13345 34207 13348
rect 34149 13339 34207 13345
rect 29733 13311 29791 13317
rect 29733 13308 29745 13311
rect 29144 13280 29745 13308
rect 29144 13268 29150 13280
rect 29733 13277 29745 13280
rect 29779 13277 29791 13311
rect 29733 13271 29791 13277
rect 29825 13311 29883 13317
rect 29825 13277 29837 13311
rect 29871 13277 29883 13311
rect 29825 13271 29883 13277
rect 30101 13311 30159 13317
rect 30101 13277 30113 13311
rect 30147 13308 30159 13311
rect 31294 13308 31300 13320
rect 30147 13280 31300 13308
rect 30147 13277 30159 13280
rect 30101 13271 30159 13277
rect 31294 13268 31300 13280
rect 31352 13268 31358 13320
rect 31938 13308 31944 13320
rect 31851 13280 31944 13308
rect 31938 13268 31944 13280
rect 31996 13308 32002 13320
rect 34164 13308 34192 13339
rect 34422 13336 34428 13348
rect 34480 13336 34486 13388
rect 34808 13376 34836 13407
rect 38746 13404 38752 13416
rect 38804 13404 38810 13456
rect 34808 13348 35756 13376
rect 35342 13308 35348 13320
rect 31996 13280 34192 13308
rect 35303 13280 35348 13308
rect 31996 13268 32002 13280
rect 35342 13268 35348 13280
rect 35400 13268 35406 13320
rect 35526 13308 35532 13320
rect 35487 13280 35532 13308
rect 35526 13268 35532 13280
rect 35584 13268 35590 13320
rect 35728 13317 35756 13348
rect 36814 13336 36820 13388
rect 36872 13376 36878 13388
rect 36872 13348 38792 13376
rect 36872 13336 36878 13348
rect 38764 13320 38792 13348
rect 35621 13311 35679 13317
rect 35621 13277 35633 13311
rect 35667 13277 35679 13311
rect 35621 13271 35679 13277
rect 35713 13311 35771 13317
rect 35713 13277 35725 13311
rect 35759 13308 35771 13311
rect 36906 13308 36912 13320
rect 35759 13280 36912 13308
rect 35759 13277 35771 13280
rect 35713 13271 35771 13277
rect 19536 13212 24440 13240
rect 12406 13144 13492 13172
rect 14553 13175 14611 13181
rect 14553 13141 14565 13175
rect 14599 13172 14611 13175
rect 14826 13172 14832 13184
rect 14599 13144 14832 13172
rect 14599 13141 14611 13144
rect 14553 13135 14611 13141
rect 14826 13132 14832 13144
rect 14884 13132 14890 13184
rect 19150 13132 19156 13184
rect 19208 13172 19214 13184
rect 19245 13175 19303 13181
rect 19245 13172 19257 13175
rect 19208 13144 19257 13172
rect 19208 13132 19214 13144
rect 19245 13141 19257 13144
rect 19291 13141 19303 13175
rect 19245 13135 19303 13141
rect 20625 13175 20683 13181
rect 20625 13141 20637 13175
rect 20671 13172 20683 13175
rect 20714 13172 20720 13184
rect 20671 13144 20720 13172
rect 20671 13141 20683 13144
rect 20625 13135 20683 13141
rect 20714 13132 20720 13144
rect 20772 13132 20778 13184
rect 22097 13175 22155 13181
rect 22097 13141 22109 13175
rect 22143 13172 22155 13175
rect 22278 13172 22284 13184
rect 22143 13144 22284 13172
rect 22143 13141 22155 13144
rect 22097 13135 22155 13141
rect 22278 13132 22284 13144
rect 22336 13172 22342 13184
rect 22554 13172 22560 13184
rect 22336 13144 22560 13172
rect 22336 13132 22342 13144
rect 22554 13132 22560 13144
rect 22612 13132 22618 13184
rect 24412 13172 24440 13212
rect 26050 13200 26056 13252
rect 26108 13240 26114 13252
rect 26482 13243 26540 13249
rect 26482 13240 26494 13243
rect 26108 13212 26494 13240
rect 26108 13200 26114 13212
rect 26482 13209 26494 13212
rect 26528 13209 26540 13243
rect 26482 13203 26540 13209
rect 28813 13243 28871 13249
rect 28813 13209 28825 13243
rect 28859 13240 28871 13243
rect 29178 13240 29184 13252
rect 28859 13212 29184 13240
rect 28859 13209 28871 13212
rect 28813 13203 28871 13209
rect 29178 13200 29184 13212
rect 29236 13240 29242 13252
rect 29914 13240 29920 13252
rect 29236 13212 29920 13240
rect 29236 13200 29242 13212
rect 29914 13200 29920 13212
rect 29972 13200 29978 13252
rect 31696 13243 31754 13249
rect 31696 13209 31708 13243
rect 31742 13240 31754 13243
rect 32398 13240 32404 13252
rect 31742 13212 32404 13240
rect 31742 13209 31754 13212
rect 31696 13203 31754 13209
rect 32398 13200 32404 13212
rect 32456 13200 32462 13252
rect 33134 13200 33140 13252
rect 33192 13240 33198 13252
rect 33882 13243 33940 13249
rect 33882 13240 33894 13243
rect 33192 13212 33894 13240
rect 33192 13200 33198 13212
rect 33882 13209 33894 13212
rect 33928 13209 33940 13243
rect 35636 13240 35664 13271
rect 36906 13268 36912 13280
rect 36964 13268 36970 13320
rect 37550 13268 37556 13320
rect 37608 13308 37614 13320
rect 37829 13311 37887 13317
rect 37829 13308 37841 13311
rect 37608 13280 37841 13308
rect 37608 13268 37614 13280
rect 37829 13277 37841 13280
rect 37875 13277 37887 13311
rect 38010 13308 38016 13320
rect 37971 13280 38016 13308
rect 37829 13271 37887 13277
rect 38010 13268 38016 13280
rect 38068 13268 38074 13320
rect 38105 13311 38163 13317
rect 38105 13277 38117 13311
rect 38151 13277 38163 13311
rect 38105 13271 38163 13277
rect 38197 13311 38255 13317
rect 38197 13277 38209 13311
rect 38243 13308 38255 13311
rect 38286 13308 38292 13320
rect 38243 13280 38292 13308
rect 38243 13277 38255 13280
rect 38197 13271 38255 13277
rect 35986 13240 35992 13252
rect 35636 13212 35992 13240
rect 33882 13203 33940 13209
rect 35986 13200 35992 13212
rect 36044 13200 36050 13252
rect 38120 13184 38148 13271
rect 38286 13268 38292 13280
rect 38344 13268 38350 13320
rect 38746 13268 38752 13320
rect 38804 13308 38810 13320
rect 39301 13311 39359 13317
rect 39301 13308 39313 13311
rect 38804 13280 39313 13308
rect 38804 13268 38810 13280
rect 39301 13277 39313 13280
rect 39347 13308 39359 13311
rect 40221 13311 40279 13317
rect 40221 13308 40233 13311
rect 39347 13280 40233 13308
rect 39347 13277 39359 13280
rect 39301 13271 39359 13277
rect 40221 13277 40233 13280
rect 40267 13277 40279 13311
rect 68094 13308 68100 13320
rect 68055 13280 68100 13308
rect 40221 13271 40279 13277
rect 68094 13268 68100 13280
rect 68152 13268 68158 13320
rect 26786 13172 26792 13184
rect 24412 13144 26792 13172
rect 26786 13132 26792 13144
rect 26844 13132 26850 13184
rect 27246 13132 27252 13184
rect 27304 13172 27310 13184
rect 27617 13175 27675 13181
rect 27617 13172 27629 13175
rect 27304 13144 27629 13172
rect 27304 13132 27310 13144
rect 27617 13141 27629 13144
rect 27663 13141 27675 13175
rect 27617 13135 27675 13141
rect 28258 13132 28264 13184
rect 28316 13172 28322 13184
rect 28445 13175 28503 13181
rect 28445 13172 28457 13175
rect 28316 13144 28457 13172
rect 28316 13132 28322 13144
rect 28445 13141 28457 13144
rect 28491 13141 28503 13175
rect 29546 13172 29552 13184
rect 29507 13144 29552 13172
rect 28445 13135 28503 13141
rect 29546 13132 29552 13144
rect 29604 13132 29610 13184
rect 32766 13172 32772 13184
rect 32727 13144 32772 13172
rect 32766 13132 32772 13144
rect 32824 13132 32830 13184
rect 38102 13132 38108 13184
rect 38160 13132 38166 13184
rect 38470 13172 38476 13184
rect 38431 13144 38476 13172
rect 38470 13132 38476 13144
rect 38528 13132 38534 13184
rect 41230 13132 41236 13184
rect 41288 13172 41294 13184
rect 41509 13175 41567 13181
rect 41509 13172 41521 13175
rect 41288 13144 41521 13172
rect 41288 13132 41294 13144
rect 41509 13141 41521 13144
rect 41555 13141 41567 13175
rect 41509 13135 41567 13141
rect 1104 13082 68816 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 68816 13082
rect 1104 13008 68816 13030
rect 2222 12928 2228 12980
rect 2280 12968 2286 12980
rect 4525 12971 4583 12977
rect 4525 12968 4537 12971
rect 2280 12940 4537 12968
rect 2280 12928 2286 12940
rect 4525 12937 4537 12940
rect 4571 12937 4583 12971
rect 5258 12968 5264 12980
rect 5219 12940 5264 12968
rect 4525 12931 4583 12937
rect 3786 12900 3792 12912
rect 2700 12872 3792 12900
rect 2700 12841 2728 12872
rect 3786 12860 3792 12872
rect 3844 12860 3850 12912
rect 4540 12900 4568 12931
rect 5258 12928 5264 12940
rect 5316 12928 5322 12980
rect 5810 12928 5816 12980
rect 5868 12968 5874 12980
rect 6457 12971 6515 12977
rect 6457 12968 6469 12971
rect 5868 12940 6469 12968
rect 5868 12928 5874 12940
rect 6457 12937 6469 12940
rect 6503 12968 6515 12971
rect 6546 12968 6552 12980
rect 6503 12940 6552 12968
rect 6503 12937 6515 12940
rect 6457 12931 6515 12937
rect 6546 12928 6552 12940
rect 6604 12928 6610 12980
rect 8570 12928 8576 12980
rect 8628 12968 8634 12980
rect 9766 12968 9772 12980
rect 8628 12940 9772 12968
rect 8628 12928 8634 12940
rect 9766 12928 9772 12940
rect 9824 12928 9830 12980
rect 16298 12968 16304 12980
rect 12728 12940 16304 12968
rect 4540 12872 9444 12900
rect 2685 12835 2743 12841
rect 2685 12801 2697 12835
rect 2731 12801 2743 12835
rect 3142 12832 3148 12844
rect 3103 12804 3148 12832
rect 2685 12795 2743 12801
rect 3142 12792 3148 12804
rect 3200 12792 3206 12844
rect 3234 12792 3240 12844
rect 3292 12832 3298 12844
rect 3401 12835 3459 12841
rect 3401 12832 3413 12835
rect 3292 12804 3413 12832
rect 3292 12792 3298 12804
rect 3401 12801 3413 12804
rect 3447 12801 3459 12835
rect 6638 12832 6644 12844
rect 6599 12804 6644 12832
rect 3401 12795 3459 12801
rect 6638 12792 6644 12804
rect 6696 12792 6702 12844
rect 7929 12835 7987 12841
rect 7929 12801 7941 12835
rect 7975 12832 7987 12835
rect 8018 12832 8024 12844
rect 7975 12804 8024 12832
rect 7975 12801 7987 12804
rect 7929 12795 7987 12801
rect 8018 12792 8024 12804
rect 8076 12792 8082 12844
rect 8202 12792 8208 12844
rect 8260 12832 8266 12844
rect 8645 12835 8703 12841
rect 8645 12832 8657 12835
rect 8260 12804 8657 12832
rect 8260 12792 8266 12804
rect 8645 12801 8657 12804
rect 8691 12801 8703 12835
rect 8645 12795 8703 12801
rect 2222 12724 2228 12776
rect 2280 12764 2286 12776
rect 2409 12767 2467 12773
rect 2409 12764 2421 12767
rect 2280 12736 2421 12764
rect 2280 12724 2286 12736
rect 2409 12733 2421 12736
rect 2455 12733 2467 12767
rect 2409 12727 2467 12733
rect 5813 12767 5871 12773
rect 5813 12733 5825 12767
rect 5859 12764 5871 12767
rect 7466 12764 7472 12776
rect 5859 12736 7472 12764
rect 5859 12733 5871 12736
rect 5813 12727 5871 12733
rect 7466 12724 7472 12736
rect 7524 12724 7530 12776
rect 7653 12767 7711 12773
rect 7653 12733 7665 12767
rect 7699 12764 7711 12767
rect 7742 12764 7748 12776
rect 7699 12736 7748 12764
rect 7699 12733 7711 12736
rect 7653 12727 7711 12733
rect 7742 12724 7748 12736
rect 7800 12724 7806 12776
rect 8386 12764 8392 12776
rect 8347 12736 8392 12764
rect 8386 12724 8392 12736
rect 8444 12724 8450 12776
rect 9416 12764 9444 12872
rect 10502 12860 10508 12912
rect 10560 12900 10566 12912
rect 11698 12900 11704 12912
rect 10560 12872 10605 12900
rect 11659 12872 11704 12900
rect 10560 12860 10566 12872
rect 11698 12860 11704 12872
rect 11756 12860 11762 12912
rect 10134 12792 10140 12844
rect 10192 12832 10198 12844
rect 10229 12835 10287 12841
rect 10229 12832 10241 12835
rect 10192 12804 10241 12832
rect 10192 12792 10198 12804
rect 10229 12801 10241 12804
rect 10275 12801 10287 12835
rect 10410 12832 10416 12844
rect 10371 12804 10416 12832
rect 10229 12795 10287 12801
rect 10410 12792 10416 12804
rect 10468 12792 10474 12844
rect 10594 12832 10600 12844
rect 10555 12804 10600 12832
rect 10594 12792 10600 12804
rect 10652 12792 10658 12844
rect 11514 12832 11520 12844
rect 11475 12804 11520 12832
rect 11514 12792 11520 12804
rect 11572 12792 11578 12844
rect 11793 12835 11851 12841
rect 11793 12801 11805 12835
rect 11839 12801 11851 12835
rect 11793 12795 11851 12801
rect 11808 12764 11836 12795
rect 11882 12792 11888 12844
rect 11940 12832 11946 12844
rect 12728 12841 12756 12940
rect 16298 12928 16304 12940
rect 16356 12968 16362 12980
rect 17954 12968 17960 12980
rect 16356 12940 17960 12968
rect 16356 12928 16362 12940
rect 17954 12928 17960 12940
rect 18012 12928 18018 12980
rect 18049 12971 18107 12977
rect 18049 12937 18061 12971
rect 18095 12968 18107 12971
rect 18138 12968 18144 12980
rect 18095 12940 18144 12968
rect 18095 12937 18107 12940
rect 18049 12931 18107 12937
rect 18138 12928 18144 12940
rect 18196 12928 18202 12980
rect 19242 12968 19248 12980
rect 18248 12940 19248 12968
rect 15194 12900 15200 12912
rect 12912 12872 15200 12900
rect 12912 12841 12940 12872
rect 15194 12860 15200 12872
rect 15252 12860 15258 12912
rect 12713 12835 12771 12841
rect 11940 12804 11985 12832
rect 11940 12792 11946 12804
rect 12713 12801 12725 12835
rect 12759 12801 12771 12835
rect 12713 12795 12771 12801
rect 12897 12835 12955 12841
rect 12897 12801 12909 12835
rect 12943 12801 12955 12835
rect 12897 12795 12955 12801
rect 13725 12835 13783 12841
rect 13725 12801 13737 12835
rect 13771 12832 13783 12835
rect 13814 12832 13820 12844
rect 13771 12804 13820 12832
rect 13771 12801 13783 12804
rect 13725 12795 13783 12801
rect 13814 12792 13820 12804
rect 13872 12832 13878 12844
rect 14182 12832 14188 12844
rect 13872 12804 14188 12832
rect 13872 12792 13878 12804
rect 14182 12792 14188 12804
rect 14240 12792 14246 12844
rect 15289 12835 15347 12841
rect 15289 12801 15301 12835
rect 15335 12832 15347 12835
rect 15378 12832 15384 12844
rect 15335 12804 15384 12832
rect 15335 12801 15347 12804
rect 15289 12795 15347 12801
rect 15378 12792 15384 12804
rect 15436 12832 15442 12844
rect 15562 12832 15568 12844
rect 15436 12804 15568 12832
rect 15436 12792 15442 12804
rect 15562 12792 15568 12804
rect 15620 12792 15626 12844
rect 17589 12835 17647 12841
rect 17589 12801 17601 12835
rect 17635 12832 17647 12835
rect 18248 12832 18276 12940
rect 19242 12928 19248 12940
rect 19300 12928 19306 12980
rect 20073 12971 20131 12977
rect 20073 12937 20085 12971
rect 20119 12968 20131 12971
rect 20162 12968 20168 12980
rect 20119 12940 20168 12968
rect 20119 12937 20131 12940
rect 20073 12931 20131 12937
rect 20162 12928 20168 12940
rect 20220 12928 20226 12980
rect 22094 12928 22100 12980
rect 22152 12968 22158 12980
rect 22373 12971 22431 12977
rect 22373 12968 22385 12971
rect 22152 12940 22385 12968
rect 22152 12928 22158 12940
rect 22373 12937 22385 12940
rect 22419 12937 22431 12971
rect 22373 12931 22431 12937
rect 23382 12928 23388 12980
rect 23440 12968 23446 12980
rect 24121 12971 24179 12977
rect 24121 12968 24133 12971
rect 23440 12940 24133 12968
rect 23440 12928 23446 12940
rect 24121 12937 24133 12940
rect 24167 12937 24179 12971
rect 24121 12931 24179 12937
rect 24949 12971 25007 12977
rect 24949 12937 24961 12971
rect 24995 12968 25007 12971
rect 25222 12968 25228 12980
rect 24995 12940 25228 12968
rect 24995 12937 25007 12940
rect 24949 12931 25007 12937
rect 25222 12928 25228 12940
rect 25280 12928 25286 12980
rect 26050 12968 26056 12980
rect 26011 12940 26056 12968
rect 26050 12928 26056 12940
rect 26108 12928 26114 12980
rect 26973 12971 27031 12977
rect 26973 12937 26985 12971
rect 27019 12968 27031 12971
rect 27154 12968 27160 12980
rect 27019 12940 27160 12968
rect 27019 12937 27031 12940
rect 26973 12931 27031 12937
rect 27154 12928 27160 12940
rect 27212 12928 27218 12980
rect 27706 12928 27712 12980
rect 27764 12968 27770 12980
rect 28077 12971 28135 12977
rect 28077 12968 28089 12971
rect 27764 12940 28089 12968
rect 27764 12928 27770 12940
rect 28077 12937 28089 12940
rect 28123 12968 28135 12971
rect 28902 12968 28908 12980
rect 28123 12940 28908 12968
rect 28123 12937 28135 12940
rect 28077 12931 28135 12937
rect 28902 12928 28908 12940
rect 28960 12928 28966 12980
rect 38930 12928 38936 12980
rect 38988 12968 38994 12980
rect 39853 12971 39911 12977
rect 39853 12968 39865 12971
rect 38988 12940 39865 12968
rect 38988 12928 38994 12940
rect 39853 12937 39865 12940
rect 39899 12937 39911 12971
rect 39853 12931 39911 12937
rect 19518 12900 19524 12912
rect 18432 12872 19524 12900
rect 18432 12841 18460 12872
rect 19518 12860 19524 12872
rect 19576 12900 19582 12912
rect 19576 12872 19748 12900
rect 19576 12860 19582 12872
rect 17635 12804 18276 12832
rect 18325 12835 18383 12841
rect 17635 12801 17647 12804
rect 17589 12795 17647 12801
rect 18325 12801 18337 12835
rect 18371 12801 18383 12835
rect 18325 12795 18383 12801
rect 18417 12835 18475 12841
rect 18417 12801 18429 12835
rect 18463 12801 18475 12835
rect 18417 12795 18475 12801
rect 16850 12764 16856 12776
rect 9416 12736 11836 12764
rect 13556 12736 16856 12764
rect 9766 12696 9772 12708
rect 9679 12668 9772 12696
rect 9766 12656 9772 12668
rect 9824 12696 9830 12708
rect 11514 12696 11520 12708
rect 9824 12668 11520 12696
rect 9824 12656 9830 12668
rect 11514 12656 11520 12668
rect 11572 12656 11578 12708
rect 12066 12696 12072 12708
rect 12027 12668 12072 12696
rect 12066 12656 12072 12668
rect 12124 12656 12130 12708
rect 12802 12656 12808 12708
rect 12860 12696 12866 12708
rect 13556 12705 13584 12736
rect 16850 12724 16856 12736
rect 16908 12724 16914 12776
rect 17494 12764 17500 12776
rect 17455 12736 17500 12764
rect 17494 12724 17500 12736
rect 17552 12724 17558 12776
rect 18340 12764 18368 12795
rect 18506 12792 18512 12844
rect 18564 12832 18570 12844
rect 18564 12804 18609 12832
rect 18564 12792 18570 12804
rect 18690 12792 18696 12844
rect 18748 12832 18754 12844
rect 19426 12832 19432 12844
rect 18748 12804 19432 12832
rect 18748 12792 18754 12804
rect 19426 12792 19432 12804
rect 19484 12792 19490 12844
rect 19720 12841 19748 12872
rect 19886 12860 19892 12912
rect 19944 12900 19950 12912
rect 19944 12872 20024 12900
rect 19944 12860 19950 12872
rect 19613 12835 19671 12841
rect 19613 12832 19625 12835
rect 19536 12804 19625 12832
rect 19058 12764 19064 12776
rect 18340 12736 19064 12764
rect 19058 12724 19064 12736
rect 19116 12724 19122 12776
rect 19536 12764 19564 12804
rect 19613 12801 19625 12804
rect 19659 12801 19671 12835
rect 19613 12795 19671 12801
rect 19705 12835 19763 12841
rect 19705 12801 19717 12835
rect 19751 12801 19763 12835
rect 19705 12795 19763 12801
rect 19794 12792 19800 12844
rect 19852 12832 19858 12844
rect 19996 12832 20024 12872
rect 20254 12860 20260 12912
rect 20312 12900 20318 12912
rect 22002 12900 22008 12912
rect 20312 12872 21864 12900
rect 21963 12872 22008 12900
rect 20312 12860 20318 12872
rect 20533 12835 20591 12841
rect 20533 12832 20545 12835
rect 19852 12804 19897 12832
rect 19996 12804 20545 12832
rect 19852 12792 19858 12804
rect 20533 12801 20545 12804
rect 20579 12801 20591 12835
rect 20533 12795 20591 12801
rect 20717 12835 20775 12841
rect 20717 12801 20729 12835
rect 20763 12832 20775 12835
rect 21266 12832 21272 12844
rect 20763 12804 21272 12832
rect 20763 12801 20775 12804
rect 20717 12795 20775 12801
rect 21266 12792 21272 12804
rect 21324 12832 21330 12844
rect 21836 12841 21864 12872
rect 22002 12860 22008 12872
rect 22060 12860 22066 12912
rect 22554 12860 22560 12912
rect 22612 12900 22618 12912
rect 24765 12903 24823 12909
rect 24765 12900 24777 12903
rect 22612 12872 24777 12900
rect 22612 12860 22618 12872
rect 24765 12869 24777 12872
rect 24811 12869 24823 12903
rect 24765 12863 24823 12869
rect 25498 12860 25504 12912
rect 25556 12900 25562 12912
rect 27246 12900 27252 12912
rect 25556 12872 25728 12900
rect 25556 12860 25562 12872
rect 21821 12835 21879 12841
rect 21324 12804 21772 12832
rect 21324 12792 21330 12804
rect 20901 12767 20959 12773
rect 20901 12764 20913 12767
rect 19536 12736 20913 12764
rect 20901 12733 20913 12736
rect 20947 12733 20959 12767
rect 20901 12727 20959 12733
rect 12897 12699 12955 12705
rect 12897 12696 12909 12699
rect 12860 12668 12909 12696
rect 12860 12656 12866 12668
rect 12897 12665 12909 12668
rect 12943 12665 12955 12699
rect 12897 12659 12955 12665
rect 13541 12699 13599 12705
rect 13541 12665 13553 12699
rect 13587 12665 13599 12699
rect 13541 12659 13599 12665
rect 14642 12656 14648 12708
rect 14700 12696 14706 12708
rect 15102 12696 15108 12708
rect 14700 12668 15108 12696
rect 14700 12656 14706 12668
rect 15102 12656 15108 12668
rect 15160 12696 15166 12708
rect 15565 12699 15623 12705
rect 15565 12696 15577 12699
rect 15160 12668 15577 12696
rect 15160 12656 15166 12668
rect 15565 12665 15577 12668
rect 15611 12665 15623 12699
rect 15746 12696 15752 12708
rect 15707 12668 15752 12696
rect 15565 12659 15623 12665
rect 15746 12656 15752 12668
rect 15804 12656 15810 12708
rect 21744 12696 21772 12804
rect 21821 12801 21833 12835
rect 21867 12801 21879 12835
rect 21821 12795 21879 12801
rect 22094 12792 22100 12844
rect 22152 12832 22158 12844
rect 22235 12835 22293 12841
rect 22152 12804 22197 12832
rect 22152 12792 22158 12804
rect 22235 12801 22247 12835
rect 22281 12832 22293 12835
rect 22370 12832 22376 12844
rect 22281 12804 22376 12832
rect 22281 12801 22293 12804
rect 22235 12795 22293 12801
rect 22370 12792 22376 12804
rect 22428 12792 22434 12844
rect 23474 12792 23480 12844
rect 23532 12832 23538 12844
rect 23661 12835 23719 12841
rect 23661 12832 23673 12835
rect 23532 12804 23673 12832
rect 23532 12792 23538 12804
rect 23661 12801 23673 12804
rect 23707 12801 23719 12835
rect 23934 12832 23940 12844
rect 23895 12804 23940 12832
rect 23661 12795 23719 12801
rect 23934 12792 23940 12804
rect 23992 12792 23998 12844
rect 24302 12792 24308 12844
rect 24360 12832 24366 12844
rect 24581 12835 24639 12841
rect 24581 12832 24593 12835
rect 24360 12804 24593 12832
rect 24360 12792 24366 12804
rect 24581 12801 24593 12804
rect 24627 12801 24639 12835
rect 24581 12795 24639 12801
rect 25314 12792 25320 12844
rect 25372 12832 25378 12844
rect 25409 12835 25467 12841
rect 25409 12832 25421 12835
rect 25372 12804 25421 12832
rect 25372 12792 25378 12804
rect 25409 12801 25421 12804
rect 25455 12801 25467 12835
rect 25590 12832 25596 12844
rect 25551 12804 25596 12832
rect 25409 12795 25467 12801
rect 25590 12792 25596 12804
rect 25648 12792 25654 12844
rect 25700 12841 25728 12872
rect 26988 12872 27252 12900
rect 26988 12844 27016 12872
rect 27246 12860 27252 12872
rect 27304 12860 27310 12912
rect 27341 12903 27399 12909
rect 27341 12869 27353 12903
rect 27387 12900 27399 12903
rect 27798 12900 27804 12912
rect 27387 12872 27804 12900
rect 27387 12869 27399 12872
rect 27341 12863 27399 12869
rect 27798 12860 27804 12872
rect 27856 12860 27862 12912
rect 29454 12860 29460 12912
rect 29512 12900 29518 12912
rect 32401 12903 32459 12909
rect 32401 12900 32413 12903
rect 29512 12872 32413 12900
rect 29512 12860 29518 12872
rect 32401 12869 32413 12872
rect 32447 12900 32459 12903
rect 32766 12900 32772 12912
rect 32447 12872 32772 12900
rect 32447 12869 32459 12872
rect 32401 12863 32459 12869
rect 32766 12860 32772 12872
rect 32824 12860 32830 12912
rect 35434 12860 35440 12912
rect 35492 12900 35498 12912
rect 35710 12900 35716 12912
rect 35492 12872 35716 12900
rect 35492 12860 35498 12872
rect 35710 12860 35716 12872
rect 35768 12860 35774 12912
rect 38470 12860 38476 12912
rect 38528 12900 38534 12912
rect 40966 12903 41024 12909
rect 40966 12900 40978 12903
rect 38528 12872 40978 12900
rect 38528 12860 38534 12872
rect 40966 12869 40978 12872
rect 41012 12869 41024 12903
rect 40966 12863 41024 12869
rect 25685 12835 25743 12841
rect 25685 12801 25697 12835
rect 25731 12801 25743 12835
rect 25685 12795 25743 12801
rect 25777 12835 25835 12841
rect 25777 12801 25789 12835
rect 25823 12832 25835 12835
rect 26878 12832 26884 12844
rect 25823 12804 26884 12832
rect 25823 12801 25835 12804
rect 25777 12795 25835 12801
rect 26878 12792 26884 12804
rect 26936 12792 26942 12844
rect 26970 12792 26976 12844
rect 27028 12792 27034 12844
rect 27157 12835 27215 12841
rect 27157 12801 27169 12835
rect 27203 12801 27215 12835
rect 27157 12795 27215 12801
rect 27525 12835 27583 12841
rect 27525 12801 27537 12835
rect 27571 12801 27583 12835
rect 27525 12795 27583 12801
rect 23750 12764 23756 12776
rect 23711 12736 23756 12764
rect 23750 12724 23756 12736
rect 23808 12724 23814 12776
rect 23860 12736 24072 12764
rect 23860 12696 23888 12736
rect 21744 12668 23888 12696
rect 24044 12696 24072 12736
rect 26326 12724 26332 12776
rect 26384 12764 26390 12776
rect 27172 12764 27200 12795
rect 26384 12736 27200 12764
rect 26384 12724 26390 12736
rect 27540 12696 27568 12795
rect 27982 12792 27988 12844
rect 28040 12832 28046 12844
rect 28813 12835 28871 12841
rect 28813 12832 28825 12835
rect 28040 12804 28825 12832
rect 28040 12792 28046 12804
rect 28813 12801 28825 12804
rect 28859 12801 28871 12835
rect 29086 12832 29092 12844
rect 29047 12804 29092 12832
rect 28813 12795 28871 12801
rect 29086 12792 29092 12804
rect 29144 12792 29150 12844
rect 31846 12792 31852 12844
rect 31904 12832 31910 12844
rect 32122 12832 32128 12844
rect 31904 12804 32128 12832
rect 31904 12792 31910 12804
rect 32122 12792 32128 12804
rect 32180 12832 32186 12844
rect 32217 12835 32275 12841
rect 32217 12832 32229 12835
rect 32180 12804 32229 12832
rect 32180 12792 32186 12804
rect 32217 12801 32229 12804
rect 32263 12801 32275 12835
rect 35894 12832 35900 12844
rect 35807 12804 35900 12832
rect 32217 12795 32275 12801
rect 35894 12792 35900 12804
rect 35952 12832 35958 12844
rect 37550 12832 37556 12844
rect 35952 12804 37412 12832
rect 37511 12804 37556 12832
rect 35952 12792 35958 12804
rect 35250 12724 35256 12776
rect 35308 12764 35314 12776
rect 35434 12764 35440 12776
rect 35308 12736 35440 12764
rect 35308 12724 35314 12736
rect 35434 12724 35440 12736
rect 35492 12724 35498 12776
rect 37274 12764 37280 12776
rect 37235 12736 37280 12764
rect 37274 12724 37280 12736
rect 37332 12724 37338 12776
rect 37384 12764 37412 12804
rect 37550 12792 37556 12804
rect 37608 12792 37614 12844
rect 38654 12792 38660 12844
rect 38712 12832 38718 12844
rect 38749 12835 38807 12841
rect 38749 12832 38761 12835
rect 38712 12804 38761 12832
rect 38712 12792 38718 12804
rect 38749 12801 38761 12804
rect 38795 12801 38807 12835
rect 38749 12795 38807 12801
rect 38838 12792 38844 12844
rect 38896 12832 38902 12844
rect 38933 12835 38991 12841
rect 38933 12832 38945 12835
rect 38896 12804 38945 12832
rect 38896 12792 38902 12804
rect 38933 12801 38945 12804
rect 38979 12801 38991 12835
rect 41230 12832 41236 12844
rect 41191 12804 41236 12832
rect 38933 12795 38991 12801
rect 41230 12792 41236 12804
rect 41288 12792 41294 12844
rect 38856 12764 38884 12792
rect 37384 12736 38884 12764
rect 36538 12696 36544 12708
rect 24044 12668 27568 12696
rect 34900 12668 36544 12696
rect 10778 12628 10784 12640
rect 10739 12600 10784 12628
rect 10778 12588 10784 12600
rect 10836 12588 10842 12640
rect 11054 12588 11060 12640
rect 11112 12628 11118 12640
rect 11882 12628 11888 12640
rect 11112 12600 11888 12628
rect 11112 12588 11118 12600
rect 11882 12588 11888 12600
rect 11940 12588 11946 12640
rect 14182 12628 14188 12640
rect 14143 12600 14188 12628
rect 14182 12588 14188 12600
rect 14240 12588 14246 12640
rect 17218 12628 17224 12640
rect 17179 12600 17224 12628
rect 17218 12588 17224 12600
rect 17276 12588 17282 12640
rect 17589 12631 17647 12637
rect 17589 12597 17601 12631
rect 17635 12628 17647 12631
rect 17862 12628 17868 12640
rect 17635 12600 17868 12628
rect 17635 12597 17647 12600
rect 17589 12591 17647 12597
rect 17862 12588 17868 12600
rect 17920 12588 17926 12640
rect 23937 12631 23995 12637
rect 23937 12597 23949 12631
rect 23983 12628 23995 12631
rect 25774 12628 25780 12640
rect 23983 12600 25780 12628
rect 23983 12597 23995 12600
rect 23937 12591 23995 12597
rect 25774 12588 25780 12600
rect 25832 12588 25838 12640
rect 27614 12588 27620 12640
rect 27672 12628 27678 12640
rect 30650 12628 30656 12640
rect 27672 12600 30656 12628
rect 27672 12588 27678 12600
rect 30650 12588 30656 12600
rect 30708 12588 30714 12640
rect 32585 12631 32643 12637
rect 32585 12597 32597 12631
rect 32631 12628 32643 12631
rect 32674 12628 32680 12640
rect 32631 12600 32680 12628
rect 32631 12597 32643 12600
rect 32585 12591 32643 12597
rect 32674 12588 32680 12600
rect 32732 12588 32738 12640
rect 34790 12588 34796 12640
rect 34848 12628 34854 12640
rect 34900 12637 34928 12668
rect 36538 12656 36544 12668
rect 36596 12656 36602 12708
rect 34885 12631 34943 12637
rect 34885 12628 34897 12631
rect 34848 12600 34897 12628
rect 34848 12588 34854 12600
rect 34885 12597 34897 12600
rect 34931 12597 34943 12631
rect 35526 12628 35532 12640
rect 35487 12600 35532 12628
rect 34885 12591 34943 12597
rect 35526 12588 35532 12600
rect 35584 12588 35590 12640
rect 37826 12588 37832 12640
rect 37884 12628 37890 12640
rect 38565 12631 38623 12637
rect 38565 12628 38577 12631
rect 37884 12600 38577 12628
rect 37884 12588 37890 12600
rect 38565 12597 38577 12600
rect 38611 12597 38623 12631
rect 38565 12591 38623 12597
rect 1104 12538 68816 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 65654 12538
rect 65706 12486 65718 12538
rect 65770 12486 65782 12538
rect 65834 12486 65846 12538
rect 65898 12486 65910 12538
rect 65962 12486 68816 12538
rect 1104 12464 68816 12486
rect 2593 12427 2651 12433
rect 2593 12393 2605 12427
rect 2639 12424 2651 12427
rect 3234 12424 3240 12436
rect 2639 12396 3240 12424
rect 2639 12393 2651 12396
rect 2593 12387 2651 12393
rect 3234 12384 3240 12396
rect 3292 12384 3298 12436
rect 5721 12427 5779 12433
rect 5721 12393 5733 12427
rect 5767 12424 5779 12427
rect 5902 12424 5908 12436
rect 5767 12396 5908 12424
rect 5767 12393 5779 12396
rect 5721 12387 5779 12393
rect 5902 12384 5908 12396
rect 5960 12384 5966 12436
rect 8202 12424 8208 12436
rect 8163 12396 8208 12424
rect 8202 12384 8208 12396
rect 8260 12384 8266 12436
rect 11698 12384 11704 12436
rect 11756 12424 11762 12436
rect 13081 12427 13139 12433
rect 13081 12424 13093 12427
rect 11756 12396 13093 12424
rect 11756 12384 11762 12396
rect 13081 12393 13093 12396
rect 13127 12393 13139 12427
rect 16206 12424 16212 12436
rect 13081 12387 13139 12393
rect 15120 12396 16212 12424
rect 2314 12316 2320 12368
rect 2372 12356 2378 12368
rect 3789 12359 3847 12365
rect 3789 12356 3801 12359
rect 2372 12328 3801 12356
rect 2372 12316 2378 12328
rect 3789 12325 3801 12328
rect 3835 12325 3847 12359
rect 7742 12356 7748 12368
rect 3789 12319 3847 12325
rect 6564 12328 7748 12356
rect 2038 12288 2044 12300
rect 1964 12260 2044 12288
rect 1964 12229 1992 12260
rect 2038 12248 2044 12260
rect 2096 12248 2102 12300
rect 1949 12223 2007 12229
rect 1949 12189 1961 12223
rect 1995 12189 2007 12223
rect 2130 12220 2136 12232
rect 2091 12192 2136 12220
rect 1949 12183 2007 12189
rect 2130 12180 2136 12192
rect 2188 12180 2194 12232
rect 2222 12180 2228 12232
rect 2280 12220 2286 12232
rect 2363 12223 2421 12229
rect 2280 12192 2325 12220
rect 2280 12180 2286 12192
rect 2363 12189 2375 12223
rect 2409 12220 2421 12223
rect 2498 12220 2504 12232
rect 2409 12192 2504 12220
rect 2409 12189 2421 12192
rect 2363 12183 2421 12189
rect 2498 12180 2504 12192
rect 2556 12220 2562 12232
rect 3053 12223 3111 12229
rect 3053 12220 3065 12223
rect 2556 12192 3065 12220
rect 2556 12180 2562 12192
rect 3053 12189 3065 12192
rect 3099 12189 3111 12223
rect 3053 12183 3111 12189
rect 3973 12223 4031 12229
rect 3973 12189 3985 12223
rect 4019 12220 4031 12223
rect 4614 12220 4620 12232
rect 4019 12192 4620 12220
rect 4019 12189 4031 12192
rect 3973 12183 4031 12189
rect 4614 12180 4620 12192
rect 4672 12180 4678 12232
rect 6362 12220 6368 12232
rect 5000 12192 6368 12220
rect 2774 12112 2780 12164
rect 2832 12152 2838 12164
rect 5000 12152 5028 12192
rect 6362 12180 6368 12192
rect 6420 12220 6426 12232
rect 6564 12229 6592 12328
rect 6457 12223 6515 12229
rect 6457 12220 6469 12223
rect 6420 12192 6469 12220
rect 6420 12180 6426 12192
rect 6457 12189 6469 12192
rect 6503 12189 6515 12223
rect 6457 12183 6515 12189
rect 6549 12223 6607 12229
rect 6549 12189 6561 12223
rect 6595 12189 6607 12223
rect 6549 12183 6607 12189
rect 6638 12180 6644 12232
rect 6696 12220 6702 12232
rect 6825 12223 6883 12229
rect 6696 12192 6741 12220
rect 6696 12180 6702 12192
rect 6825 12189 6837 12223
rect 6871 12220 6883 12223
rect 7190 12220 7196 12232
rect 6871 12192 7196 12220
rect 6871 12189 6883 12192
rect 6825 12183 6883 12189
rect 2832 12124 5028 12152
rect 5169 12155 5227 12161
rect 2832 12112 2838 12124
rect 5169 12121 5181 12155
rect 5215 12152 5227 12155
rect 6840 12152 6868 12183
rect 7190 12180 7196 12192
rect 7248 12220 7254 12232
rect 7561 12223 7619 12229
rect 7561 12220 7573 12223
rect 7248 12192 7573 12220
rect 7248 12180 7254 12192
rect 7561 12189 7573 12192
rect 7607 12189 7619 12223
rect 7561 12183 7619 12189
rect 5215 12124 6868 12152
rect 7668 12152 7696 12328
rect 7742 12316 7748 12328
rect 7800 12316 7806 12368
rect 9858 12316 9864 12368
rect 9916 12316 9922 12368
rect 14274 12316 14280 12368
rect 14332 12356 14338 12368
rect 14369 12359 14427 12365
rect 14369 12356 14381 12359
rect 14332 12328 14381 12356
rect 14332 12316 14338 12328
rect 14369 12325 14381 12328
rect 14415 12325 14427 12359
rect 14369 12319 14427 12325
rect 8294 12288 8300 12300
rect 7760 12260 8300 12288
rect 7760 12229 7788 12260
rect 8294 12248 8300 12260
rect 8352 12248 8358 12300
rect 9876 12288 9904 12316
rect 9508 12260 9904 12288
rect 10505 12291 10563 12297
rect 7724 12223 7788 12229
rect 7724 12189 7736 12223
rect 7770 12192 7788 12223
rect 7840 12220 7898 12226
rect 7840 12196 7852 12220
rect 7770 12189 7782 12192
rect 7724 12183 7782 12189
rect 7839 12186 7852 12196
rect 7886 12186 7898 12220
rect 7839 12180 7898 12186
rect 7926 12180 7932 12232
rect 7984 12220 7990 12232
rect 9508 12229 9536 12260
rect 10505 12257 10517 12291
rect 10551 12288 10563 12291
rect 11054 12288 11060 12300
rect 10551 12260 11060 12288
rect 10551 12257 10563 12260
rect 10505 12251 10563 12257
rect 11054 12248 11060 12260
rect 11112 12248 11118 12300
rect 13096 12260 14688 12288
rect 13096 12232 13124 12260
rect 9493 12223 9551 12229
rect 7984 12192 8029 12220
rect 7984 12180 7990 12192
rect 9493 12189 9505 12223
rect 9539 12189 9551 12223
rect 9769 12223 9827 12229
rect 9769 12220 9781 12223
rect 9493 12183 9551 12189
rect 9600 12192 9781 12220
rect 7839 12168 7880 12180
rect 7839 12152 7867 12168
rect 9600 12152 9628 12192
rect 9769 12189 9781 12192
rect 9815 12189 9827 12223
rect 9769 12183 9827 12189
rect 9861 12223 9919 12229
rect 9861 12189 9873 12223
rect 9907 12220 9919 12223
rect 10594 12220 10600 12232
rect 9907 12192 10600 12220
rect 9907 12189 9919 12192
rect 9861 12183 9919 12189
rect 10594 12180 10600 12192
rect 10652 12220 10658 12232
rect 12618 12229 12624 12232
rect 10781 12223 10839 12229
rect 10781 12220 10793 12223
rect 10652 12192 10793 12220
rect 10652 12180 10658 12192
rect 10781 12189 10793 12192
rect 10827 12189 10839 12223
rect 10781 12183 10839 12189
rect 11885 12223 11943 12229
rect 11885 12189 11897 12223
rect 11931 12220 11943 12223
rect 12614 12220 12624 12229
rect 11931 12192 12624 12220
rect 11931 12189 11943 12192
rect 11885 12183 11943 12189
rect 12614 12183 12624 12192
rect 12618 12180 12624 12183
rect 12676 12180 12682 12232
rect 13078 12220 13084 12232
rect 13039 12192 13084 12220
rect 13078 12180 13084 12192
rect 13136 12180 13142 12232
rect 13265 12223 13323 12229
rect 13265 12189 13277 12223
rect 13311 12220 13323 12223
rect 14093 12223 14151 12229
rect 14093 12220 14105 12223
rect 13311 12192 14105 12220
rect 13311 12189 13323 12192
rect 13265 12183 13323 12189
rect 14093 12189 14105 12192
rect 14139 12189 14151 12223
rect 14366 12220 14372 12232
rect 14327 12192 14372 12220
rect 14093 12183 14151 12189
rect 7668 12124 7867 12152
rect 8128 12124 9628 12152
rect 9677 12155 9735 12161
rect 5215 12121 5227 12124
rect 5169 12115 5227 12121
rect 4617 12087 4675 12093
rect 4617 12053 4629 12087
rect 4663 12084 4675 12087
rect 5184 12084 5212 12115
rect 6178 12084 6184 12096
rect 4663 12056 5212 12084
rect 6139 12056 6184 12084
rect 4663 12053 4675 12056
rect 4617 12047 4675 12053
rect 6178 12044 6184 12056
rect 6236 12044 6242 12096
rect 6454 12044 6460 12096
rect 6512 12084 6518 12096
rect 8128 12084 8156 12124
rect 9677 12121 9689 12155
rect 9723 12121 9735 12155
rect 10410 12152 10416 12164
rect 9677 12115 9735 12121
rect 9876 12124 10416 12152
rect 9030 12084 9036 12096
rect 6512 12056 8156 12084
rect 8991 12056 9036 12084
rect 6512 12044 6518 12056
rect 9030 12044 9036 12056
rect 9088 12044 9094 12096
rect 9692 12084 9720 12115
rect 9876 12084 9904 12124
rect 10410 12112 10416 12124
rect 10468 12112 10474 12164
rect 12894 12112 12900 12164
rect 12952 12152 12958 12164
rect 13280 12152 13308 12183
rect 14366 12180 14372 12192
rect 14424 12220 14430 12232
rect 14550 12220 14556 12232
rect 14424 12192 14556 12220
rect 14424 12180 14430 12192
rect 14550 12180 14556 12192
rect 14608 12180 14614 12232
rect 12952 12124 13308 12152
rect 14660 12152 14688 12260
rect 15120 12220 15148 12396
rect 16206 12384 16212 12396
rect 16264 12384 16270 12436
rect 17773 12427 17831 12433
rect 17773 12393 17785 12427
rect 17819 12424 17831 12427
rect 18506 12424 18512 12436
rect 17819 12396 18512 12424
rect 17819 12393 17831 12396
rect 17773 12387 17831 12393
rect 18506 12384 18512 12396
rect 18564 12384 18570 12436
rect 19794 12384 19800 12436
rect 19852 12424 19858 12436
rect 20254 12424 20260 12436
rect 19852 12396 20260 12424
rect 19852 12384 19858 12396
rect 20254 12384 20260 12396
rect 20312 12384 20318 12436
rect 22186 12384 22192 12436
rect 22244 12424 22250 12436
rect 22281 12427 22339 12433
rect 22281 12424 22293 12427
rect 22244 12396 22293 12424
rect 22244 12384 22250 12396
rect 22281 12393 22293 12396
rect 22327 12393 22339 12427
rect 24397 12427 24455 12433
rect 24397 12424 24409 12427
rect 22281 12387 22339 12393
rect 23860 12396 24409 12424
rect 15197 12359 15255 12365
rect 15197 12325 15209 12359
rect 15243 12356 15255 12359
rect 15286 12356 15292 12368
rect 15243 12328 15292 12356
rect 15243 12325 15255 12328
rect 15197 12319 15255 12325
rect 15286 12316 15292 12328
rect 15344 12316 15350 12368
rect 15470 12316 15476 12368
rect 15528 12356 15534 12368
rect 23860 12356 23888 12396
rect 24397 12393 24409 12396
rect 24443 12424 24455 12427
rect 24946 12424 24952 12436
rect 24443 12396 24952 12424
rect 24443 12393 24455 12396
rect 24397 12387 24455 12393
rect 24946 12384 24952 12396
rect 25004 12384 25010 12436
rect 25317 12427 25375 12433
rect 25317 12393 25329 12427
rect 25363 12424 25375 12427
rect 25590 12424 25596 12436
rect 25363 12396 25596 12424
rect 25363 12393 25375 12396
rect 25317 12387 25375 12393
rect 25590 12384 25596 12396
rect 25648 12384 25654 12436
rect 25866 12384 25872 12436
rect 25924 12424 25930 12436
rect 28258 12424 28264 12436
rect 25924 12396 27752 12424
rect 28219 12396 28264 12424
rect 25924 12384 25930 12396
rect 15528 12328 23888 12356
rect 15528 12316 15534 12328
rect 23934 12316 23940 12368
rect 23992 12356 23998 12368
rect 27614 12356 27620 12368
rect 23992 12328 27620 12356
rect 23992 12316 23998 12328
rect 27614 12316 27620 12328
rect 27672 12316 27678 12368
rect 27724 12356 27752 12396
rect 28258 12384 28264 12396
rect 28316 12384 28322 12436
rect 33134 12424 33140 12436
rect 31726 12396 32996 12424
rect 33095 12396 33140 12424
rect 31726 12356 31754 12396
rect 32674 12356 32680 12368
rect 27724 12328 31754 12356
rect 32600 12328 32680 12356
rect 16301 12291 16359 12297
rect 16301 12257 16313 12291
rect 16347 12288 16359 12291
rect 27890 12288 27896 12300
rect 16347 12260 27896 12288
rect 16347 12257 16359 12260
rect 16301 12251 16359 12257
rect 27890 12248 27896 12260
rect 27948 12248 27954 12300
rect 28074 12288 28080 12300
rect 28035 12260 28080 12288
rect 28074 12248 28080 12260
rect 28132 12248 28138 12300
rect 28166 12248 28172 12300
rect 28224 12288 28230 12300
rect 31941 12291 31999 12297
rect 31941 12288 31953 12291
rect 28224 12260 31953 12288
rect 28224 12248 28230 12260
rect 31941 12257 31953 12260
rect 31987 12257 31999 12291
rect 31941 12251 31999 12257
rect 15197 12223 15255 12229
rect 15197 12220 15209 12223
rect 15120 12192 15209 12220
rect 15197 12189 15209 12192
rect 15243 12189 15255 12223
rect 15197 12183 15255 12189
rect 15473 12223 15531 12229
rect 15473 12189 15485 12223
rect 15519 12189 15531 12223
rect 15473 12183 15531 12189
rect 15933 12223 15991 12229
rect 15933 12189 15945 12223
rect 15979 12189 15991 12223
rect 16206 12220 16212 12232
rect 16119 12192 16212 12220
rect 15933 12183 15991 12189
rect 15378 12152 15384 12164
rect 14660 12124 15384 12152
rect 12952 12112 12958 12124
rect 15378 12112 15384 12124
rect 15436 12152 15442 12164
rect 15497 12152 15525 12183
rect 15436 12124 15525 12152
rect 15436 12112 15442 12124
rect 10042 12084 10048 12096
rect 9692 12056 9904 12084
rect 10003 12056 10048 12084
rect 10042 12044 10048 12056
rect 10100 12044 10106 12096
rect 10962 12044 10968 12096
rect 11020 12084 11026 12096
rect 12437 12087 12495 12093
rect 12437 12084 12449 12087
rect 11020 12056 12449 12084
rect 11020 12044 11026 12056
rect 12437 12053 12449 12056
rect 12483 12053 12495 12087
rect 12437 12047 12495 12053
rect 13170 12044 13176 12096
rect 13228 12084 13234 12096
rect 15948 12084 15976 12183
rect 16206 12180 16212 12192
rect 16264 12220 16270 12232
rect 17862 12220 17868 12232
rect 16264 12192 17868 12220
rect 16264 12180 16270 12192
rect 17862 12180 17868 12192
rect 17920 12180 17926 12232
rect 17957 12223 18015 12229
rect 17957 12189 17969 12223
rect 18003 12220 18015 12223
rect 19334 12220 19340 12232
rect 18003 12192 19340 12220
rect 18003 12189 18015 12192
rect 17957 12183 18015 12189
rect 19334 12180 19340 12192
rect 19392 12180 19398 12232
rect 19705 12223 19763 12229
rect 19705 12189 19717 12223
rect 19751 12220 19763 12223
rect 19794 12220 19800 12232
rect 19751 12192 19800 12220
rect 19751 12189 19763 12192
rect 19705 12183 19763 12189
rect 18138 12152 18144 12164
rect 18051 12124 18144 12152
rect 18138 12112 18144 12124
rect 18196 12152 18202 12164
rect 19720 12152 19748 12183
rect 19794 12180 19800 12192
rect 19852 12180 19858 12232
rect 20254 12180 20260 12232
rect 20312 12220 20318 12232
rect 21729 12223 21787 12229
rect 21729 12220 21741 12223
rect 20312 12192 21741 12220
rect 20312 12180 20318 12192
rect 21729 12189 21741 12192
rect 21775 12189 21787 12223
rect 21729 12183 21787 12189
rect 22097 12223 22155 12229
rect 22097 12189 22109 12223
rect 22143 12220 22155 12223
rect 22370 12220 22376 12232
rect 22143 12192 22376 12220
rect 22143 12189 22155 12192
rect 22097 12183 22155 12189
rect 22370 12180 22376 12192
rect 22428 12220 22434 12232
rect 23014 12220 23020 12232
rect 22428 12192 23020 12220
rect 22428 12180 22434 12192
rect 23014 12180 23020 12192
rect 23072 12180 23078 12232
rect 25133 12223 25191 12229
rect 25133 12189 25145 12223
rect 25179 12220 25191 12223
rect 26970 12220 26976 12232
rect 25179 12192 26976 12220
rect 25179 12189 25191 12192
rect 25133 12183 25191 12189
rect 26970 12180 26976 12192
rect 27028 12180 27034 12232
rect 27982 12220 27988 12232
rect 27943 12192 27988 12220
rect 27982 12180 27988 12192
rect 28040 12180 28046 12232
rect 28258 12220 28264 12232
rect 28219 12192 28264 12220
rect 28258 12180 28264 12192
rect 28316 12180 28322 12232
rect 29086 12180 29092 12232
rect 29144 12220 29150 12232
rect 29733 12223 29791 12229
rect 29733 12220 29745 12223
rect 29144 12192 29745 12220
rect 29144 12180 29150 12192
rect 29733 12189 29745 12192
rect 29779 12189 29791 12223
rect 29914 12220 29920 12232
rect 29875 12192 29920 12220
rect 29733 12183 29791 12189
rect 29914 12180 29920 12192
rect 29972 12180 29978 12232
rect 30098 12220 30104 12232
rect 30059 12192 30104 12220
rect 30098 12180 30104 12192
rect 30156 12180 30162 12232
rect 18196 12124 19748 12152
rect 19889 12155 19947 12161
rect 18196 12112 18202 12124
rect 19889 12121 19901 12155
rect 19935 12152 19947 12155
rect 21266 12152 21272 12164
rect 19935 12124 21272 12152
rect 19935 12121 19947 12124
rect 19889 12115 19947 12121
rect 21266 12112 21272 12124
rect 21324 12112 21330 12164
rect 21542 12112 21548 12164
rect 21600 12152 21606 12164
rect 21910 12152 21916 12164
rect 21600 12124 21916 12152
rect 21600 12112 21606 12124
rect 21910 12112 21916 12124
rect 21968 12112 21974 12164
rect 22005 12155 22063 12161
rect 22005 12121 22017 12155
rect 22051 12152 22063 12155
rect 22278 12152 22284 12164
rect 22051 12124 22284 12152
rect 22051 12121 22063 12124
rect 22005 12115 22063 12121
rect 22278 12112 22284 12124
rect 22336 12112 22342 12164
rect 24302 12112 24308 12164
rect 24360 12152 24366 12164
rect 24949 12155 25007 12161
rect 24949 12152 24961 12155
rect 24360 12124 24961 12152
rect 24360 12112 24366 12124
rect 24949 12121 24961 12124
rect 24995 12121 25007 12155
rect 24949 12115 25007 12121
rect 25777 12155 25835 12161
rect 25777 12121 25789 12155
rect 25823 12152 25835 12155
rect 27614 12152 27620 12164
rect 25823 12124 27620 12152
rect 25823 12121 25835 12124
rect 25777 12115 25835 12121
rect 27614 12112 27620 12124
rect 27672 12112 27678 12164
rect 29825 12155 29883 12161
rect 29825 12121 29837 12155
rect 29871 12121 29883 12155
rect 31956 12152 31984 12251
rect 32306 12180 32312 12232
rect 32364 12220 32370 12232
rect 32493 12223 32551 12229
rect 32493 12220 32505 12223
rect 32364 12192 32505 12220
rect 32364 12180 32370 12192
rect 32493 12189 32505 12192
rect 32539 12189 32551 12223
rect 32600 12220 32628 12328
rect 32674 12316 32680 12328
rect 32732 12316 32738 12368
rect 32766 12316 32772 12368
rect 32824 12316 32830 12368
rect 32781 12229 32809 12316
rect 32968 12288 32996 12396
rect 33134 12384 33140 12396
rect 33192 12384 33198 12436
rect 34514 12384 34520 12436
rect 34572 12424 34578 12436
rect 35342 12424 35348 12436
rect 34572 12396 35348 12424
rect 34572 12384 34578 12396
rect 35342 12384 35348 12396
rect 35400 12384 35406 12436
rect 34790 12288 34796 12300
rect 32968 12260 34796 12288
rect 34790 12248 34796 12260
rect 34848 12248 34854 12300
rect 35360 12288 35388 12384
rect 37093 12291 37151 12297
rect 35360 12260 35756 12288
rect 32656 12223 32714 12229
rect 32656 12220 32668 12223
rect 32600 12192 32668 12220
rect 32493 12183 32551 12189
rect 32656 12189 32668 12192
rect 32702 12189 32714 12223
rect 32656 12183 32714 12189
rect 32769 12223 32827 12229
rect 32769 12189 32781 12223
rect 32815 12189 32827 12223
rect 32769 12183 32827 12189
rect 32861 12223 32919 12229
rect 32861 12189 32873 12223
rect 32907 12189 32919 12223
rect 34808 12220 34836 12248
rect 35345 12223 35403 12229
rect 35345 12220 35357 12223
rect 34808 12192 35357 12220
rect 32861 12183 32919 12189
rect 35345 12189 35357 12192
rect 35391 12189 35403 12223
rect 35345 12183 35403 12189
rect 35437 12223 35495 12229
rect 35437 12189 35449 12223
rect 35483 12189 35495 12223
rect 35437 12183 35495 12189
rect 32876 12152 32904 12183
rect 31956 12124 32904 12152
rect 35452 12152 35480 12183
rect 35526 12180 35532 12232
rect 35584 12220 35590 12232
rect 35728 12229 35756 12260
rect 37093 12257 37105 12291
rect 37139 12288 37151 12291
rect 37274 12288 37280 12300
rect 37139 12260 37280 12288
rect 37139 12257 37151 12260
rect 37093 12251 37151 12257
rect 37274 12248 37280 12260
rect 37332 12248 37338 12300
rect 35713 12223 35771 12229
rect 35584 12192 35629 12220
rect 35584 12180 35590 12192
rect 35713 12189 35725 12223
rect 35759 12189 35771 12223
rect 35713 12183 35771 12189
rect 36817 12223 36875 12229
rect 36817 12189 36829 12223
rect 36863 12220 36875 12223
rect 37458 12220 37464 12232
rect 36863 12192 37464 12220
rect 36863 12189 36875 12192
rect 36817 12183 36875 12189
rect 37458 12180 37464 12192
rect 37516 12180 37522 12232
rect 37550 12180 37556 12232
rect 37608 12220 37614 12232
rect 37645 12223 37703 12229
rect 37645 12220 37657 12223
rect 37608 12192 37657 12220
rect 37608 12180 37614 12192
rect 37645 12189 37657 12192
rect 37691 12189 37703 12223
rect 37826 12220 37832 12232
rect 37787 12192 37832 12220
rect 37645 12183 37703 12189
rect 37826 12180 37832 12192
rect 37884 12180 37890 12232
rect 37921 12223 37979 12229
rect 37921 12189 37933 12223
rect 37967 12189 37979 12223
rect 37921 12183 37979 12189
rect 35986 12152 35992 12164
rect 35452 12124 35992 12152
rect 29825 12115 29883 12121
rect 13228 12056 15976 12084
rect 18693 12087 18751 12093
rect 13228 12044 13234 12056
rect 18693 12053 18705 12087
rect 18739 12084 18751 12087
rect 18966 12084 18972 12096
rect 18739 12056 18972 12084
rect 18739 12053 18751 12056
rect 18693 12047 18751 12053
rect 18966 12044 18972 12056
rect 19024 12044 19030 12096
rect 19334 12044 19340 12096
rect 19392 12084 19398 12096
rect 19518 12084 19524 12096
rect 19392 12056 19524 12084
rect 19392 12044 19398 12056
rect 19518 12044 19524 12056
rect 19576 12044 19582 12096
rect 20070 12084 20076 12096
rect 20031 12056 20076 12084
rect 20070 12044 20076 12056
rect 20128 12044 20134 12096
rect 24762 12044 24768 12096
rect 24820 12084 24826 12096
rect 25866 12084 25872 12096
rect 24820 12056 25872 12084
rect 24820 12044 24826 12056
rect 25866 12044 25872 12056
rect 25924 12044 25930 12096
rect 26234 12044 26240 12096
rect 26292 12084 26298 12096
rect 26510 12084 26516 12096
rect 26292 12056 26516 12084
rect 26292 12044 26298 12056
rect 26510 12044 26516 12056
rect 26568 12084 26574 12096
rect 27065 12087 27123 12093
rect 27065 12084 27077 12087
rect 26568 12056 27077 12084
rect 26568 12044 26574 12056
rect 27065 12053 27077 12056
rect 27111 12053 27123 12087
rect 28442 12084 28448 12096
rect 28403 12056 28448 12084
rect 27065 12047 27123 12053
rect 28442 12044 28448 12056
rect 28500 12044 28506 12096
rect 29178 12044 29184 12096
rect 29236 12084 29242 12096
rect 29549 12087 29607 12093
rect 29549 12084 29561 12087
rect 29236 12056 29561 12084
rect 29236 12044 29242 12056
rect 29549 12053 29561 12056
rect 29595 12053 29607 12087
rect 29840 12084 29868 12115
rect 35986 12112 35992 12124
rect 36044 12152 36050 12164
rect 37182 12152 37188 12164
rect 36044 12124 37188 12152
rect 36044 12112 36050 12124
rect 37182 12112 37188 12124
rect 37240 12152 37246 12164
rect 37936 12152 37964 12183
rect 38010 12180 38016 12232
rect 38068 12220 38074 12232
rect 38194 12220 38200 12232
rect 38068 12192 38200 12220
rect 38068 12180 38074 12192
rect 38194 12180 38200 12192
rect 38252 12220 38258 12232
rect 38749 12223 38807 12229
rect 38749 12220 38761 12223
rect 38252 12192 38761 12220
rect 38252 12180 38258 12192
rect 38749 12189 38761 12192
rect 38795 12189 38807 12223
rect 38749 12183 38807 12189
rect 40494 12180 40500 12232
rect 40552 12220 40558 12232
rect 41230 12220 41236 12232
rect 40552 12192 41236 12220
rect 40552 12180 40558 12192
rect 41230 12180 41236 12192
rect 41288 12180 41294 12232
rect 38102 12152 38108 12164
rect 37240 12124 38108 12152
rect 37240 12112 37246 12124
rect 38102 12112 38108 12124
rect 38160 12112 38166 12164
rect 38289 12155 38347 12161
rect 38289 12121 38301 12155
rect 38335 12152 38347 12155
rect 40966 12155 41024 12161
rect 40966 12152 40978 12155
rect 38335 12124 40978 12152
rect 38335 12121 38347 12124
rect 38289 12115 38347 12121
rect 40966 12121 40978 12124
rect 41012 12121 41024 12155
rect 40966 12115 41024 12121
rect 33410 12084 33416 12096
rect 29840 12056 33416 12084
rect 29549 12047 29607 12053
rect 33410 12044 33416 12056
rect 33468 12044 33474 12096
rect 35066 12084 35072 12096
rect 35027 12056 35072 12084
rect 35066 12044 35072 12056
rect 35124 12044 35130 12096
rect 38654 12044 38660 12096
rect 38712 12084 38718 12096
rect 39853 12087 39911 12093
rect 39853 12084 39865 12087
rect 38712 12056 39865 12084
rect 38712 12044 38718 12056
rect 39853 12053 39865 12056
rect 39899 12053 39911 12087
rect 39853 12047 39911 12053
rect 1104 11994 68816 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 68816 11994
rect 1104 11920 68816 11942
rect 5445 11883 5503 11889
rect 5445 11849 5457 11883
rect 5491 11880 5503 11883
rect 6638 11880 6644 11892
rect 5491 11852 6644 11880
rect 5491 11849 5503 11852
rect 5445 11843 5503 11849
rect 6638 11840 6644 11852
rect 6696 11840 6702 11892
rect 13354 11840 13360 11892
rect 13412 11880 13418 11892
rect 13449 11883 13507 11889
rect 13449 11880 13461 11883
rect 13412 11852 13461 11880
rect 13412 11840 13418 11852
rect 13449 11849 13461 11852
rect 13495 11849 13507 11883
rect 14182 11880 14188 11892
rect 14143 11852 14188 11880
rect 13449 11843 13507 11849
rect 14182 11840 14188 11852
rect 14240 11840 14246 11892
rect 14921 11883 14979 11889
rect 14921 11849 14933 11883
rect 14967 11880 14979 11883
rect 14967 11852 16160 11880
rect 14967 11849 14979 11852
rect 14921 11843 14979 11849
rect 2593 11815 2651 11821
rect 2593 11781 2605 11815
rect 2639 11812 2651 11815
rect 3390 11815 3448 11821
rect 3390 11812 3402 11815
rect 2639 11784 3402 11812
rect 2639 11781 2651 11784
rect 2593 11775 2651 11781
rect 3390 11781 3402 11784
rect 3436 11781 3448 11815
rect 3390 11775 3448 11781
rect 5166 11772 5172 11824
rect 5224 11812 5230 11824
rect 5629 11815 5687 11821
rect 5629 11812 5641 11815
rect 5224 11784 5641 11812
rect 5224 11772 5230 11784
rect 5629 11781 5641 11784
rect 5675 11812 5687 11815
rect 12621 11815 12679 11821
rect 12621 11812 12633 11815
rect 5675 11784 11560 11812
rect 5675 11781 5687 11784
rect 5629 11775 5687 11781
rect 1762 11704 1768 11756
rect 1820 11744 1826 11756
rect 1949 11747 2007 11753
rect 1949 11744 1961 11747
rect 1820 11716 1961 11744
rect 1820 11704 1826 11716
rect 1949 11713 1961 11716
rect 1995 11713 2007 11747
rect 2130 11744 2136 11756
rect 2091 11716 2136 11744
rect 1949 11707 2007 11713
rect 2130 11704 2136 11716
rect 2188 11704 2194 11756
rect 2222 11704 2228 11756
rect 2280 11744 2286 11756
rect 2363 11747 2421 11753
rect 2280 11716 2325 11744
rect 2280 11704 2286 11716
rect 2363 11713 2375 11747
rect 2409 11744 2421 11747
rect 2774 11744 2780 11756
rect 2409 11716 2780 11744
rect 2409 11713 2421 11716
rect 2363 11707 2421 11713
rect 2774 11704 2780 11716
rect 2832 11704 2838 11756
rect 5810 11744 5816 11756
rect 5771 11716 5816 11744
rect 5810 11704 5816 11716
rect 5868 11704 5874 11756
rect 6730 11744 6736 11756
rect 6643 11716 6736 11744
rect 6730 11704 6736 11716
rect 6788 11744 6794 11756
rect 8941 11747 8999 11753
rect 8941 11744 8953 11747
rect 6788 11716 8953 11744
rect 6788 11704 6794 11716
rect 8941 11713 8953 11716
rect 8987 11713 8999 11747
rect 10410 11744 10416 11756
rect 10371 11716 10416 11744
rect 8941 11707 8999 11713
rect 10410 11704 10416 11716
rect 10468 11704 10474 11756
rect 11532 11753 11560 11784
rect 12406 11784 12633 11812
rect 11517 11747 11575 11753
rect 11517 11713 11529 11747
rect 11563 11713 11575 11747
rect 11698 11744 11704 11756
rect 11611 11716 11704 11744
rect 11517 11707 11575 11713
rect 11698 11704 11704 11716
rect 11756 11704 11762 11756
rect 11793 11747 11851 11753
rect 11793 11713 11805 11747
rect 11839 11713 11851 11747
rect 11793 11707 11851 11713
rect 3142 11676 3148 11688
rect 3103 11648 3148 11676
rect 3142 11636 3148 11648
rect 3200 11636 3206 11688
rect 6362 11636 6368 11688
rect 6420 11676 6426 11688
rect 9490 11676 9496 11688
rect 6420 11648 9496 11676
rect 6420 11636 6426 11648
rect 9490 11636 9496 11648
rect 9548 11636 9554 11688
rect 10137 11679 10195 11685
rect 10137 11645 10149 11679
rect 10183 11676 10195 11679
rect 11716 11676 11744 11704
rect 10183 11648 11744 11676
rect 10183 11645 10195 11648
rect 10137 11639 10195 11645
rect 4525 11611 4583 11617
rect 4525 11577 4537 11611
rect 4571 11608 4583 11611
rect 11808 11608 11836 11707
rect 11882 11704 11888 11756
rect 11940 11744 11946 11756
rect 12406 11744 12434 11784
rect 12621 11781 12633 11784
rect 12667 11781 12679 11815
rect 12621 11775 12679 11781
rect 11940 11716 12434 11744
rect 12529 11747 12587 11753
rect 11940 11704 11946 11716
rect 12529 11713 12541 11747
rect 12575 11713 12587 11747
rect 12529 11707 12587 11713
rect 12713 11747 12771 11753
rect 12713 11713 12725 11747
rect 12759 11744 12771 11747
rect 12894 11744 12900 11756
rect 12759 11716 12900 11744
rect 12759 11713 12771 11716
rect 12713 11707 12771 11713
rect 12544 11676 12572 11707
rect 12894 11704 12900 11716
rect 12952 11704 12958 11756
rect 13633 11747 13691 11753
rect 13633 11713 13645 11747
rect 13679 11713 13691 11747
rect 13633 11707 13691 11713
rect 13170 11676 13176 11688
rect 12544 11648 13176 11676
rect 13170 11636 13176 11648
rect 13228 11636 13234 11688
rect 13648 11676 13676 11707
rect 13722 11704 13728 11756
rect 13780 11744 13786 11756
rect 14369 11747 14427 11753
rect 14369 11744 14381 11747
rect 13780 11716 14381 11744
rect 13780 11704 13786 11716
rect 14369 11713 14381 11716
rect 14415 11744 14427 11747
rect 14936 11744 14964 11843
rect 15838 11812 15844 11824
rect 15799 11784 15844 11812
rect 15838 11772 15844 11784
rect 15896 11772 15902 11824
rect 14415 11716 14964 11744
rect 16025 11747 16083 11753
rect 14415 11713 14427 11716
rect 14369 11707 14427 11713
rect 16025 11713 16037 11747
rect 16071 11713 16083 11747
rect 16025 11707 16083 11713
rect 16040 11676 16068 11707
rect 13648 11648 16068 11676
rect 16132 11676 16160 11852
rect 16390 11840 16396 11892
rect 16448 11880 16454 11892
rect 21266 11880 21272 11892
rect 16448 11852 20300 11880
rect 21227 11852 21272 11880
rect 16448 11840 16454 11852
rect 17862 11772 17868 11824
rect 17920 11812 17926 11824
rect 18325 11815 18383 11821
rect 18325 11812 18337 11815
rect 17920 11784 18337 11812
rect 17920 11772 17926 11784
rect 18325 11781 18337 11784
rect 18371 11812 18383 11815
rect 19702 11812 19708 11824
rect 18371 11784 19708 11812
rect 18371 11781 18383 11784
rect 18325 11775 18383 11781
rect 19702 11772 19708 11784
rect 19760 11772 19766 11824
rect 19794 11772 19800 11824
rect 19852 11812 19858 11824
rect 20134 11815 20192 11821
rect 20134 11812 20146 11815
rect 19852 11784 20146 11812
rect 19852 11772 19858 11784
rect 20134 11781 20146 11784
rect 20180 11781 20192 11815
rect 20272 11812 20300 11852
rect 21266 11840 21272 11852
rect 21324 11840 21330 11892
rect 22094 11840 22100 11892
rect 22152 11880 22158 11892
rect 22465 11883 22523 11889
rect 22465 11880 22477 11883
rect 22152 11852 22477 11880
rect 22152 11840 22158 11852
rect 22465 11849 22477 11852
rect 22511 11880 22523 11883
rect 22511 11852 24532 11880
rect 22511 11849 22523 11852
rect 22465 11843 22523 11849
rect 22186 11812 22192 11824
rect 20272 11784 22192 11812
rect 20134 11775 20192 11781
rect 22186 11772 22192 11784
rect 22244 11772 22250 11824
rect 24504 11821 24532 11852
rect 25498 11840 25504 11892
rect 25556 11840 25562 11892
rect 26786 11840 26792 11892
rect 26844 11880 26850 11892
rect 27433 11883 27491 11889
rect 27433 11880 27445 11883
rect 26844 11852 27445 11880
rect 26844 11840 26850 11852
rect 27433 11849 27445 11852
rect 27479 11849 27491 11883
rect 27433 11843 27491 11849
rect 27522 11840 27528 11892
rect 27580 11880 27586 11892
rect 28166 11880 28172 11892
rect 27580 11852 28172 11880
rect 27580 11840 27586 11852
rect 28166 11840 28172 11852
rect 28224 11840 28230 11892
rect 32122 11880 32128 11892
rect 29288 11852 32128 11880
rect 24489 11815 24547 11821
rect 24489 11781 24501 11815
rect 24535 11781 24547 11815
rect 24489 11775 24547 11781
rect 25038 11772 25044 11824
rect 25096 11812 25102 11824
rect 25516 11812 25544 11840
rect 29288 11812 29316 11852
rect 32122 11840 32128 11852
rect 32180 11840 32186 11892
rect 32306 11840 32312 11892
rect 32364 11880 32370 11892
rect 34057 11883 34115 11889
rect 32364 11852 32904 11880
rect 32364 11840 32370 11852
rect 29454 11812 29460 11824
rect 25096 11784 25636 11812
rect 25096 11772 25102 11784
rect 18138 11744 18144 11756
rect 18099 11716 18144 11744
rect 18138 11704 18144 11716
rect 18196 11704 18202 11756
rect 19886 11744 19892 11756
rect 19847 11716 19892 11744
rect 19886 11704 19892 11716
rect 19944 11704 19950 11756
rect 21450 11744 21456 11756
rect 19996 11716 21456 11744
rect 18874 11676 18880 11688
rect 16132 11648 18880 11676
rect 12066 11608 12072 11620
rect 4571 11580 11836 11608
rect 12027 11580 12072 11608
rect 4571 11577 4583 11580
rect 4525 11571 4583 11577
rect 2498 11500 2504 11552
rect 2556 11540 2562 11552
rect 4540 11540 4568 11571
rect 12066 11568 12072 11580
rect 12124 11568 12130 11620
rect 2556 11512 4568 11540
rect 2556 11500 2562 11512
rect 7558 11500 7564 11552
rect 7616 11540 7622 11552
rect 8021 11543 8079 11549
rect 8021 11540 8033 11543
rect 7616 11512 8033 11540
rect 7616 11500 7622 11512
rect 8021 11509 8033 11512
rect 8067 11509 8079 11543
rect 8021 11503 8079 11509
rect 9490 11500 9496 11552
rect 9548 11540 9554 11552
rect 13354 11540 13360 11552
rect 9548 11512 13360 11540
rect 9548 11500 9554 11512
rect 13354 11500 13360 11512
rect 13412 11500 13418 11552
rect 15838 11500 15844 11552
rect 15896 11540 15902 11552
rect 16040 11540 16068 11648
rect 18874 11636 18880 11648
rect 18932 11636 18938 11688
rect 18966 11636 18972 11688
rect 19024 11676 19030 11688
rect 19996 11676 20024 11716
rect 21450 11704 21456 11716
rect 21508 11704 21514 11756
rect 23589 11747 23647 11753
rect 23589 11713 23601 11747
rect 23635 11744 23647 11747
rect 24210 11744 24216 11756
rect 23635 11716 24216 11744
rect 23635 11713 23647 11716
rect 23589 11707 23647 11713
rect 24210 11704 24216 11716
rect 24268 11704 24274 11756
rect 24302 11704 24308 11756
rect 24360 11744 24366 11756
rect 25314 11744 25320 11756
rect 24360 11716 24405 11744
rect 25275 11716 25320 11744
rect 24360 11704 24366 11716
rect 25314 11704 25320 11716
rect 25372 11704 25378 11756
rect 25498 11744 25504 11756
rect 25459 11716 25504 11744
rect 25498 11704 25504 11716
rect 25556 11704 25562 11756
rect 25608 11753 25636 11784
rect 27264 11784 29316 11812
rect 29415 11784 29460 11812
rect 25593 11747 25651 11753
rect 25593 11713 25605 11747
rect 25639 11713 25651 11747
rect 25593 11707 25651 11713
rect 25682 11704 25688 11756
rect 25740 11744 25746 11756
rect 26970 11744 26976 11756
rect 25740 11716 25785 11744
rect 26931 11716 26976 11744
rect 25740 11704 25746 11716
rect 26970 11704 26976 11716
rect 27028 11704 27034 11756
rect 27264 11753 27292 11784
rect 29454 11772 29460 11784
rect 29512 11772 29518 11824
rect 29549 11815 29607 11821
rect 29549 11781 29561 11815
rect 29595 11812 29607 11815
rect 29914 11812 29920 11824
rect 29595 11784 29920 11812
rect 29595 11781 29607 11784
rect 29549 11775 29607 11781
rect 29914 11772 29920 11784
rect 29972 11772 29978 11824
rect 31328 11815 31386 11821
rect 31328 11781 31340 11815
rect 31374 11812 31386 11815
rect 32217 11815 32275 11821
rect 32217 11812 32229 11815
rect 31374 11784 32229 11812
rect 31374 11781 31386 11784
rect 31328 11775 31386 11781
rect 32217 11781 32229 11784
rect 32263 11781 32275 11815
rect 32766 11812 32772 11824
rect 32217 11775 32275 11781
rect 32600 11784 32772 11812
rect 27249 11747 27307 11753
rect 27249 11713 27261 11747
rect 27295 11713 27307 11747
rect 27249 11707 27307 11713
rect 27890 11704 27896 11756
rect 27948 11744 27954 11756
rect 27985 11747 28043 11753
rect 27985 11744 27997 11747
rect 27948 11716 27997 11744
rect 27948 11704 27954 11716
rect 27985 11713 27997 11716
rect 28031 11744 28043 11747
rect 28629 11747 28687 11753
rect 28629 11744 28641 11747
rect 28031 11716 28641 11744
rect 28031 11713 28043 11716
rect 27985 11707 28043 11713
rect 28629 11713 28641 11716
rect 28675 11713 28687 11747
rect 28629 11707 28687 11713
rect 29086 11704 29092 11756
rect 29144 11744 29150 11756
rect 29362 11744 29368 11756
rect 29144 11716 29368 11744
rect 29144 11704 29150 11716
rect 29362 11704 29368 11716
rect 29420 11704 29426 11756
rect 29733 11747 29791 11753
rect 29733 11713 29745 11747
rect 29779 11744 29791 11747
rect 30466 11744 30472 11756
rect 29779 11716 30472 11744
rect 29779 11713 29791 11716
rect 29733 11707 29791 11713
rect 30466 11704 30472 11716
rect 30524 11704 30530 11756
rect 31573 11747 31631 11753
rect 31573 11713 31585 11747
rect 31619 11744 31631 11747
rect 31938 11744 31944 11756
rect 31619 11716 31944 11744
rect 31619 11713 31631 11716
rect 31573 11707 31631 11713
rect 31938 11704 31944 11716
rect 31996 11704 32002 11756
rect 32490 11744 32496 11756
rect 32451 11716 32496 11744
rect 32490 11704 32496 11716
rect 32548 11704 32554 11756
rect 32600 11753 32628 11784
rect 32766 11772 32772 11784
rect 32824 11772 32830 11824
rect 32585 11747 32643 11753
rect 32585 11713 32597 11747
rect 32631 11713 32643 11747
rect 32585 11707 32643 11713
rect 32674 11704 32680 11756
rect 32732 11744 32738 11756
rect 32876 11753 32904 11852
rect 34057 11849 34069 11883
rect 34103 11880 34115 11883
rect 35710 11880 35716 11892
rect 34103 11852 35716 11880
rect 34103 11849 34115 11852
rect 34057 11843 34115 11849
rect 35710 11840 35716 11852
rect 35768 11840 35774 11892
rect 37366 11880 37372 11892
rect 36372 11852 37372 11880
rect 35066 11772 35072 11824
rect 35124 11812 35130 11824
rect 35170 11815 35228 11821
rect 35170 11812 35182 11815
rect 35124 11784 35182 11812
rect 35124 11772 35130 11784
rect 35170 11781 35182 11784
rect 35216 11781 35228 11815
rect 35170 11775 35228 11781
rect 36372 11753 36400 11852
rect 37366 11840 37372 11852
rect 37424 11840 37430 11892
rect 36464 11784 40540 11812
rect 32861 11747 32919 11753
rect 32732 11716 32777 11744
rect 32732 11704 32738 11716
rect 32861 11713 32873 11747
rect 32907 11713 32919 11747
rect 32861 11707 32919 11713
rect 35437 11747 35495 11753
rect 35437 11713 35449 11747
rect 35483 11713 35495 11747
rect 35437 11707 35495 11713
rect 36357 11747 36415 11753
rect 36357 11713 36369 11747
rect 36403 11713 36415 11747
rect 36357 11707 36415 11713
rect 19024 11648 20024 11676
rect 19024 11636 19030 11648
rect 23842 11636 23848 11688
rect 23900 11676 23906 11688
rect 26510 11676 26516 11688
rect 23900 11648 26516 11676
rect 23900 11636 23906 11648
rect 26510 11636 26516 11648
rect 26568 11636 26574 11688
rect 27062 11676 27068 11688
rect 27023 11648 27068 11676
rect 27062 11636 27068 11648
rect 27120 11636 27126 11688
rect 35452 11676 35480 11707
rect 36464 11676 36492 11784
rect 40512 11756 40540 11784
rect 36541 11747 36599 11753
rect 36541 11713 36553 11747
rect 36587 11719 36676 11747
rect 36587 11713 36599 11719
rect 36541 11707 36599 11713
rect 35452 11648 36492 11676
rect 28166 11608 28172 11620
rect 28127 11580 28172 11608
rect 28166 11568 28172 11580
rect 28224 11568 28230 11620
rect 28258 11568 28264 11620
rect 28316 11608 28322 11620
rect 36648 11608 36676 11719
rect 37458 11704 37464 11756
rect 37516 11744 37522 11756
rect 37645 11747 37703 11753
rect 37516 11716 37561 11744
rect 37516 11704 37522 11716
rect 37645 11713 37657 11747
rect 37691 11713 37703 11747
rect 37645 11707 37703 11713
rect 37737 11747 37795 11753
rect 37737 11713 37749 11747
rect 37783 11713 37795 11747
rect 37737 11707 37795 11713
rect 37829 11747 37887 11753
rect 37829 11713 37841 11747
rect 37875 11744 37887 11747
rect 38010 11744 38016 11756
rect 37875 11716 38016 11744
rect 37875 11713 37887 11716
rect 37829 11707 37887 11713
rect 36725 11679 36783 11685
rect 36725 11645 36737 11679
rect 36771 11676 36783 11679
rect 37660 11676 37688 11707
rect 36771 11648 37688 11676
rect 37752 11676 37780 11707
rect 38010 11704 38016 11716
rect 38068 11704 38074 11756
rect 40230 11747 40288 11753
rect 40230 11744 40242 11747
rect 38120 11716 40242 11744
rect 37918 11676 37924 11688
rect 37752 11648 37924 11676
rect 36771 11645 36783 11648
rect 36725 11639 36783 11645
rect 37918 11636 37924 11648
rect 37976 11636 37982 11688
rect 38120 11685 38148 11716
rect 40230 11713 40242 11716
rect 40276 11713 40288 11747
rect 40494 11744 40500 11756
rect 40407 11716 40500 11744
rect 40230 11707 40288 11713
rect 40494 11704 40500 11716
rect 40552 11704 40558 11756
rect 38105 11679 38163 11685
rect 38105 11645 38117 11679
rect 38151 11645 38163 11679
rect 38105 11639 38163 11645
rect 67634 11608 67640 11620
rect 28316 11580 30420 11608
rect 36648 11580 37320 11608
rect 67595 11580 67640 11608
rect 28316 11568 28322 11580
rect 16669 11543 16727 11549
rect 16669 11540 16681 11543
rect 15896 11512 16681 11540
rect 15896 11500 15902 11512
rect 16669 11509 16681 11512
rect 16715 11509 16727 11543
rect 16669 11503 16727 11509
rect 17034 11500 17040 11552
rect 17092 11540 17098 11552
rect 17589 11543 17647 11549
rect 17589 11540 17601 11543
rect 17092 11512 17601 11540
rect 17092 11500 17098 11512
rect 17589 11509 17601 11512
rect 17635 11509 17647 11543
rect 18506 11540 18512 11552
rect 18467 11512 18512 11540
rect 17589 11503 17647 11509
rect 18506 11500 18512 11512
rect 18564 11500 18570 11552
rect 19337 11543 19395 11549
rect 19337 11509 19349 11543
rect 19383 11540 19395 11543
rect 20162 11540 20168 11552
rect 19383 11512 20168 11540
rect 19383 11509 19395 11512
rect 19337 11503 19395 11509
rect 20162 11500 20168 11512
rect 20220 11500 20226 11552
rect 21266 11500 21272 11552
rect 21324 11540 21330 11552
rect 22370 11540 22376 11552
rect 21324 11512 22376 11540
rect 21324 11500 21330 11512
rect 22370 11500 22376 11512
rect 22428 11500 22434 11552
rect 24673 11543 24731 11549
rect 24673 11509 24685 11543
rect 24719 11540 24731 11543
rect 25130 11540 25136 11552
rect 24719 11512 25136 11540
rect 24719 11509 24731 11512
rect 24673 11503 24731 11509
rect 25130 11500 25136 11512
rect 25188 11500 25194 11552
rect 25961 11543 26019 11549
rect 25961 11509 25973 11543
rect 26007 11540 26019 11543
rect 26602 11540 26608 11552
rect 26007 11512 26608 11540
rect 26007 11509 26019 11512
rect 25961 11503 26019 11509
rect 26602 11500 26608 11512
rect 26660 11500 26666 11552
rect 27249 11543 27307 11549
rect 27249 11509 27261 11543
rect 27295 11540 27307 11543
rect 27338 11540 27344 11552
rect 27295 11512 27344 11540
rect 27295 11509 27307 11512
rect 27249 11503 27307 11509
rect 27338 11500 27344 11512
rect 27396 11500 27402 11552
rect 27798 11500 27804 11552
rect 27856 11540 27862 11552
rect 28534 11540 28540 11552
rect 27856 11512 28540 11540
rect 27856 11500 27862 11512
rect 28534 11500 28540 11512
rect 28592 11500 28598 11552
rect 29086 11500 29092 11552
rect 29144 11540 29150 11552
rect 29181 11543 29239 11549
rect 29181 11540 29193 11543
rect 29144 11512 29193 11540
rect 29144 11500 29150 11512
rect 29181 11509 29193 11512
rect 29227 11509 29239 11543
rect 29181 11503 29239 11509
rect 30193 11543 30251 11549
rect 30193 11509 30205 11543
rect 30239 11540 30251 11543
rect 30282 11540 30288 11552
rect 30239 11512 30288 11540
rect 30239 11509 30251 11512
rect 30193 11503 30251 11509
rect 30282 11500 30288 11512
rect 30340 11500 30346 11552
rect 30392 11540 30420 11580
rect 37292 11552 37320 11580
rect 67634 11568 67640 11580
rect 67692 11568 67698 11620
rect 36906 11540 36912 11552
rect 30392 11512 36912 11540
rect 36906 11500 36912 11512
rect 36964 11500 36970 11552
rect 37274 11500 37280 11552
rect 37332 11540 37338 11552
rect 39117 11543 39175 11549
rect 39117 11540 39129 11543
rect 37332 11512 39129 11540
rect 37332 11500 37338 11512
rect 39117 11509 39129 11512
rect 39163 11509 39175 11543
rect 39117 11503 39175 11509
rect 1104 11450 68816 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 65654 11450
rect 65706 11398 65718 11450
rect 65770 11398 65782 11450
rect 65834 11398 65846 11450
rect 65898 11398 65910 11450
rect 65962 11398 68816 11450
rect 1104 11376 68816 11398
rect 1949 11339 2007 11345
rect 1949 11305 1961 11339
rect 1995 11336 2007 11339
rect 2130 11336 2136 11348
rect 1995 11308 2136 11336
rect 1995 11305 2007 11308
rect 1949 11299 2007 11305
rect 2130 11296 2136 11308
rect 2188 11296 2194 11348
rect 2774 11336 2780 11348
rect 2735 11308 2780 11336
rect 2774 11296 2780 11308
rect 2832 11296 2838 11348
rect 5166 11336 5172 11348
rect 5127 11308 5172 11336
rect 5166 11296 5172 11308
rect 5224 11296 5230 11348
rect 7193 11339 7251 11345
rect 7193 11305 7205 11339
rect 7239 11336 7251 11339
rect 7926 11336 7932 11348
rect 7239 11308 7932 11336
rect 7239 11305 7251 11308
rect 7193 11299 7251 11305
rect 7926 11296 7932 11308
rect 7984 11296 7990 11348
rect 13357 11339 13415 11345
rect 13357 11305 13369 11339
rect 13403 11336 13415 11339
rect 13446 11336 13452 11348
rect 13403 11308 13452 11336
rect 13403 11305 13415 11308
rect 13357 11299 13415 11305
rect 13446 11296 13452 11308
rect 13504 11296 13510 11348
rect 16390 11336 16396 11348
rect 14476 11308 16396 11336
rect 12434 11228 12440 11280
rect 12492 11268 12498 11280
rect 12529 11271 12587 11277
rect 12529 11268 12541 11271
rect 12492 11240 12541 11268
rect 12492 11228 12498 11240
rect 12529 11237 12541 11240
rect 12575 11268 12587 11271
rect 14476 11268 14504 11308
rect 16390 11296 16396 11308
rect 16448 11296 16454 11348
rect 17773 11339 17831 11345
rect 17773 11305 17785 11339
rect 17819 11336 17831 11339
rect 17862 11336 17868 11348
rect 17819 11308 17868 11336
rect 17819 11305 17831 11308
rect 17773 11299 17831 11305
rect 17862 11296 17868 11308
rect 17920 11296 17926 11348
rect 18414 11336 18420 11348
rect 18375 11308 18420 11336
rect 18414 11296 18420 11308
rect 18472 11296 18478 11348
rect 19794 11296 19800 11348
rect 19852 11336 19858 11348
rect 20349 11339 20407 11345
rect 20349 11336 20361 11339
rect 19852 11308 20361 11336
rect 19852 11296 19858 11308
rect 20349 11305 20361 11308
rect 20395 11305 20407 11339
rect 20349 11299 20407 11305
rect 22005 11339 22063 11345
rect 22005 11305 22017 11339
rect 22051 11336 22063 11339
rect 22186 11336 22192 11348
rect 22051 11308 22192 11336
rect 22051 11305 22063 11308
rect 22005 11299 22063 11305
rect 22186 11296 22192 11308
rect 22244 11296 22250 11348
rect 23845 11339 23903 11345
rect 23845 11305 23857 11339
rect 23891 11336 23903 11339
rect 23934 11336 23940 11348
rect 23891 11308 23940 11336
rect 23891 11305 23903 11308
rect 23845 11299 23903 11305
rect 23934 11296 23940 11308
rect 23992 11296 23998 11348
rect 24210 11296 24216 11348
rect 24268 11336 24274 11348
rect 24673 11339 24731 11345
rect 24673 11336 24685 11339
rect 24268 11308 24685 11336
rect 24268 11296 24274 11308
rect 24673 11305 24685 11308
rect 24719 11305 24731 11339
rect 24673 11299 24731 11305
rect 24854 11296 24860 11348
rect 24912 11336 24918 11348
rect 25590 11336 25596 11348
rect 24912 11308 25596 11336
rect 24912 11296 24918 11308
rect 25590 11296 25596 11308
rect 25648 11296 25654 11348
rect 25682 11296 25688 11348
rect 25740 11336 25746 11348
rect 25777 11339 25835 11345
rect 25777 11336 25789 11339
rect 25740 11308 25789 11336
rect 25740 11296 25746 11308
rect 25777 11305 25789 11308
rect 25823 11305 25835 11339
rect 25777 11299 25835 11305
rect 26142 11296 26148 11348
rect 26200 11336 26206 11348
rect 27893 11339 27951 11345
rect 27893 11336 27905 11339
rect 26200 11308 27905 11336
rect 26200 11296 26206 11308
rect 27893 11305 27905 11308
rect 27939 11305 27951 11339
rect 27893 11299 27951 11305
rect 19886 11268 19892 11280
rect 12575 11240 14504 11268
rect 18708 11240 19892 11268
rect 12575 11237 12587 11240
rect 12529 11231 12587 11237
rect 8386 11200 8392 11212
rect 7576 11172 8392 11200
rect 7576 11144 7604 11172
rect 8386 11160 8392 11172
rect 8444 11200 8450 11212
rect 8941 11203 8999 11209
rect 8941 11200 8953 11203
rect 8444 11172 8953 11200
rect 8444 11160 8450 11172
rect 8941 11169 8953 11172
rect 8987 11169 8999 11203
rect 8941 11163 8999 11169
rect 11977 11203 12035 11209
rect 11977 11169 11989 11203
rect 12023 11200 12035 11203
rect 18708 11200 18736 11240
rect 19886 11228 19892 11240
rect 19944 11228 19950 11280
rect 20070 11268 20076 11280
rect 19996 11240 20076 11268
rect 19610 11200 19616 11212
rect 12023 11172 13216 11200
rect 12023 11169 12035 11172
rect 11977 11163 12035 11169
rect 2133 11135 2191 11141
rect 2133 11101 2145 11135
rect 2179 11132 2191 11135
rect 2498 11132 2504 11144
rect 2179 11104 2504 11132
rect 2179 11101 2191 11104
rect 2133 11095 2191 11101
rect 2498 11092 2504 11104
rect 2556 11092 2562 11144
rect 3142 11092 3148 11144
rect 3200 11132 3206 11144
rect 6549 11135 6607 11141
rect 6549 11132 6561 11135
rect 3200 11104 6561 11132
rect 3200 11092 3206 11104
rect 6549 11101 6561 11104
rect 6595 11132 6607 11135
rect 7558 11132 7564 11144
rect 6595 11104 7564 11132
rect 6595 11101 6607 11104
rect 6549 11095 6607 11101
rect 7558 11092 7564 11104
rect 7616 11092 7622 11144
rect 7653 11135 7711 11141
rect 7653 11101 7665 11135
rect 7699 11101 7711 11135
rect 7653 11095 7711 11101
rect 2314 11064 2320 11076
rect 2275 11036 2320 11064
rect 2314 11024 2320 11036
rect 2372 11024 2378 11076
rect 6178 11024 6184 11076
rect 6236 11064 6242 11076
rect 6282 11067 6340 11073
rect 6282 11064 6294 11067
rect 6236 11036 6294 11064
rect 6236 11024 6242 11036
rect 6282 11033 6294 11036
rect 6328 11033 6340 11067
rect 6282 11027 6340 11033
rect 7006 11024 7012 11076
rect 7064 11064 7070 11076
rect 7668 11064 7696 11095
rect 7742 11092 7748 11144
rect 7800 11132 7806 11144
rect 7837 11135 7895 11141
rect 7837 11132 7849 11135
rect 7800 11104 7849 11132
rect 7800 11092 7806 11104
rect 7837 11101 7849 11104
rect 7883 11101 7895 11135
rect 7837 11095 7895 11101
rect 7926 11092 7932 11144
rect 7984 11132 7990 11144
rect 8067 11135 8125 11141
rect 7984 11104 8029 11132
rect 7984 11092 7990 11104
rect 8067 11101 8079 11135
rect 8113 11132 8125 11135
rect 8754 11132 8760 11144
rect 8113 11104 8760 11132
rect 8113 11101 8125 11104
rect 8067 11095 8125 11101
rect 8754 11092 8760 11104
rect 8812 11092 8818 11144
rect 13188 11141 13216 11172
rect 18432 11172 18736 11200
rect 19306 11172 19616 11200
rect 12713 11135 12771 11141
rect 12713 11101 12725 11135
rect 12759 11101 12771 11135
rect 12713 11095 12771 11101
rect 13173 11135 13231 11141
rect 13173 11101 13185 11135
rect 13219 11132 13231 11135
rect 13722 11132 13728 11144
rect 13219 11104 13728 11132
rect 13219 11101 13231 11104
rect 13173 11095 13231 11101
rect 7064 11036 7696 11064
rect 8297 11067 8355 11073
rect 7064 11024 7070 11036
rect 8297 11033 8309 11067
rect 8343 11064 8355 11067
rect 9186 11067 9244 11073
rect 9186 11064 9198 11067
rect 8343 11036 9198 11064
rect 8343 11033 8355 11036
rect 8297 11027 8355 11033
rect 9186 11033 9198 11036
rect 9232 11033 9244 11067
rect 12728 11064 12756 11095
rect 13722 11092 13728 11104
rect 13780 11092 13786 11144
rect 15749 11135 15807 11141
rect 15749 11101 15761 11135
rect 15795 11132 15807 11135
rect 16393 11135 16451 11141
rect 16393 11132 16405 11135
rect 15795 11104 16405 11132
rect 15795 11101 15807 11104
rect 15749 11095 15807 11101
rect 16393 11101 16405 11104
rect 16439 11132 16451 11135
rect 18432 11132 18460 11172
rect 16439 11104 18460 11132
rect 18509 11135 18567 11141
rect 16439 11101 16451 11104
rect 16393 11095 16451 11101
rect 18509 11101 18521 11135
rect 18555 11101 18567 11135
rect 18509 11095 18567 11101
rect 18601 11135 18659 11141
rect 18601 11101 18613 11135
rect 18647 11132 18659 11135
rect 19306 11132 19334 11172
rect 19610 11160 19616 11172
rect 19668 11160 19674 11212
rect 19794 11160 19800 11212
rect 19852 11160 19858 11212
rect 18647 11104 19334 11132
rect 18647 11101 18659 11104
rect 18601 11095 18659 11101
rect 13262 11064 13268 11076
rect 9186 11027 9244 11033
rect 10060 11036 10456 11064
rect 12728 11036 13268 11064
rect 9030 10956 9036 11008
rect 9088 10996 9094 11008
rect 10060 10996 10088 11036
rect 9088 10968 10088 10996
rect 9088 10956 9094 10968
rect 10134 10956 10140 11008
rect 10192 10996 10198 11008
rect 10321 10999 10379 11005
rect 10321 10996 10333 10999
rect 10192 10968 10333 10996
rect 10192 10956 10198 10968
rect 10321 10965 10333 10968
rect 10367 10965 10379 10999
rect 10428 10996 10456 11036
rect 13262 11024 13268 11036
rect 13320 11024 13326 11076
rect 15194 11024 15200 11076
rect 15252 11064 15258 11076
rect 15482 11067 15540 11073
rect 15482 11064 15494 11067
rect 15252 11036 15494 11064
rect 15252 11024 15258 11036
rect 15482 11033 15494 11036
rect 15528 11033 15540 11067
rect 15482 11027 15540 11033
rect 16660 11067 16718 11073
rect 16660 11033 16672 11067
rect 16706 11064 16718 11067
rect 18046 11064 18052 11076
rect 16706 11036 18052 11064
rect 16706 11033 16718 11036
rect 16660 11027 16718 11033
rect 18046 11024 18052 11036
rect 18104 11024 18110 11076
rect 18524 11064 18552 11095
rect 19426 11092 19432 11144
rect 19484 11132 19490 11144
rect 19705 11135 19763 11141
rect 19705 11132 19717 11135
rect 19484 11104 19717 11132
rect 19484 11092 19490 11104
rect 19705 11101 19717 11104
rect 19751 11101 19763 11135
rect 19705 11095 19763 11101
rect 19812 11126 19840 11160
rect 19996 11141 20024 11240
rect 20070 11228 20076 11240
rect 20128 11228 20134 11280
rect 20162 11228 20168 11280
rect 20220 11268 20226 11280
rect 20714 11268 20720 11280
rect 20220 11240 20720 11268
rect 20220 11228 20226 11240
rect 20714 11228 20720 11240
rect 20772 11228 20778 11280
rect 21450 11160 21456 11212
rect 21508 11200 21514 11212
rect 22465 11203 22523 11209
rect 22465 11200 22477 11203
rect 21508 11172 22477 11200
rect 21508 11160 21514 11172
rect 22465 11169 22477 11172
rect 22511 11169 22523 11203
rect 27908 11200 27936 11299
rect 29270 11296 29276 11348
rect 29328 11336 29334 11348
rect 29549 11339 29607 11345
rect 29549 11336 29561 11339
rect 29328 11308 29561 11336
rect 29328 11296 29334 11308
rect 29549 11305 29561 11308
rect 29595 11305 29607 11339
rect 29549 11299 29607 11305
rect 32217 11339 32275 11345
rect 32217 11305 32229 11339
rect 32263 11336 32275 11339
rect 32674 11336 32680 11348
rect 32263 11308 32680 11336
rect 32263 11305 32275 11308
rect 32217 11299 32275 11305
rect 32674 11296 32680 11308
rect 32732 11296 32738 11348
rect 33962 11296 33968 11348
rect 34020 11336 34026 11348
rect 34057 11339 34115 11345
rect 34057 11336 34069 11339
rect 34020 11308 34069 11336
rect 34020 11296 34026 11308
rect 34057 11305 34069 11308
rect 34103 11336 34115 11339
rect 34514 11336 34520 11348
rect 34103 11308 34520 11336
rect 34103 11305 34115 11308
rect 34057 11299 34115 11305
rect 34514 11296 34520 11308
rect 34572 11296 34578 11348
rect 38010 11336 38016 11348
rect 37971 11308 38016 11336
rect 38010 11296 38016 11308
rect 38068 11296 38074 11348
rect 28905 11271 28963 11277
rect 28905 11237 28917 11271
rect 28951 11268 28963 11271
rect 29454 11268 29460 11280
rect 28951 11240 29460 11268
rect 28951 11237 28963 11240
rect 28905 11231 28963 11237
rect 29454 11228 29460 11240
rect 29512 11228 29518 11280
rect 30650 11228 30656 11280
rect 30708 11268 30714 11280
rect 37001 11271 37059 11277
rect 37001 11268 37013 11271
rect 30708 11240 37013 11268
rect 30708 11228 30714 11240
rect 37001 11237 37013 11240
rect 37047 11237 37059 11271
rect 37001 11231 37059 11237
rect 30282 11200 30288 11212
rect 27908 11172 28672 11200
rect 22465 11163 22523 11169
rect 19884 11132 19942 11138
rect 19884 11126 19896 11132
rect 19812 11098 19896 11126
rect 19930 11098 19942 11132
rect 19884 11092 19942 11098
rect 19984 11135 20042 11141
rect 19984 11101 19996 11135
rect 20030 11101 20042 11135
rect 19984 11095 20042 11101
rect 20119 11135 20177 11141
rect 20119 11101 20131 11135
rect 20165 11132 20177 11135
rect 21358 11132 21364 11144
rect 20165 11104 21364 11132
rect 20165 11101 20208 11104
rect 20119 11095 20177 11101
rect 21358 11092 21364 11104
rect 21416 11092 21422 11144
rect 22480 11132 22508 11163
rect 23109 11135 23167 11141
rect 23109 11132 23121 11135
rect 22480 11104 23121 11132
rect 23109 11101 23121 11104
rect 23155 11101 23167 11135
rect 23109 11095 23167 11101
rect 23293 11135 23351 11141
rect 23293 11101 23305 11135
rect 23339 11132 23351 11135
rect 24762 11132 24768 11144
rect 23339 11104 24768 11132
rect 23339 11101 23351 11104
rect 23293 11095 23351 11101
rect 24762 11092 24768 11104
rect 24820 11132 24826 11144
rect 24903 11135 24961 11141
rect 24903 11132 24915 11135
rect 24820 11104 24915 11132
rect 24820 11092 24826 11104
rect 24903 11101 24915 11104
rect 24949 11101 24961 11135
rect 25038 11132 25044 11144
rect 24999 11104 25044 11132
rect 24903 11095 24961 11101
rect 25038 11092 25044 11104
rect 25096 11092 25102 11144
rect 25130 11092 25136 11144
rect 25188 11132 25194 11144
rect 25188 11104 25233 11132
rect 25188 11092 25194 11104
rect 25314 11092 25320 11144
rect 25372 11132 25378 11144
rect 26510 11132 26516 11144
rect 25372 11104 25417 11132
rect 26471 11104 26516 11132
rect 25372 11092 25378 11104
rect 26510 11092 26516 11104
rect 26568 11092 26574 11144
rect 26602 11092 26608 11144
rect 26660 11132 26666 11144
rect 26769 11135 26827 11141
rect 26769 11132 26781 11135
rect 26660 11104 26781 11132
rect 26660 11092 26666 11104
rect 26769 11101 26781 11104
rect 26815 11101 26827 11135
rect 26769 11095 26827 11101
rect 28353 11135 28411 11141
rect 28353 11101 28365 11135
rect 28399 11101 28411 11135
rect 28534 11132 28540 11144
rect 28495 11104 28540 11132
rect 28353 11095 28411 11101
rect 19242 11064 19248 11076
rect 18524 11036 19248 11064
rect 19242 11024 19248 11036
rect 19300 11024 19306 11076
rect 22370 11024 22376 11076
rect 22428 11064 22434 11076
rect 28368 11064 28396 11095
rect 28534 11092 28540 11104
rect 28592 11092 28598 11144
rect 28644 11141 28672 11172
rect 29840 11172 30288 11200
rect 28629 11135 28687 11141
rect 28629 11101 28641 11135
rect 28675 11101 28687 11135
rect 28629 11095 28687 11101
rect 28721 11135 28779 11141
rect 28721 11101 28733 11135
rect 28767 11101 28779 11135
rect 28721 11095 28779 11101
rect 22428 11036 28396 11064
rect 22428 11024 22434 11036
rect 28442 11024 28448 11076
rect 28500 11064 28506 11076
rect 28736 11064 28764 11095
rect 29362 11092 29368 11144
rect 29420 11132 29426 11144
rect 29840 11141 29868 11172
rect 30282 11160 30288 11172
rect 30340 11200 30346 11212
rect 30340 11172 32076 11200
rect 30340 11160 30346 11172
rect 29733 11135 29791 11141
rect 29733 11132 29745 11135
rect 29420 11104 29745 11132
rect 29420 11092 29426 11104
rect 29733 11101 29745 11104
rect 29779 11101 29791 11135
rect 29733 11095 29791 11101
rect 29825 11135 29883 11141
rect 29825 11101 29837 11135
rect 29871 11101 29883 11135
rect 29825 11095 29883 11101
rect 29914 11092 29920 11144
rect 29972 11132 29978 11144
rect 30101 11135 30159 11141
rect 29972 11104 30017 11132
rect 29972 11092 29978 11104
rect 30101 11101 30113 11135
rect 30147 11132 30159 11135
rect 30190 11132 30196 11144
rect 30147 11104 30196 11132
rect 30147 11101 30159 11104
rect 30101 11095 30159 11101
rect 30190 11092 30196 11104
rect 30248 11092 30254 11144
rect 31846 11132 31852 11144
rect 31807 11104 31852 11132
rect 31846 11092 31852 11104
rect 31904 11092 31910 11144
rect 32048 11141 32076 11172
rect 32214 11160 32220 11212
rect 32272 11200 32278 11212
rect 32490 11200 32496 11212
rect 32272 11172 32496 11200
rect 32272 11160 32278 11172
rect 32490 11160 32496 11172
rect 32548 11200 32554 11212
rect 32677 11203 32735 11209
rect 32677 11200 32689 11203
rect 32548 11172 32689 11200
rect 32548 11160 32554 11172
rect 32677 11169 32689 11172
rect 32723 11169 32735 11203
rect 32677 11163 32735 11169
rect 34514 11160 34520 11212
rect 34572 11200 34578 11212
rect 35069 11203 35127 11209
rect 35069 11200 35081 11203
rect 34572 11172 35081 11200
rect 34572 11160 34578 11172
rect 35069 11169 35081 11172
rect 35115 11169 35127 11203
rect 35069 11163 35127 11169
rect 32033 11135 32091 11141
rect 32033 11101 32045 11135
rect 32079 11101 32091 11135
rect 32033 11095 32091 11101
rect 34885 11135 34943 11141
rect 34885 11101 34897 11135
rect 34931 11101 34943 11135
rect 34885 11095 34943 11101
rect 28500 11036 28764 11064
rect 28500 11024 28506 11036
rect 32582 11024 32588 11076
rect 32640 11064 32646 11076
rect 33413 11067 33471 11073
rect 33413 11064 33425 11067
rect 32640 11036 33425 11064
rect 32640 11024 32646 11036
rect 33413 11033 33425 11036
rect 33459 11033 33471 11067
rect 33413 11027 33471 11033
rect 33597 11067 33655 11073
rect 33597 11033 33609 11067
rect 33643 11064 33655 11067
rect 34698 11064 34704 11076
rect 33643 11036 34704 11064
rect 33643 11033 33655 11036
rect 33597 11027 33655 11033
rect 34698 11024 34704 11036
rect 34756 11024 34762 11076
rect 34900 11064 34928 11095
rect 34974 11092 34980 11144
rect 35032 11132 35038 11144
rect 35529 11135 35587 11141
rect 35529 11132 35541 11135
rect 35032 11104 35541 11132
rect 35032 11092 35038 11104
rect 35529 11101 35541 11104
rect 35575 11101 35587 11135
rect 35529 11095 35587 11101
rect 35713 11135 35771 11141
rect 35713 11101 35725 11135
rect 35759 11132 35771 11135
rect 35802 11132 35808 11144
rect 35759 11104 35808 11132
rect 35759 11101 35771 11104
rect 35713 11095 35771 11101
rect 35342 11064 35348 11076
rect 34900 11036 35348 11064
rect 35342 11024 35348 11036
rect 35400 11024 35406 11076
rect 35544 11064 35572 11095
rect 35802 11092 35808 11104
rect 35860 11092 35866 11144
rect 37090 11092 37096 11144
rect 37148 11132 37154 11144
rect 37185 11135 37243 11141
rect 37185 11132 37197 11135
rect 37148 11104 37197 11132
rect 37148 11092 37154 11104
rect 37185 11101 37197 11104
rect 37231 11101 37243 11135
rect 37185 11095 37243 11101
rect 37274 11092 37280 11144
rect 37332 11132 37338 11144
rect 37553 11135 37611 11141
rect 37332 11104 37377 11132
rect 37332 11092 37338 11104
rect 37553 11101 37565 11135
rect 37599 11132 37611 11135
rect 38654 11132 38660 11144
rect 37599 11104 38660 11132
rect 37599 11101 37611 11104
rect 37553 11095 37611 11101
rect 38654 11092 38660 11104
rect 38712 11092 38718 11144
rect 36173 11067 36231 11073
rect 36173 11064 36185 11067
rect 35544 11036 36185 11064
rect 36173 11033 36185 11036
rect 36219 11033 36231 11067
rect 36173 11027 36231 11033
rect 37369 11067 37427 11073
rect 37369 11033 37381 11067
rect 37415 11033 37427 11067
rect 37369 11027 37427 11033
rect 13814 10996 13820 11008
rect 10428 10968 13820 10996
rect 10321 10959 10379 10965
rect 13814 10956 13820 10968
rect 13872 10956 13878 11008
rect 14274 10956 14280 11008
rect 14332 10996 14338 11008
rect 14369 10999 14427 11005
rect 14369 10996 14381 10999
rect 14332 10968 14381 10996
rect 14332 10956 14338 10968
rect 14369 10965 14381 10968
rect 14415 10965 14427 10999
rect 18230 10996 18236 11008
rect 18191 10968 18236 10996
rect 14369 10959 14427 10965
rect 18230 10956 18236 10968
rect 18288 10956 18294 11008
rect 20806 10996 20812 11008
rect 20767 10968 20812 10996
rect 20806 10956 20812 10968
rect 20864 10996 20870 11008
rect 21082 10996 21088 11008
rect 20864 10968 21088 10996
rect 20864 10956 20870 10968
rect 21082 10956 21088 10968
rect 21140 10956 21146 11008
rect 33229 10999 33287 11005
rect 33229 10965 33241 10999
rect 33275 10996 33287 10999
rect 33686 10996 33692 11008
rect 33275 10968 33692 10996
rect 33275 10965 33287 10968
rect 33229 10959 33287 10965
rect 33686 10956 33692 10968
rect 33744 10956 33750 11008
rect 35526 10996 35532 11008
rect 35487 10968 35532 10996
rect 35526 10956 35532 10968
rect 35584 10956 35590 11008
rect 37274 10956 37280 11008
rect 37332 10996 37338 11008
rect 37384 10996 37412 11027
rect 37332 10968 37412 10996
rect 37332 10956 37338 10968
rect 38378 10956 38384 11008
rect 38436 10996 38442 11008
rect 38565 10999 38623 11005
rect 38565 10996 38577 10999
rect 38436 10968 38577 10996
rect 38436 10956 38442 10968
rect 38565 10965 38577 10968
rect 38611 10965 38623 10999
rect 38565 10959 38623 10965
rect 1104 10906 68816 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 68816 10906
rect 1104 10832 68816 10854
rect 4522 10792 4528 10804
rect 4435 10764 4528 10792
rect 4522 10752 4528 10764
rect 4580 10792 4586 10804
rect 7742 10792 7748 10804
rect 4580 10764 7328 10792
rect 7703 10764 7748 10792
rect 4580 10752 4586 10764
rect 2222 10724 2228 10736
rect 2056 10696 2228 10724
rect 1762 10656 1768 10668
rect 1723 10628 1768 10656
rect 1762 10616 1768 10628
rect 1820 10616 1826 10668
rect 1854 10616 1860 10668
rect 1912 10656 1918 10668
rect 2056 10665 2084 10696
rect 2222 10684 2228 10696
rect 2280 10684 2286 10736
rect 2409 10727 2467 10733
rect 2409 10693 2421 10727
rect 2455 10724 2467 10727
rect 3390 10727 3448 10733
rect 3390 10724 3402 10727
rect 2455 10696 3402 10724
rect 2455 10693 2467 10696
rect 2409 10687 2467 10693
rect 3390 10693 3402 10696
rect 3436 10693 3448 10727
rect 3390 10687 3448 10693
rect 5810 10684 5816 10736
rect 5868 10724 5874 10736
rect 7300 10724 7328 10764
rect 7742 10752 7748 10764
rect 7800 10752 7806 10804
rect 10410 10792 10416 10804
rect 7852 10764 10272 10792
rect 7852 10724 7880 10764
rect 5868 10696 7236 10724
rect 7300 10696 7880 10724
rect 7929 10727 7987 10733
rect 5868 10684 5874 10696
rect 1949 10659 2007 10665
rect 1949 10656 1961 10659
rect 1912 10628 1961 10656
rect 1912 10616 1918 10628
rect 1949 10625 1961 10628
rect 1995 10625 2007 10659
rect 1949 10619 2007 10625
rect 2041 10659 2099 10665
rect 2041 10625 2053 10659
rect 2087 10625 2099 10659
rect 2041 10619 2099 10625
rect 2130 10616 2136 10668
rect 2188 10656 2194 10668
rect 3142 10656 3148 10668
rect 2188 10628 2233 10656
rect 3103 10628 3148 10656
rect 2188 10616 2194 10628
rect 3142 10616 3148 10628
rect 3200 10616 3206 10668
rect 3234 10616 3240 10668
rect 3292 10656 3298 10668
rect 6641 10659 6699 10665
rect 3292 10628 5856 10656
rect 3292 10616 3298 10628
rect 5828 10597 5856 10628
rect 6641 10625 6653 10659
rect 6687 10625 6699 10659
rect 6641 10619 6699 10625
rect 6733 10659 6791 10665
rect 6733 10625 6745 10659
rect 6779 10625 6791 10659
rect 6733 10619 6791 10625
rect 5813 10591 5871 10597
rect 5813 10557 5825 10591
rect 5859 10588 5871 10591
rect 6656 10588 6684 10619
rect 5859 10560 6684 10588
rect 6748 10588 6776 10619
rect 6822 10616 6828 10668
rect 6880 10656 6886 10668
rect 6880 10628 6925 10656
rect 6880 10616 6886 10628
rect 7006 10616 7012 10668
rect 7064 10656 7070 10668
rect 7208 10656 7236 10696
rect 7929 10693 7941 10727
rect 7975 10724 7987 10727
rect 7975 10696 9674 10724
rect 7975 10693 7987 10696
rect 7929 10687 7987 10693
rect 8113 10659 8171 10665
rect 8113 10656 8125 10659
rect 7064 10628 7109 10656
rect 7208 10628 8125 10656
rect 7064 10616 7070 10628
rect 8113 10625 8125 10628
rect 8159 10625 8171 10659
rect 8113 10619 8171 10625
rect 8573 10659 8631 10665
rect 8573 10625 8585 10659
rect 8619 10656 8631 10659
rect 8754 10656 8760 10668
rect 8619 10628 8760 10656
rect 8619 10625 8631 10628
rect 8573 10619 8631 10625
rect 8754 10616 8760 10628
rect 8812 10616 8818 10668
rect 9646 10656 9674 10696
rect 10134 10656 10140 10668
rect 9646 10628 10140 10656
rect 10134 10616 10140 10628
rect 10192 10616 10198 10668
rect 10244 10656 10272 10764
rect 10336 10764 10416 10792
rect 10336 10733 10364 10764
rect 10410 10752 10416 10764
rect 10468 10752 10474 10804
rect 12158 10752 12164 10804
rect 12216 10792 12222 10804
rect 14461 10795 14519 10801
rect 12216 10764 13768 10792
rect 12216 10752 12222 10764
rect 10321 10727 10379 10733
rect 10321 10693 10333 10727
rect 10367 10693 10379 10727
rect 10321 10687 10379 10693
rect 12526 10684 12532 10736
rect 12584 10724 12590 10736
rect 13740 10724 13768 10764
rect 14461 10761 14473 10795
rect 14507 10792 14519 10795
rect 15194 10792 15200 10804
rect 14507 10764 15200 10792
rect 14507 10761 14519 10764
rect 14461 10755 14519 10761
rect 15194 10752 15200 10764
rect 15252 10752 15258 10804
rect 18049 10795 18107 10801
rect 18049 10761 18061 10795
rect 18095 10792 18107 10795
rect 18414 10792 18420 10804
rect 18095 10764 18420 10792
rect 18095 10761 18107 10764
rect 18049 10755 18107 10761
rect 18414 10752 18420 10764
rect 18472 10752 18478 10804
rect 19242 10752 19248 10804
rect 19300 10792 19306 10804
rect 22281 10795 22339 10801
rect 19300 10764 22094 10792
rect 19300 10752 19306 10764
rect 16390 10724 16396 10736
rect 12584 10696 12940 10724
rect 12584 10684 12590 10696
rect 10413 10659 10471 10665
rect 10413 10656 10425 10659
rect 10244 10628 10425 10656
rect 10413 10625 10425 10628
rect 10459 10625 10471 10659
rect 10413 10619 10471 10625
rect 10505 10659 10563 10665
rect 10505 10625 10517 10659
rect 10551 10656 10563 10659
rect 10594 10656 10600 10668
rect 10551 10628 10600 10656
rect 10551 10625 10563 10628
rect 10505 10619 10563 10625
rect 10594 10616 10600 10628
rect 10652 10616 10658 10668
rect 11422 10616 11428 10668
rect 11480 10656 11486 10668
rect 12912 10665 12940 10696
rect 13740 10696 16396 10724
rect 13740 10665 13768 10696
rect 16390 10684 16396 10696
rect 16448 10684 16454 10736
rect 17126 10684 17132 10736
rect 17184 10724 17190 10736
rect 18509 10727 18567 10733
rect 18509 10724 18521 10727
rect 17184 10696 18521 10724
rect 17184 10684 17190 10696
rect 18509 10693 18521 10696
rect 18555 10693 18567 10727
rect 18509 10687 18567 10693
rect 19794 10684 19800 10736
rect 19852 10724 19858 10736
rect 22066 10724 22094 10764
rect 22281 10761 22293 10795
rect 22327 10792 22339 10795
rect 23934 10792 23940 10804
rect 22327 10764 23940 10792
rect 22327 10761 22339 10764
rect 22281 10755 22339 10761
rect 23934 10752 23940 10764
rect 23992 10752 23998 10804
rect 24762 10792 24768 10804
rect 24723 10764 24768 10792
rect 24762 10752 24768 10764
rect 24820 10752 24826 10804
rect 25498 10752 25504 10804
rect 25556 10792 25562 10804
rect 25685 10795 25743 10801
rect 25685 10792 25697 10795
rect 25556 10764 25697 10792
rect 25556 10752 25562 10764
rect 25685 10761 25697 10764
rect 25731 10761 25743 10795
rect 26234 10792 26240 10804
rect 26195 10764 26240 10792
rect 25685 10755 25743 10761
rect 26234 10752 26240 10764
rect 26292 10792 26298 10804
rect 26602 10792 26608 10804
rect 26292 10764 26608 10792
rect 26292 10752 26298 10764
rect 26602 10752 26608 10764
rect 26660 10752 26666 10804
rect 29825 10795 29883 10801
rect 29825 10761 29837 10795
rect 29871 10761 29883 10795
rect 32674 10792 32680 10804
rect 32635 10764 32680 10792
rect 29825 10755 29883 10761
rect 29840 10724 29868 10755
rect 32674 10752 32680 10764
rect 32732 10752 32738 10804
rect 34514 10792 34520 10804
rect 34475 10764 34520 10792
rect 34514 10752 34520 10764
rect 34572 10792 34578 10804
rect 34572 10764 35112 10792
rect 34572 10752 34578 10764
rect 19852 10696 21956 10724
rect 22066 10696 29868 10724
rect 19852 10684 19858 10696
rect 12630 10659 12688 10665
rect 12630 10656 12642 10659
rect 11480 10628 12642 10656
rect 11480 10616 11486 10628
rect 12630 10625 12642 10628
rect 12676 10625 12688 10659
rect 12630 10619 12688 10625
rect 12897 10659 12955 10665
rect 12897 10625 12909 10659
rect 12943 10625 12955 10659
rect 12897 10619 12955 10625
rect 13725 10659 13783 10665
rect 13725 10625 13737 10659
rect 13771 10625 13783 10659
rect 13906 10656 13912 10668
rect 13867 10628 13912 10656
rect 13725 10619 13783 10625
rect 13906 10616 13912 10628
rect 13964 10616 13970 10668
rect 14274 10656 14280 10668
rect 14235 10628 14280 10656
rect 14274 10616 14280 10628
rect 14332 10616 14338 10668
rect 15933 10659 15991 10665
rect 15933 10625 15945 10659
rect 15979 10656 15991 10659
rect 16298 10656 16304 10668
rect 15979 10628 16304 10656
rect 15979 10625 15991 10628
rect 15933 10619 15991 10625
rect 7926 10588 7932 10600
rect 6748 10560 7932 10588
rect 5859 10557 5871 10560
rect 5813 10551 5871 10557
rect 6656 10520 6684 10560
rect 7926 10548 7932 10560
rect 7984 10548 7990 10600
rect 13998 10588 14004 10600
rect 8036 10560 11652 10588
rect 13959 10560 14004 10588
rect 8036 10520 8064 10560
rect 10686 10520 10692 10532
rect 6656 10492 8064 10520
rect 10647 10492 10692 10520
rect 10686 10480 10692 10492
rect 10744 10480 10750 10532
rect 2038 10412 2044 10464
rect 2096 10452 2102 10464
rect 4522 10452 4528 10464
rect 2096 10424 4528 10452
rect 2096 10412 2102 10424
rect 4522 10412 4528 10424
rect 4580 10412 4586 10464
rect 6362 10452 6368 10464
rect 6323 10424 6368 10452
rect 6362 10412 6368 10424
rect 6420 10412 6426 10464
rect 11514 10452 11520 10464
rect 11475 10424 11520 10452
rect 11514 10412 11520 10424
rect 11572 10412 11578 10464
rect 11624 10452 11652 10560
rect 13998 10548 14004 10560
rect 14056 10548 14062 10600
rect 14090 10548 14096 10600
rect 14148 10588 14154 10600
rect 14148 10560 14193 10588
rect 14148 10548 14154 10560
rect 13262 10480 13268 10532
rect 13320 10520 13326 10532
rect 15948 10520 15976 10619
rect 16298 10616 16304 10628
rect 16356 10656 16362 10668
rect 17037 10659 17095 10665
rect 17037 10656 17049 10659
rect 16356 10628 17049 10656
rect 16356 10616 16362 10628
rect 17037 10625 17049 10628
rect 17083 10625 17095 10659
rect 17037 10619 17095 10625
rect 19978 10616 19984 10668
rect 20036 10656 20042 10668
rect 20073 10659 20131 10665
rect 20073 10656 20085 10659
rect 20036 10628 20085 10656
rect 20036 10616 20042 10628
rect 20073 10625 20085 10628
rect 20119 10625 20131 10659
rect 20073 10619 20131 10625
rect 20901 10659 20959 10665
rect 20901 10625 20913 10659
rect 20947 10656 20959 10659
rect 21542 10656 21548 10668
rect 20947 10628 21548 10656
rect 20947 10625 20959 10628
rect 20901 10619 20959 10625
rect 21542 10616 21548 10628
rect 21600 10616 21606 10668
rect 16117 10591 16175 10597
rect 16117 10557 16129 10591
rect 16163 10588 16175 10591
rect 20806 10588 20812 10600
rect 16163 10560 20812 10588
rect 16163 10557 16175 10560
rect 16117 10551 16175 10557
rect 20806 10548 20812 10560
rect 20864 10588 20870 10600
rect 21085 10591 21143 10597
rect 21085 10588 21097 10591
rect 20864 10560 21097 10588
rect 20864 10548 20870 10560
rect 21085 10557 21097 10560
rect 21131 10557 21143 10591
rect 21928 10588 21956 10696
rect 30742 10684 30748 10736
rect 30800 10724 30806 10736
rect 34974 10724 34980 10736
rect 30800 10696 34980 10724
rect 30800 10684 30806 10696
rect 34532 10668 34560 10696
rect 34974 10684 34980 10696
rect 35032 10684 35038 10736
rect 22186 10656 22192 10668
rect 22147 10628 22192 10656
rect 22186 10616 22192 10628
rect 22244 10616 22250 10668
rect 23014 10656 23020 10668
rect 22927 10628 23020 10656
rect 23014 10616 23020 10628
rect 23072 10656 23078 10668
rect 24029 10659 24087 10665
rect 24029 10656 24041 10659
rect 23072 10628 24041 10656
rect 23072 10616 23078 10628
rect 24029 10625 24041 10628
rect 24075 10625 24087 10659
rect 24029 10619 24087 10625
rect 22830 10588 22836 10600
rect 21928 10560 22836 10588
rect 21085 10551 21143 10557
rect 22830 10548 22836 10560
rect 22888 10548 22894 10600
rect 13320 10492 15976 10520
rect 17221 10523 17279 10529
rect 13320 10480 13326 10492
rect 17221 10489 17233 10523
rect 17267 10520 17279 10523
rect 20530 10520 20536 10532
rect 17267 10492 20536 10520
rect 17267 10489 17279 10492
rect 17221 10483 17279 10489
rect 20530 10480 20536 10492
rect 20588 10480 20594 10532
rect 13446 10452 13452 10464
rect 11624 10424 13452 10452
rect 13446 10412 13452 10424
rect 13504 10412 13510 10464
rect 20717 10455 20775 10461
rect 20717 10421 20729 10455
rect 20763 10452 20775 10455
rect 21082 10452 21088 10464
rect 20763 10424 21088 10452
rect 20763 10421 20775 10424
rect 20717 10415 20775 10421
rect 21082 10412 21088 10424
rect 21140 10412 21146 10464
rect 23201 10455 23259 10461
rect 23201 10421 23213 10455
rect 23247 10452 23259 10455
rect 23566 10452 23572 10464
rect 23247 10424 23572 10452
rect 23247 10421 23259 10424
rect 23201 10415 23259 10421
rect 23566 10412 23572 10424
rect 23624 10412 23630 10464
rect 24044 10452 24072 10619
rect 24118 10616 24124 10668
rect 24176 10656 24182 10668
rect 24213 10659 24271 10665
rect 24213 10656 24225 10659
rect 24176 10628 24225 10656
rect 24176 10616 24182 10628
rect 24213 10625 24225 10628
rect 24259 10625 24271 10659
rect 24213 10619 24271 10625
rect 25317 10659 25375 10665
rect 25317 10625 25329 10659
rect 25363 10656 25375 10659
rect 25406 10656 25412 10668
rect 25363 10628 25412 10656
rect 25363 10625 25375 10628
rect 25317 10619 25375 10625
rect 25406 10616 25412 10628
rect 25464 10616 25470 10668
rect 25501 10659 25559 10665
rect 25501 10625 25513 10659
rect 25547 10656 25559 10659
rect 26142 10656 26148 10668
rect 25547 10628 26148 10656
rect 25547 10625 25559 10628
rect 25501 10619 25559 10625
rect 26142 10616 26148 10628
rect 26200 10616 26206 10668
rect 28810 10656 28816 10668
rect 28771 10628 28816 10656
rect 28810 10616 28816 10628
rect 28868 10656 28874 10668
rect 29365 10659 29423 10665
rect 29365 10656 29377 10659
rect 28868 10628 29377 10656
rect 28868 10616 28874 10628
rect 29365 10625 29377 10628
rect 29411 10625 29423 10659
rect 29365 10619 29423 10625
rect 29641 10659 29699 10665
rect 29641 10625 29653 10659
rect 29687 10656 29699 10659
rect 30650 10656 30656 10668
rect 29687 10628 30656 10656
rect 29687 10625 29699 10628
rect 29641 10619 29699 10625
rect 30650 10616 30656 10628
rect 30708 10616 30714 10668
rect 32674 10616 32680 10668
rect 32732 10656 32738 10668
rect 33505 10659 33563 10665
rect 33505 10656 33517 10659
rect 32732 10628 33517 10656
rect 32732 10616 32738 10628
rect 33505 10625 33517 10628
rect 33551 10625 33563 10659
rect 33505 10619 33563 10625
rect 33597 10659 33655 10665
rect 33597 10625 33609 10659
rect 33643 10625 33655 10659
rect 33597 10619 33655 10625
rect 29454 10588 29460 10600
rect 29415 10560 29460 10588
rect 29454 10548 29460 10560
rect 29512 10548 29518 10600
rect 33612 10588 33640 10619
rect 33686 10616 33692 10668
rect 33744 10656 33750 10668
rect 33744 10628 33789 10656
rect 33744 10616 33750 10628
rect 33870 10616 33876 10668
rect 33928 10656 33934 10668
rect 33928 10628 33973 10656
rect 33928 10616 33934 10628
rect 34514 10616 34520 10668
rect 34572 10616 34578 10668
rect 35084 10665 35112 10764
rect 35434 10724 35440 10736
rect 35347 10696 35440 10724
rect 35434 10684 35440 10696
rect 35492 10724 35498 10736
rect 38657 10727 38715 10733
rect 35492 10696 37320 10724
rect 35492 10684 35498 10696
rect 35069 10659 35127 10665
rect 35069 10625 35081 10659
rect 35115 10625 35127 10659
rect 35069 10619 35127 10625
rect 35253 10659 35311 10665
rect 35253 10625 35265 10659
rect 35299 10656 35311 10659
rect 35802 10656 35808 10668
rect 35299 10628 35808 10656
rect 35299 10625 35311 10628
rect 35253 10619 35311 10625
rect 35802 10616 35808 10628
rect 35860 10616 35866 10668
rect 37292 10665 37320 10696
rect 38657 10693 38669 10727
rect 38703 10724 38715 10727
rect 40230 10727 40288 10733
rect 40230 10724 40242 10727
rect 38703 10696 40242 10724
rect 38703 10693 38715 10696
rect 38657 10687 38715 10693
rect 40230 10693 40242 10696
rect 40276 10693 40288 10727
rect 40230 10687 40288 10693
rect 37277 10659 37335 10665
rect 37277 10625 37289 10659
rect 37323 10625 37335 10659
rect 37277 10619 37335 10625
rect 37458 10616 37464 10668
rect 37516 10656 37522 10668
rect 38010 10656 38016 10668
rect 37516 10628 38016 10656
rect 37516 10616 37522 10628
rect 38010 10616 38016 10628
rect 38068 10616 38074 10668
rect 38194 10656 38200 10668
rect 38155 10628 38200 10656
rect 38194 10616 38200 10628
rect 38252 10616 38258 10668
rect 38289 10659 38347 10665
rect 38289 10625 38301 10659
rect 38335 10625 38347 10659
rect 38289 10619 38347 10625
rect 34790 10588 34796 10600
rect 33612 10560 34796 10588
rect 34790 10548 34796 10560
rect 34848 10548 34854 10600
rect 35526 10548 35532 10600
rect 35584 10588 35590 10600
rect 35897 10591 35955 10597
rect 35897 10588 35909 10591
rect 35584 10560 35909 10588
rect 35584 10548 35590 10560
rect 35897 10557 35909 10560
rect 35943 10557 35955 10591
rect 35897 10551 35955 10557
rect 36173 10591 36231 10597
rect 36173 10557 36185 10591
rect 36219 10588 36231 10591
rect 37918 10588 37924 10600
rect 36219 10560 37924 10588
rect 36219 10557 36231 10560
rect 36173 10551 36231 10557
rect 37918 10548 37924 10560
rect 37976 10588 37982 10600
rect 38304 10588 38332 10619
rect 38378 10616 38384 10668
rect 38436 10656 38442 10668
rect 40494 10656 40500 10668
rect 38436 10628 38481 10656
rect 40455 10628 40500 10656
rect 38436 10616 38442 10628
rect 40494 10616 40500 10628
rect 40552 10616 40558 10668
rect 37976 10560 38332 10588
rect 37976 10548 37982 10560
rect 24121 10523 24179 10529
rect 24121 10489 24133 10523
rect 24167 10520 24179 10523
rect 24854 10520 24860 10532
rect 24167 10492 24860 10520
rect 24167 10489 24179 10492
rect 24121 10483 24179 10489
rect 24854 10480 24860 10492
rect 24912 10480 24918 10532
rect 28718 10480 28724 10532
rect 28776 10520 28782 10532
rect 36814 10520 36820 10532
rect 28776 10492 36820 10520
rect 28776 10480 28782 10492
rect 36814 10480 36820 10492
rect 36872 10480 36878 10532
rect 26142 10452 26148 10464
rect 24044 10424 26148 10452
rect 26142 10412 26148 10424
rect 26200 10412 26206 10464
rect 29546 10452 29552 10464
rect 29507 10424 29552 10452
rect 29546 10412 29552 10424
rect 29604 10412 29610 10464
rect 33226 10452 33232 10464
rect 33187 10424 33232 10452
rect 33226 10412 33232 10424
rect 33284 10412 33290 10464
rect 37366 10412 37372 10464
rect 37424 10452 37430 10464
rect 37461 10455 37519 10461
rect 37461 10452 37473 10455
rect 37424 10424 37473 10452
rect 37424 10412 37430 10424
rect 37461 10421 37473 10424
rect 37507 10452 37519 10455
rect 37918 10452 37924 10464
rect 37507 10424 37924 10452
rect 37507 10421 37519 10424
rect 37461 10415 37519 10421
rect 37918 10412 37924 10424
rect 37976 10412 37982 10464
rect 38102 10412 38108 10464
rect 38160 10452 38166 10464
rect 39117 10455 39175 10461
rect 39117 10452 39129 10455
rect 38160 10424 39129 10452
rect 38160 10412 38166 10424
rect 39117 10421 39129 10424
rect 39163 10421 39175 10455
rect 67634 10452 67640 10464
rect 67595 10424 67640 10452
rect 39117 10415 39175 10421
rect 67634 10412 67640 10424
rect 67692 10412 67698 10464
rect 1104 10362 68816 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 65654 10362
rect 65706 10310 65718 10362
rect 65770 10310 65782 10362
rect 65834 10310 65846 10362
rect 65898 10310 65910 10362
rect 65962 10310 68816 10362
rect 1104 10288 68816 10310
rect 1854 10248 1860 10260
rect 1815 10220 1860 10248
rect 1854 10208 1860 10220
rect 1912 10208 1918 10260
rect 6549 10251 6607 10257
rect 6549 10217 6561 10251
rect 6595 10248 6607 10251
rect 6822 10248 6828 10260
rect 6595 10220 6828 10248
rect 6595 10217 6607 10220
rect 6549 10211 6607 10217
rect 6822 10208 6828 10220
rect 6880 10208 6886 10260
rect 9033 10251 9091 10257
rect 9033 10217 9045 10251
rect 9079 10248 9091 10251
rect 10962 10248 10968 10260
rect 9079 10220 10968 10248
rect 9079 10217 9091 10220
rect 9033 10211 9091 10217
rect 2130 10140 2136 10192
rect 2188 10180 2194 10192
rect 2777 10183 2835 10189
rect 2777 10180 2789 10183
rect 2188 10152 2789 10180
rect 2188 10140 2194 10152
rect 2777 10149 2789 10152
rect 2823 10180 2835 10183
rect 8754 10180 8760 10192
rect 2823 10152 8760 10180
rect 2823 10149 2835 10152
rect 2777 10143 2835 10149
rect 8754 10140 8760 10152
rect 8812 10140 8818 10192
rect 7926 10112 7932 10124
rect 7760 10084 7932 10112
rect 2038 10044 2044 10056
rect 1999 10016 2044 10044
rect 2038 10004 2044 10016
rect 2096 10004 2102 10056
rect 2225 10047 2283 10053
rect 2225 10013 2237 10047
rect 2271 10044 2283 10047
rect 2406 10044 2412 10056
rect 2271 10016 2412 10044
rect 2271 10013 2283 10016
rect 2225 10007 2283 10013
rect 2406 10004 2412 10016
rect 2464 10044 2470 10056
rect 3786 10044 3792 10056
rect 2464 10016 3792 10044
rect 2464 10004 2470 10016
rect 3786 10004 3792 10016
rect 3844 10004 3850 10056
rect 5810 10004 5816 10056
rect 5868 10044 5874 10056
rect 6181 10047 6239 10053
rect 6181 10044 6193 10047
rect 5868 10016 6193 10044
rect 5868 10004 5874 10016
rect 6181 10013 6193 10016
rect 6227 10013 6239 10047
rect 6181 10007 6239 10013
rect 7006 10004 7012 10056
rect 7064 10044 7070 10056
rect 7469 10047 7527 10053
rect 7469 10044 7481 10047
rect 7064 10016 7481 10044
rect 7064 10004 7070 10016
rect 7469 10013 7481 10016
rect 7515 10013 7527 10047
rect 7650 10044 7656 10056
rect 7611 10016 7656 10044
rect 7469 10007 7527 10013
rect 7650 10004 7656 10016
rect 7708 10004 7714 10056
rect 7760 10053 7788 10084
rect 7926 10072 7932 10084
rect 7984 10072 7990 10124
rect 7745 10047 7803 10053
rect 7745 10013 7757 10047
rect 7791 10013 7803 10047
rect 7745 10007 7803 10013
rect 7834 10004 7840 10056
rect 7892 10044 7898 10056
rect 9048 10044 9076 10211
rect 10962 10208 10968 10220
rect 11020 10208 11026 10260
rect 11422 10248 11428 10260
rect 11383 10220 11428 10248
rect 11422 10208 11428 10220
rect 11480 10208 11486 10260
rect 13998 10248 14004 10260
rect 12406 10220 14004 10248
rect 9674 10140 9680 10192
rect 9732 10180 9738 10192
rect 12406 10180 12434 10220
rect 13998 10208 14004 10220
rect 14056 10208 14062 10260
rect 17494 10248 17500 10260
rect 17455 10220 17500 10248
rect 17494 10208 17500 10220
rect 17552 10208 17558 10260
rect 18046 10248 18052 10260
rect 18007 10220 18052 10248
rect 18046 10208 18052 10220
rect 18104 10208 18110 10260
rect 19337 10251 19395 10257
rect 19337 10217 19349 10251
rect 19383 10248 19395 10251
rect 20162 10248 20168 10260
rect 19383 10220 20168 10248
rect 19383 10217 19395 10220
rect 19337 10211 19395 10217
rect 20162 10208 20168 10220
rect 20220 10208 20226 10260
rect 20622 10208 20628 10260
rect 20680 10248 20686 10260
rect 22830 10248 22836 10260
rect 20680 10220 22094 10248
rect 22791 10220 22836 10248
rect 20680 10208 20686 10220
rect 9732 10152 12434 10180
rect 9732 10140 9738 10152
rect 12618 10140 12624 10192
rect 12676 10180 12682 10192
rect 17221 10183 17279 10189
rect 17221 10180 17233 10183
rect 12676 10152 17233 10180
rect 12676 10140 12682 10152
rect 17221 10149 17233 10152
rect 17267 10149 17279 10183
rect 18230 10180 18236 10192
rect 17221 10143 17279 10149
rect 17328 10152 18236 10180
rect 10134 10112 10140 10124
rect 9876 10084 10140 10112
rect 7892 10016 9076 10044
rect 7892 10004 7898 10016
rect 9398 10004 9404 10056
rect 9456 10044 9462 10056
rect 9876 10053 9904 10084
rect 10134 10072 10140 10084
rect 10192 10112 10198 10124
rect 10410 10112 10416 10124
rect 10192 10084 10416 10112
rect 10192 10072 10198 10084
rect 10410 10072 10416 10084
rect 10468 10072 10474 10124
rect 10686 10072 10692 10124
rect 10744 10112 10750 10124
rect 11885 10115 11943 10121
rect 11885 10112 11897 10115
rect 10744 10084 11897 10112
rect 10744 10072 10750 10084
rect 11885 10081 11897 10084
rect 11931 10081 11943 10115
rect 17328 10112 17356 10152
rect 18230 10140 18236 10152
rect 18288 10140 18294 10192
rect 19518 10140 19524 10192
rect 19576 10180 19582 10192
rect 22066 10180 22094 10220
rect 22830 10208 22836 10220
rect 22888 10208 22894 10260
rect 23845 10251 23903 10257
rect 23845 10217 23857 10251
rect 23891 10248 23903 10251
rect 24302 10248 24308 10260
rect 23891 10220 24308 10248
rect 23891 10217 23903 10220
rect 23845 10211 23903 10217
rect 24302 10208 24308 10220
rect 24360 10248 24366 10260
rect 25406 10248 25412 10260
rect 24360 10220 25412 10248
rect 24360 10208 24366 10220
rect 25406 10208 25412 10220
rect 25464 10208 25470 10260
rect 27801 10251 27859 10257
rect 27801 10217 27813 10251
rect 27847 10248 27859 10251
rect 28074 10248 28080 10260
rect 27847 10220 28080 10248
rect 27847 10217 27859 10220
rect 27801 10211 27859 10217
rect 28074 10208 28080 10220
rect 28132 10208 28138 10260
rect 28905 10251 28963 10257
rect 28905 10217 28917 10251
rect 28951 10248 28963 10251
rect 29178 10248 29184 10260
rect 28951 10220 29184 10248
rect 28951 10217 28963 10220
rect 28905 10211 28963 10217
rect 29178 10208 29184 10220
rect 29236 10208 29242 10260
rect 31386 10208 31392 10260
rect 31444 10248 31450 10260
rect 32582 10248 32588 10260
rect 31444 10220 32588 10248
rect 31444 10208 31450 10220
rect 32582 10208 32588 10220
rect 32640 10208 32646 10260
rect 34790 10248 34796 10260
rect 34751 10220 34796 10248
rect 34790 10208 34796 10220
rect 34848 10208 34854 10260
rect 36906 10248 36912 10260
rect 36867 10220 36912 10248
rect 36906 10208 36912 10220
rect 36964 10208 36970 10260
rect 38194 10208 38200 10260
rect 38252 10248 38258 10260
rect 38289 10251 38347 10257
rect 38289 10248 38301 10251
rect 38252 10220 38301 10248
rect 38252 10208 38258 10220
rect 38289 10217 38301 10220
rect 38335 10217 38347 10251
rect 38289 10211 38347 10217
rect 22373 10183 22431 10189
rect 22373 10180 22385 10183
rect 19576 10152 19932 10180
rect 22066 10152 22385 10180
rect 19576 10140 19582 10152
rect 11885 10075 11943 10081
rect 11992 10084 17356 10112
rect 17497 10115 17555 10121
rect 9677 10047 9735 10053
rect 9677 10044 9689 10047
rect 9456 10016 9689 10044
rect 9456 10004 9462 10016
rect 9677 10013 9689 10016
rect 9723 10013 9735 10047
rect 9677 10007 9735 10013
rect 9861 10047 9919 10053
rect 9861 10013 9873 10047
rect 9907 10013 9919 10047
rect 9861 10007 9919 10013
rect 10045 10047 10103 10053
rect 10045 10013 10057 10047
rect 10091 10044 10103 10047
rect 10594 10044 10600 10056
rect 10091 10016 10600 10044
rect 10091 10013 10103 10016
rect 10045 10007 10103 10013
rect 10594 10004 10600 10016
rect 10652 10004 10658 10056
rect 11606 10044 11612 10056
rect 11567 10016 11612 10044
rect 11606 10004 11612 10016
rect 11664 10004 11670 10056
rect 11992 10053 12020 10084
rect 17497 10081 17509 10115
rect 17543 10112 17555 10115
rect 19702 10112 19708 10124
rect 17543 10084 19708 10112
rect 17543 10081 17555 10084
rect 17497 10075 17555 10081
rect 19702 10072 19708 10084
rect 19760 10072 19766 10124
rect 19904 10112 19932 10152
rect 22373 10149 22385 10152
rect 22419 10180 22431 10183
rect 28534 10180 28540 10192
rect 22419 10152 27292 10180
rect 28495 10152 28540 10180
rect 22419 10149 22431 10152
rect 22373 10143 22431 10149
rect 19904 10084 20024 10112
rect 11793 10047 11851 10053
rect 11793 10013 11805 10047
rect 11839 10013 11851 10047
rect 11793 10007 11851 10013
rect 11977 10047 12035 10053
rect 11977 10013 11989 10047
rect 12023 10013 12035 10047
rect 12158 10044 12164 10056
rect 12119 10016 12164 10044
rect 11977 10007 12035 10013
rect 3970 9976 3976 9988
rect 3883 9948 3976 9976
rect 3970 9936 3976 9948
rect 4028 9976 4034 9988
rect 6365 9979 6423 9985
rect 4028 9948 6040 9976
rect 4028 9936 4034 9948
rect 4154 9908 4160 9920
rect 4115 9880 4160 9908
rect 4154 9868 4160 9880
rect 4212 9868 4218 9920
rect 4709 9911 4767 9917
rect 4709 9877 4721 9911
rect 4755 9908 4767 9911
rect 5442 9908 5448 9920
rect 4755 9880 5448 9908
rect 4755 9877 4767 9880
rect 4709 9871 4767 9877
rect 5442 9868 5448 9880
rect 5500 9868 5506 9920
rect 6012 9908 6040 9948
rect 6365 9945 6377 9979
rect 6411 9976 6423 9979
rect 6914 9976 6920 9988
rect 6411 9948 6920 9976
rect 6411 9945 6423 9948
rect 6365 9939 6423 9945
rect 6914 9936 6920 9948
rect 6972 9936 6978 9988
rect 9953 9979 10011 9985
rect 9953 9976 9965 9979
rect 7024 9948 9965 9976
rect 7024 9908 7052 9948
rect 9953 9945 9965 9948
rect 9999 9945 10011 9979
rect 11808 9976 11836 10007
rect 12158 10004 12164 10016
rect 12216 10004 12222 10056
rect 14090 10044 14096 10056
rect 12406 10016 14096 10044
rect 12406 9976 12434 10016
rect 14090 10004 14096 10016
rect 14148 10004 14154 10056
rect 14185 10047 14243 10053
rect 14185 10013 14197 10047
rect 14231 10044 14243 10047
rect 15838 10044 15844 10056
rect 14231 10016 15844 10044
rect 14231 10013 14243 10016
rect 14185 10007 14243 10013
rect 15838 10004 15844 10016
rect 15896 10004 15902 10056
rect 16298 10044 16304 10056
rect 16259 10016 16304 10044
rect 16298 10004 16304 10016
rect 16356 10004 16362 10056
rect 17586 10004 17592 10056
rect 17644 10044 17650 10056
rect 18322 10044 18328 10056
rect 17644 10016 17689 10044
rect 18283 10016 18328 10044
rect 17644 10004 17650 10016
rect 18322 10004 18328 10016
rect 18380 10004 18386 10056
rect 18417 10047 18475 10053
rect 18417 10013 18429 10047
rect 18463 10013 18475 10047
rect 18417 10007 18475 10013
rect 11808 9948 12434 9976
rect 9953 9939 10011 9945
rect 11992 9920 12020 9948
rect 13814 9936 13820 9988
rect 13872 9976 13878 9988
rect 18432 9976 18460 10007
rect 18506 10004 18512 10056
rect 18564 10044 18570 10056
rect 18693 10047 18751 10053
rect 18564 10016 18609 10044
rect 18564 10004 18570 10016
rect 18693 10013 18705 10047
rect 18739 10044 18751 10047
rect 19426 10044 19432 10056
rect 18739 10016 19432 10044
rect 18739 10013 18751 10016
rect 18693 10007 18751 10013
rect 19426 10004 19432 10016
rect 19484 10044 19490 10056
rect 19996 10053 20024 10084
rect 20806 10072 20812 10124
rect 20864 10112 20870 10124
rect 20993 10115 21051 10121
rect 20993 10112 21005 10115
rect 20864 10084 21005 10112
rect 20864 10072 20870 10084
rect 20993 10081 21005 10084
rect 21039 10081 21051 10115
rect 24854 10112 24860 10124
rect 24815 10084 24860 10112
rect 20993 10075 21051 10081
rect 24854 10072 24860 10084
rect 24912 10072 24918 10124
rect 25038 10072 25044 10124
rect 25096 10112 25102 10124
rect 25133 10115 25191 10121
rect 25133 10112 25145 10115
rect 25096 10084 25145 10112
rect 25096 10072 25102 10084
rect 25133 10081 25145 10084
rect 25179 10112 25191 10115
rect 25179 10084 26464 10112
rect 25179 10081 25191 10084
rect 25133 10075 25191 10081
rect 19797 10047 19855 10053
rect 19797 10044 19809 10047
rect 19484 10016 19809 10044
rect 19484 10004 19490 10016
rect 19797 10013 19809 10016
rect 19843 10013 19855 10047
rect 19797 10007 19855 10013
rect 19981 10047 20039 10053
rect 19981 10013 19993 10047
rect 20027 10013 20039 10047
rect 19981 10007 20039 10013
rect 20076 10041 20134 10047
rect 20076 10007 20088 10041
rect 20122 10007 20134 10041
rect 20076 10001 20134 10007
rect 20162 10004 20168 10056
rect 20220 10053 20226 10056
rect 20220 10047 20243 10053
rect 20231 10013 20243 10047
rect 20220 10007 20243 10013
rect 20220 10004 20226 10007
rect 23566 10004 23572 10056
rect 23624 10044 23630 10056
rect 23661 10047 23719 10053
rect 23661 10044 23673 10047
rect 23624 10016 23673 10044
rect 23624 10004 23630 10016
rect 23661 10013 23673 10016
rect 23707 10044 23719 10047
rect 24394 10044 24400 10056
rect 23707 10016 24400 10044
rect 23707 10013 23719 10016
rect 23661 10007 23719 10013
rect 24394 10004 24400 10016
rect 24452 10004 24458 10056
rect 25314 10004 25320 10056
rect 25372 10044 25378 10056
rect 26145 10047 26203 10053
rect 26145 10044 26157 10047
rect 25372 10016 26157 10044
rect 25372 10004 25378 10016
rect 26145 10013 26157 10016
rect 26191 10013 26203 10047
rect 26326 10044 26332 10056
rect 26287 10016 26332 10044
rect 26145 10007 26203 10013
rect 26326 10004 26332 10016
rect 26384 10004 26390 10056
rect 26436 10053 26464 10084
rect 26421 10047 26479 10053
rect 26421 10013 26433 10047
rect 26467 10013 26479 10047
rect 26421 10007 26479 10013
rect 26513 10047 26571 10053
rect 26513 10013 26525 10047
rect 26559 10044 26571 10047
rect 26602 10044 26608 10056
rect 26559 10016 26608 10044
rect 26559 10013 26571 10016
rect 26513 10007 26571 10013
rect 26602 10004 26608 10016
rect 26660 10004 26666 10056
rect 27264 10053 27292 10152
rect 28534 10140 28540 10152
rect 28592 10140 28598 10192
rect 32953 10115 33011 10121
rect 27356 10084 31754 10112
rect 27249 10047 27307 10053
rect 27249 10013 27261 10047
rect 27295 10013 27307 10047
rect 27249 10007 27307 10013
rect 19334 9976 19340 9988
rect 13872 9948 16252 9976
rect 18432 9948 19340 9976
rect 13872 9936 13878 9948
rect 6012 9880 7052 9908
rect 7098 9868 7104 9920
rect 7156 9908 7162 9920
rect 7834 9908 7840 9920
rect 7156 9880 7840 9908
rect 7156 9868 7162 9880
rect 7834 9868 7840 9880
rect 7892 9868 7898 9920
rect 8113 9911 8171 9917
rect 8113 9877 8125 9911
rect 8159 9908 8171 9911
rect 8294 9908 8300 9920
rect 8159 9880 8300 9908
rect 8159 9877 8171 9880
rect 8113 9871 8171 9877
rect 8294 9868 8300 9880
rect 8352 9868 8358 9920
rect 10229 9911 10287 9917
rect 10229 9877 10241 9911
rect 10275 9908 10287 9911
rect 10962 9908 10968 9920
rect 10275 9880 10968 9908
rect 10275 9877 10287 9880
rect 10229 9871 10287 9877
rect 10962 9868 10968 9880
rect 11020 9868 11026 9920
rect 11974 9868 11980 9920
rect 12032 9868 12038 9920
rect 12710 9908 12716 9920
rect 12671 9880 12716 9908
rect 12710 9868 12716 9880
rect 12768 9868 12774 9920
rect 13538 9908 13544 9920
rect 13499 9880 13544 9908
rect 13538 9868 13544 9880
rect 13596 9868 13602 9920
rect 14182 9868 14188 9920
rect 14240 9908 14246 9920
rect 14645 9911 14703 9917
rect 14645 9908 14657 9911
rect 14240 9880 14657 9908
rect 14240 9868 14246 9880
rect 14645 9877 14657 9880
rect 14691 9877 14703 9911
rect 14645 9871 14703 9877
rect 15289 9911 15347 9917
rect 15289 9877 15301 9911
rect 15335 9908 15347 9911
rect 15470 9908 15476 9920
rect 15335 9880 15476 9908
rect 15335 9877 15347 9880
rect 15289 9871 15347 9877
rect 15470 9868 15476 9880
rect 15528 9868 15534 9920
rect 16224 9917 16252 9948
rect 19334 9936 19340 9948
rect 19392 9976 19398 9988
rect 19392 9948 20024 9976
rect 19392 9936 19398 9948
rect 16209 9911 16267 9917
rect 16209 9877 16221 9911
rect 16255 9908 16267 9911
rect 19794 9908 19800 9920
rect 16255 9880 19800 9908
rect 16255 9877 16267 9880
rect 16209 9871 16267 9877
rect 19794 9868 19800 9880
rect 19852 9868 19858 9920
rect 19996 9908 20024 9948
rect 20093 9920 20121 10001
rect 20441 9979 20499 9985
rect 20441 9945 20453 9979
rect 20487 9976 20499 9979
rect 21238 9979 21296 9985
rect 21238 9976 21250 9979
rect 20487 9948 21250 9976
rect 20487 9945 20499 9948
rect 20441 9939 20499 9945
rect 21238 9945 21250 9948
rect 21284 9945 21296 9979
rect 26620 9976 26648 10004
rect 27356 9976 27384 10084
rect 27522 10044 27528 10056
rect 27483 10016 27528 10044
rect 27522 10004 27528 10016
rect 27580 10004 27586 10056
rect 27617 10047 27675 10053
rect 27617 10013 27629 10047
rect 27663 10044 27675 10047
rect 28442 10044 28448 10056
rect 27663 10016 28448 10044
rect 27663 10013 27675 10016
rect 27617 10007 27675 10013
rect 28442 10004 28448 10016
rect 28500 10004 28506 10056
rect 28718 10044 28724 10056
rect 28679 10016 28724 10044
rect 28718 10004 28724 10016
rect 28776 10004 28782 10056
rect 28810 10004 28816 10056
rect 28868 10044 28874 10056
rect 28868 10016 28913 10044
rect 28868 10004 28874 10016
rect 28994 10004 29000 10056
rect 29052 10044 29058 10056
rect 29549 10047 29607 10053
rect 29549 10044 29561 10047
rect 29052 10016 29561 10044
rect 29052 10004 29058 10016
rect 29549 10013 29561 10016
rect 29595 10013 29607 10047
rect 29549 10007 29607 10013
rect 26620 9948 27384 9976
rect 27433 9979 27491 9985
rect 21238 9939 21296 9945
rect 27433 9945 27445 9979
rect 27479 9976 27491 9979
rect 27798 9976 27804 9988
rect 27479 9948 27804 9976
rect 27479 9945 27491 9948
rect 27433 9939 27491 9945
rect 27798 9936 27804 9948
rect 27856 9936 27862 9988
rect 31726 9976 31754 10084
rect 32953 10081 32965 10115
rect 32999 10112 33011 10115
rect 39022 10112 39028 10124
rect 32999 10084 39028 10112
rect 32999 10081 33011 10084
rect 32953 10075 33011 10081
rect 39022 10072 39028 10084
rect 39080 10072 39086 10124
rect 32697 10047 32755 10053
rect 32697 10013 32709 10047
rect 32743 10044 32755 10047
rect 33226 10044 33232 10056
rect 32743 10016 33232 10044
rect 32743 10013 32755 10016
rect 32697 10007 32755 10013
rect 33226 10004 33232 10016
rect 33284 10004 33290 10056
rect 34514 10004 34520 10056
rect 34572 10044 34578 10056
rect 34701 10047 34759 10053
rect 34701 10044 34713 10047
rect 34572 10016 34713 10044
rect 34572 10004 34578 10016
rect 34701 10013 34713 10016
rect 34747 10013 34759 10047
rect 34701 10007 34759 10013
rect 34885 10047 34943 10053
rect 34885 10013 34897 10047
rect 34931 10044 34943 10047
rect 35342 10044 35348 10056
rect 34931 10016 35348 10044
rect 34931 10013 34943 10016
rect 34885 10007 34943 10013
rect 35342 10004 35348 10016
rect 35400 10044 35406 10056
rect 35710 10044 35716 10056
rect 35400 10016 35716 10044
rect 35400 10004 35406 10016
rect 35710 10004 35716 10016
rect 35768 10004 35774 10056
rect 35802 10004 35808 10056
rect 35860 10044 35866 10056
rect 35897 10047 35955 10053
rect 35897 10044 35909 10047
rect 35860 10016 35909 10044
rect 35860 10004 35866 10016
rect 35897 10013 35909 10016
rect 35943 10013 35955 10047
rect 35897 10007 35955 10013
rect 36173 10047 36231 10053
rect 36173 10013 36185 10047
rect 36219 10013 36231 10047
rect 37090 10044 37096 10056
rect 37051 10016 37096 10044
rect 36173 10007 36231 10013
rect 34238 9976 34244 9988
rect 31726 9948 34244 9976
rect 34238 9936 34244 9948
rect 34296 9936 34302 9988
rect 20070 9908 20076 9920
rect 19996 9880 20076 9908
rect 20070 9868 20076 9880
rect 20128 9868 20134 9920
rect 20714 9868 20720 9920
rect 20772 9908 20778 9920
rect 21082 9908 21088 9920
rect 20772 9880 21088 9908
rect 20772 9868 20778 9880
rect 21082 9868 21088 9880
rect 21140 9868 21146 9920
rect 26786 9908 26792 9920
rect 26747 9880 26792 9908
rect 26786 9868 26792 9880
rect 26844 9868 26850 9920
rect 31386 9868 31392 9920
rect 31444 9908 31450 9920
rect 31573 9911 31631 9917
rect 31573 9908 31585 9911
rect 31444 9880 31585 9908
rect 31444 9868 31450 9880
rect 31573 9877 31585 9880
rect 31619 9877 31631 9911
rect 31573 9871 31631 9877
rect 34054 9868 34060 9920
rect 34112 9908 34118 9920
rect 34149 9911 34207 9917
rect 34149 9908 34161 9911
rect 34112 9880 34161 9908
rect 34112 9868 34118 9880
rect 34149 9877 34161 9880
rect 34195 9908 34207 9911
rect 36188 9908 36216 10007
rect 37090 10004 37096 10016
rect 37148 10004 37154 10056
rect 37185 10047 37243 10053
rect 37185 10013 37197 10047
rect 37231 10044 37243 10047
rect 37461 10047 37519 10053
rect 37231 10016 37412 10044
rect 37231 10013 37243 10016
rect 37185 10007 37243 10013
rect 36998 9936 37004 9988
rect 37056 9976 37062 9988
rect 37274 9976 37280 9988
rect 37056 9948 37280 9976
rect 37056 9936 37062 9948
rect 37274 9936 37280 9948
rect 37332 9936 37338 9988
rect 37384 9976 37412 10016
rect 37461 10013 37473 10047
rect 37507 10044 37519 10047
rect 37734 10044 37740 10056
rect 37507 10016 37740 10044
rect 37507 10013 37519 10016
rect 37461 10007 37519 10013
rect 37734 10004 37740 10016
rect 37792 10004 37798 10056
rect 38102 10044 38108 10056
rect 37844 10016 38108 10044
rect 37844 9976 37872 10016
rect 38102 10004 38108 10016
rect 38160 10004 38166 10056
rect 37384 9948 37872 9976
rect 37918 9936 37924 9988
rect 37976 9976 37982 9988
rect 37976 9948 38021 9976
rect 37976 9936 37982 9948
rect 37366 9908 37372 9920
rect 34195 9880 37372 9908
rect 34195 9877 34207 9880
rect 34149 9871 34207 9877
rect 37366 9868 37372 9880
rect 37424 9868 37430 9920
rect 1104 9818 68816 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 68816 9818
rect 1104 9744 68816 9766
rect 4154 9704 4160 9716
rect 3712 9676 4160 9704
rect 2240 9646 2452 9674
rect 2240 9636 2268 9646
rect 2235 9608 2268 9636
rect 2424 9636 2452 9646
rect 3712 9636 3740 9676
rect 4154 9664 4160 9676
rect 4212 9664 4218 9716
rect 5169 9707 5227 9713
rect 5169 9686 5181 9707
rect 5215 9686 5227 9707
rect 7561 9707 7619 9713
rect 5166 9674 5172 9686
rect 4614 9636 4620 9648
rect 2424 9608 3740 9636
rect 3804 9608 4620 9636
rect 2235 9580 2263 9608
rect 1762 9528 1768 9580
rect 1820 9568 1826 9580
rect 2041 9571 2099 9577
rect 2041 9568 2053 9571
rect 1820 9540 2053 9568
rect 1820 9528 1826 9540
rect 2041 9537 2053 9540
rect 2087 9537 2099 9571
rect 2041 9531 2099 9537
rect 2220 9574 2278 9580
rect 3804 9577 3832 9608
rect 4614 9596 4620 9608
rect 4672 9596 4678 9648
rect 5109 9646 5172 9674
rect 5166 9634 5172 9646
rect 5224 9634 5230 9686
rect 7561 9673 7573 9707
rect 7607 9704 7619 9707
rect 7650 9704 7656 9716
rect 7607 9676 7656 9704
rect 7607 9673 7619 9676
rect 7561 9667 7619 9673
rect 7650 9664 7656 9676
rect 7708 9664 7714 9716
rect 10962 9664 10968 9716
rect 11020 9704 11026 9716
rect 14274 9704 14280 9716
rect 11020 9676 14280 9704
rect 11020 9664 11026 9676
rect 14274 9664 14280 9676
rect 14332 9664 14338 9716
rect 18782 9664 18788 9716
rect 18840 9704 18846 9716
rect 19334 9704 19340 9716
rect 18840 9676 19340 9704
rect 18840 9664 18846 9676
rect 19334 9664 19340 9676
rect 19392 9664 19398 9716
rect 19518 9664 19524 9716
rect 19576 9704 19582 9716
rect 19613 9707 19671 9713
rect 19613 9704 19625 9707
rect 19576 9676 19625 9704
rect 19576 9664 19582 9676
rect 19613 9673 19625 9676
rect 19659 9673 19671 9707
rect 19613 9667 19671 9673
rect 20070 9664 20076 9716
rect 20128 9704 20134 9716
rect 20303 9707 20361 9713
rect 20303 9704 20315 9707
rect 20128 9676 20315 9704
rect 20128 9664 20134 9676
rect 20303 9673 20315 9676
rect 20349 9673 20361 9707
rect 32674 9704 32680 9716
rect 32635 9676 32680 9704
rect 20303 9667 20361 9673
rect 32674 9664 32680 9676
rect 32732 9704 32738 9716
rect 32732 9676 33456 9704
rect 32732 9664 32738 9676
rect 5258 9596 5264 9648
rect 5316 9636 5322 9648
rect 8294 9645 8300 9648
rect 8288 9636 8300 9645
rect 5316 9608 8156 9636
rect 8255 9608 8300 9636
rect 5316 9596 5322 9608
rect 4062 9577 4068 9580
rect 2220 9540 2232 9574
rect 2266 9540 2278 9574
rect 2220 9534 2278 9540
rect 2317 9571 2375 9577
rect 2317 9537 2329 9571
rect 2363 9537 2375 9571
rect 2317 9531 2375 9537
rect 2455 9571 2513 9577
rect 2455 9537 2467 9571
rect 2501 9568 2513 9571
rect 3789 9571 3847 9577
rect 2501 9540 3280 9568
rect 2501 9537 2513 9540
rect 2455 9531 2513 9537
rect 2332 9444 2360 9531
rect 2314 9392 2320 9444
rect 2372 9392 2378 9444
rect 1581 9367 1639 9373
rect 1581 9333 1593 9367
rect 1627 9364 1639 9367
rect 2406 9364 2412 9376
rect 1627 9336 2412 9364
rect 1627 9333 1639 9336
rect 1581 9327 1639 9333
rect 2406 9324 2412 9336
rect 2464 9324 2470 9376
rect 2682 9364 2688 9376
rect 2643 9336 2688 9364
rect 2682 9324 2688 9336
rect 2740 9324 2746 9376
rect 3252 9373 3280 9540
rect 3789 9537 3801 9571
rect 3835 9537 3847 9571
rect 3789 9531 3847 9537
rect 4056 9531 4068 9577
rect 4120 9568 4126 9580
rect 4120 9540 4156 9568
rect 4062 9528 4068 9531
rect 4120 9528 4126 9540
rect 5810 9528 5816 9580
rect 5868 9568 5874 9580
rect 7193 9571 7251 9577
rect 7193 9568 7205 9571
rect 5868 9540 7205 9568
rect 5868 9528 5874 9540
rect 7193 9537 7205 9540
rect 7239 9537 7251 9571
rect 7193 9531 7251 9537
rect 7377 9571 7435 9577
rect 7377 9537 7389 9571
rect 7423 9537 7435 9571
rect 7377 9531 7435 9537
rect 3237 9367 3295 9373
rect 3237 9333 3249 9367
rect 3283 9364 3295 9367
rect 7098 9364 7104 9376
rect 3283 9336 7104 9364
rect 3283 9333 3295 9336
rect 3237 9327 3295 9333
rect 7098 9324 7104 9336
rect 7156 9324 7162 9376
rect 7392 9364 7420 9531
rect 7558 9528 7564 9580
rect 7616 9568 7622 9580
rect 8021 9571 8079 9577
rect 8021 9568 8033 9571
rect 7616 9540 8033 9568
rect 7616 9528 7622 9540
rect 8021 9537 8033 9540
rect 8067 9537 8079 9571
rect 8128 9568 8156 9608
rect 8288 9599 8300 9608
rect 8294 9596 8300 9599
rect 8352 9596 8358 9648
rect 10229 9639 10287 9645
rect 10229 9636 10241 9639
rect 8404 9608 10241 9636
rect 8404 9568 8432 9608
rect 10229 9605 10241 9608
rect 10275 9605 10287 9639
rect 10229 9599 10287 9605
rect 10410 9596 10416 9648
rect 10468 9636 10474 9648
rect 17218 9636 17224 9648
rect 10468 9608 15884 9636
rect 10468 9596 10474 9608
rect 8128 9540 8432 9568
rect 8021 9531 8079 9537
rect 8754 9528 8760 9580
rect 8812 9568 8818 9580
rect 9950 9568 9956 9580
rect 8812 9540 9076 9568
rect 9911 9540 9956 9568
rect 8812 9528 8818 9540
rect 9048 9432 9076 9540
rect 9950 9528 9956 9540
rect 10008 9528 10014 9580
rect 10134 9568 10140 9580
rect 10095 9540 10140 9568
rect 10134 9528 10140 9540
rect 10192 9528 10198 9580
rect 10321 9571 10379 9577
rect 10321 9537 10333 9571
rect 10367 9568 10379 9571
rect 10594 9568 10600 9580
rect 10367 9540 10600 9568
rect 10367 9537 10379 9540
rect 10321 9531 10379 9537
rect 10594 9528 10600 9540
rect 10652 9528 10658 9580
rect 12158 9568 12164 9580
rect 12119 9540 12164 9568
rect 12158 9528 12164 9540
rect 12216 9528 12222 9580
rect 12345 9571 12403 9577
rect 12345 9537 12357 9571
rect 12391 9568 12403 9571
rect 12618 9568 12624 9580
rect 12391 9540 12624 9568
rect 12391 9537 12403 9540
rect 12345 9531 12403 9537
rect 12618 9528 12624 9540
rect 12676 9528 12682 9580
rect 12713 9571 12771 9577
rect 12713 9537 12725 9571
rect 12759 9537 12771 9571
rect 12713 9531 12771 9537
rect 12897 9571 12955 9577
rect 12897 9537 12909 9571
rect 12943 9568 12955 9571
rect 14470 9571 14528 9577
rect 14470 9568 14482 9571
rect 12943 9540 14482 9568
rect 12943 9537 12955 9540
rect 12897 9531 12955 9537
rect 14470 9537 14482 9540
rect 14516 9537 14528 9571
rect 15562 9568 15568 9580
rect 14470 9531 14528 9537
rect 14844 9540 15568 9568
rect 9858 9460 9864 9512
rect 9916 9500 9922 9512
rect 12437 9503 12495 9509
rect 12437 9500 12449 9503
rect 9916 9472 12449 9500
rect 9916 9460 9922 9472
rect 12437 9469 12449 9472
rect 12483 9469 12495 9503
rect 12437 9463 12495 9469
rect 12526 9460 12532 9512
rect 12584 9500 12590 9512
rect 12728 9500 12756 9531
rect 13354 9500 13360 9512
rect 12584 9472 12629 9500
rect 12728 9472 13360 9500
rect 12584 9460 12590 9472
rect 13354 9460 13360 9472
rect 13412 9460 13418 9512
rect 14734 9500 14740 9512
rect 14695 9472 14740 9500
rect 14734 9460 14740 9472
rect 14792 9460 14798 9512
rect 9048 9404 12434 9432
rect 9398 9364 9404 9376
rect 7392 9336 9404 9364
rect 9398 9324 9404 9336
rect 9456 9324 9462 9376
rect 10502 9364 10508 9376
rect 10463 9336 10508 9364
rect 10502 9324 10508 9336
rect 10560 9324 10566 9376
rect 11514 9364 11520 9376
rect 11475 9336 11520 9364
rect 11514 9324 11520 9336
rect 11572 9324 11578 9376
rect 12406 9364 12434 9404
rect 13188 9404 13860 9432
rect 13188 9364 13216 9404
rect 13354 9364 13360 9376
rect 12406 9336 13216 9364
rect 13315 9336 13360 9364
rect 13354 9324 13360 9336
rect 13412 9324 13418 9376
rect 13832 9364 13860 9404
rect 14844 9364 14872 9540
rect 15562 9528 15568 9540
rect 15620 9528 15626 9580
rect 15856 9577 15884 9608
rect 15948 9608 17224 9636
rect 15948 9577 15976 9608
rect 17218 9596 17224 9608
rect 17276 9596 17282 9648
rect 18046 9596 18052 9648
rect 18104 9636 18110 9648
rect 19429 9639 19487 9645
rect 18104 9608 18644 9636
rect 18104 9596 18110 9608
rect 15841 9571 15899 9577
rect 15841 9537 15853 9571
rect 15887 9537 15899 9571
rect 15841 9531 15899 9537
rect 15933 9571 15991 9577
rect 15933 9537 15945 9571
rect 15979 9537 15991 9571
rect 15933 9531 15991 9537
rect 16117 9571 16175 9577
rect 16117 9537 16129 9571
rect 16163 9568 16175 9571
rect 16390 9568 16396 9580
rect 16163 9540 16396 9568
rect 16163 9537 16175 9540
rect 16117 9531 16175 9537
rect 16390 9528 16396 9540
rect 16448 9528 16454 9580
rect 17862 9568 17868 9580
rect 17823 9540 17868 9568
rect 17862 9528 17868 9540
rect 17920 9528 17926 9580
rect 17957 9571 18015 9577
rect 17957 9537 17969 9571
rect 18003 9537 18015 9571
rect 18414 9568 18420 9580
rect 18375 9540 18420 9568
rect 17957 9531 18015 9537
rect 15286 9460 15292 9512
rect 15344 9500 15350 9512
rect 15749 9503 15807 9509
rect 15749 9500 15761 9503
rect 15344 9472 15761 9500
rect 15344 9460 15350 9472
rect 15749 9469 15761 9472
rect 15795 9500 15807 9503
rect 16942 9500 16948 9512
rect 15795 9472 16948 9500
rect 15795 9469 15807 9472
rect 15749 9463 15807 9469
rect 16942 9460 16948 9472
rect 17000 9460 17006 9512
rect 17972 9500 18000 9531
rect 18414 9528 18420 9540
rect 18472 9528 18478 9580
rect 18616 9577 18644 9608
rect 19429 9605 19441 9639
rect 19475 9636 19487 9639
rect 20622 9636 20628 9648
rect 19475 9608 20628 9636
rect 19475 9605 19487 9608
rect 19429 9599 19487 9605
rect 20622 9596 20628 9608
rect 20680 9596 20686 9648
rect 22186 9636 22192 9648
rect 21836 9608 22192 9636
rect 18601 9571 18659 9577
rect 18601 9537 18613 9571
rect 18647 9537 18659 9571
rect 18601 9531 18659 9537
rect 19245 9571 19303 9577
rect 19245 9537 19257 9571
rect 19291 9568 19303 9571
rect 19518 9568 19524 9580
rect 19291 9540 19524 9568
rect 19291 9537 19303 9540
rect 19245 9531 19303 9537
rect 19518 9528 19524 9540
rect 19576 9528 19582 9580
rect 21836 9577 21864 9608
rect 22186 9596 22192 9608
rect 22244 9636 22250 9648
rect 22465 9639 22523 9645
rect 22465 9636 22477 9639
rect 22244 9608 22477 9636
rect 22244 9596 22250 9608
rect 22465 9605 22477 9608
rect 22511 9605 22523 9639
rect 24854 9636 24860 9648
rect 22465 9599 22523 9605
rect 24504 9608 24860 9636
rect 21821 9571 21879 9577
rect 19996 9540 20300 9568
rect 19996 9500 20024 9540
rect 17972 9472 20024 9500
rect 20070 9460 20076 9512
rect 20128 9500 20134 9512
rect 20272 9500 20300 9540
rect 21821 9537 21833 9571
rect 21867 9537 21879 9571
rect 21821 9531 21879 9537
rect 22005 9571 22063 9577
rect 22005 9537 22017 9571
rect 22051 9537 22063 9571
rect 22005 9531 22063 9537
rect 20438 9500 20444 9512
rect 20128 9472 20173 9500
rect 20272 9472 20444 9500
rect 20128 9460 20134 9472
rect 20438 9460 20444 9472
rect 20496 9460 20502 9512
rect 21542 9460 21548 9512
rect 21600 9500 21606 9512
rect 22020 9500 22048 9531
rect 22922 9528 22928 9580
rect 22980 9568 22986 9580
rect 23109 9571 23167 9577
rect 23109 9568 23121 9571
rect 22980 9540 23121 9568
rect 22980 9528 22986 9540
rect 23109 9537 23121 9540
rect 23155 9568 23167 9571
rect 24302 9568 24308 9580
rect 23155 9540 24308 9568
rect 23155 9537 23167 9540
rect 23109 9531 23167 9537
rect 24302 9528 24308 9540
rect 24360 9568 24366 9580
rect 24504 9577 24532 9608
rect 24854 9596 24860 9608
rect 24912 9596 24918 9648
rect 25406 9596 25412 9648
rect 25464 9636 25470 9648
rect 25685 9639 25743 9645
rect 25685 9636 25697 9639
rect 25464 9608 25697 9636
rect 25464 9596 25470 9608
rect 25685 9605 25697 9608
rect 25731 9605 25743 9639
rect 25685 9599 25743 9605
rect 26053 9639 26111 9645
rect 26053 9605 26065 9639
rect 26099 9636 26111 9639
rect 26326 9636 26332 9648
rect 26099 9608 26332 9636
rect 26099 9605 26111 9608
rect 26053 9599 26111 9605
rect 26326 9596 26332 9608
rect 26384 9596 26390 9648
rect 26510 9596 26516 9648
rect 26568 9636 26574 9648
rect 30092 9639 30150 9645
rect 26568 9608 29868 9636
rect 26568 9596 26574 9608
rect 24397 9571 24455 9577
rect 24397 9568 24409 9571
rect 24360 9540 24409 9568
rect 24360 9528 24366 9540
rect 24397 9537 24409 9540
rect 24443 9537 24455 9571
rect 24397 9531 24455 9537
rect 24489 9571 24547 9577
rect 24489 9537 24501 9571
rect 24535 9537 24547 9571
rect 24489 9531 24547 9537
rect 24578 9528 24584 9580
rect 24636 9568 24642 9580
rect 24765 9571 24823 9577
rect 24636 9540 24681 9568
rect 24636 9528 24642 9540
rect 24765 9537 24777 9571
rect 24811 9568 24823 9571
rect 25314 9568 25320 9580
rect 24811 9540 25320 9568
rect 24811 9537 24823 9540
rect 24765 9531 24823 9537
rect 21600 9472 22048 9500
rect 23661 9503 23719 9509
rect 21600 9460 21606 9472
rect 23661 9469 23673 9503
rect 23707 9500 23719 9503
rect 24780 9500 24808 9531
rect 25314 9528 25320 9540
rect 25372 9528 25378 9580
rect 25869 9571 25927 9577
rect 25869 9537 25881 9571
rect 25915 9568 25927 9571
rect 27430 9568 27436 9580
rect 25915 9540 27436 9568
rect 25915 9537 25927 9540
rect 25869 9531 25927 9537
rect 27430 9528 27436 9540
rect 27488 9528 27494 9580
rect 27982 9568 27988 9580
rect 27943 9540 27988 9568
rect 27982 9528 27988 9540
rect 28040 9528 28046 9580
rect 28261 9571 28319 9577
rect 28261 9537 28273 9571
rect 28307 9537 28319 9571
rect 28902 9568 28908 9580
rect 28863 9540 28908 9568
rect 28261 9531 28319 9537
rect 23707 9472 24808 9500
rect 23707 9469 23719 9472
rect 23661 9463 23719 9469
rect 25590 9460 25596 9512
rect 25648 9500 25654 9512
rect 26973 9503 27031 9509
rect 26973 9500 26985 9503
rect 25648 9472 26985 9500
rect 25648 9460 25654 9472
rect 26973 9469 26985 9472
rect 27019 9469 27031 9503
rect 28074 9500 28080 9512
rect 28035 9472 28080 9500
rect 26973 9463 27031 9469
rect 28074 9460 28080 9472
rect 28132 9460 28138 9512
rect 28276 9500 28304 9531
rect 28902 9528 28908 9540
rect 28960 9528 28966 9580
rect 28994 9528 29000 9580
rect 29052 9568 29058 9580
rect 29089 9571 29147 9577
rect 29089 9568 29101 9571
rect 29052 9540 29101 9568
rect 29052 9528 29058 9540
rect 29089 9537 29101 9540
rect 29135 9537 29147 9571
rect 29089 9531 29147 9537
rect 29181 9571 29239 9577
rect 29181 9537 29193 9571
rect 29227 9568 29239 9571
rect 29730 9568 29736 9580
rect 29227 9540 29736 9568
rect 29227 9537 29239 9540
rect 29181 9531 29239 9537
rect 29730 9528 29736 9540
rect 29788 9528 29794 9580
rect 29840 9577 29868 9608
rect 30092 9605 30104 9639
rect 30138 9636 30150 9639
rect 33137 9639 33195 9645
rect 33137 9636 33149 9639
rect 30138 9608 33149 9636
rect 30138 9605 30150 9608
rect 30092 9599 30150 9605
rect 33137 9605 33149 9608
rect 33183 9605 33195 9639
rect 33137 9599 33195 9605
rect 33428 9577 33456 9676
rect 34238 9664 34244 9716
rect 34296 9704 34302 9716
rect 37277 9707 37335 9713
rect 37277 9704 37289 9707
rect 34296 9676 37289 9704
rect 34296 9664 34302 9676
rect 37277 9673 37289 9676
rect 37323 9673 37335 9707
rect 37277 9667 37335 9673
rect 34333 9639 34391 9645
rect 34333 9605 34345 9639
rect 34379 9636 34391 9639
rect 34514 9636 34520 9648
rect 34379 9608 34520 9636
rect 34379 9605 34391 9608
rect 34333 9599 34391 9605
rect 34514 9596 34520 9608
rect 34572 9596 34578 9648
rect 37292 9636 37320 9667
rect 38378 9636 38384 9648
rect 37292 9608 38384 9636
rect 29825 9571 29883 9577
rect 29825 9537 29837 9571
rect 29871 9537 29883 9571
rect 29825 9531 29883 9537
rect 33413 9571 33471 9577
rect 33413 9537 33425 9571
rect 33459 9537 33471 9571
rect 33413 9531 33471 9537
rect 33505 9571 33563 9577
rect 33505 9537 33517 9571
rect 33551 9537 33563 9571
rect 33505 9531 33563 9537
rect 29546 9500 29552 9512
rect 28276 9472 29552 9500
rect 29546 9460 29552 9472
rect 29604 9460 29610 9512
rect 18322 9432 18328 9444
rect 17144 9404 18328 9432
rect 17144 9376 17172 9404
rect 18322 9392 18328 9404
rect 18380 9392 18386 9444
rect 18693 9435 18751 9441
rect 18693 9401 18705 9435
rect 18739 9432 18751 9435
rect 28166 9432 28172 9444
rect 18739 9404 28172 9432
rect 18739 9401 18751 9404
rect 18693 9395 18751 9401
rect 28166 9392 28172 9404
rect 28224 9392 28230 9444
rect 28442 9432 28448 9444
rect 28403 9404 28448 9432
rect 28442 9392 28448 9404
rect 28500 9392 28506 9444
rect 29270 9432 29276 9444
rect 28736 9404 29276 9432
rect 15378 9364 15384 9376
rect 13832 9336 14872 9364
rect 15339 9336 15384 9364
rect 15378 9324 15384 9336
rect 15436 9324 15442 9376
rect 17126 9364 17132 9376
rect 17087 9336 17132 9364
rect 17126 9324 17132 9336
rect 17184 9324 17190 9376
rect 17310 9324 17316 9376
rect 17368 9364 17374 9376
rect 17589 9367 17647 9373
rect 17589 9364 17601 9367
rect 17368 9336 17601 9364
rect 17368 9324 17374 9336
rect 17589 9333 17601 9336
rect 17635 9333 17647 9367
rect 17770 9364 17776 9376
rect 17731 9336 17776 9364
rect 17589 9327 17647 9333
rect 17770 9324 17776 9336
rect 17828 9324 17834 9376
rect 20070 9324 20076 9376
rect 20128 9364 20134 9376
rect 21913 9367 21971 9373
rect 21913 9364 21925 9367
rect 20128 9336 21925 9364
rect 20128 9324 20134 9336
rect 21913 9333 21925 9336
rect 21959 9333 21971 9367
rect 24118 9364 24124 9376
rect 24079 9336 24124 9364
rect 21913 9327 21971 9333
rect 24118 9324 24124 9336
rect 24176 9324 24182 9376
rect 28261 9367 28319 9373
rect 28261 9333 28273 9367
rect 28307 9364 28319 9367
rect 28736 9364 28764 9404
rect 29270 9392 29276 9404
rect 29328 9392 29334 9444
rect 33520 9432 33548 9531
rect 33594 9528 33600 9580
rect 33652 9568 33658 9580
rect 33781 9571 33839 9577
rect 33652 9540 33697 9568
rect 33652 9528 33658 9540
rect 33781 9537 33793 9571
rect 33827 9568 33839 9571
rect 34422 9568 34428 9580
rect 33827 9540 34428 9568
rect 33827 9537 33839 9540
rect 33781 9531 33839 9537
rect 34422 9528 34428 9540
rect 34480 9568 34486 9580
rect 34606 9568 34612 9580
rect 34480 9540 34612 9568
rect 34480 9528 34486 9540
rect 34606 9528 34612 9540
rect 34664 9528 34670 9580
rect 34698 9528 34704 9580
rect 34756 9568 34762 9580
rect 34977 9571 35035 9577
rect 34977 9568 34989 9571
rect 34756 9540 34989 9568
rect 34756 9528 34762 9540
rect 34977 9537 34989 9540
rect 35023 9537 35035 9571
rect 35710 9568 35716 9580
rect 35671 9540 35716 9568
rect 34977 9531 35035 9537
rect 35710 9528 35716 9540
rect 35768 9528 35774 9580
rect 37550 9528 37556 9580
rect 37608 9568 37614 9580
rect 37829 9571 37887 9577
rect 37829 9568 37841 9571
rect 37608 9540 37841 9568
rect 37608 9528 37614 9540
rect 37829 9537 37841 9540
rect 37875 9537 37887 9571
rect 38010 9568 38016 9580
rect 37971 9540 38016 9568
rect 37829 9531 37887 9537
rect 38010 9528 38016 9540
rect 38068 9528 38074 9580
rect 38212 9577 38240 9608
rect 38378 9596 38384 9608
rect 38436 9596 38442 9648
rect 38473 9639 38531 9645
rect 38473 9605 38485 9639
rect 38519 9636 38531 9639
rect 39270 9639 39328 9645
rect 39270 9636 39282 9639
rect 38519 9608 39282 9636
rect 38519 9605 38531 9608
rect 38473 9599 38531 9605
rect 39270 9605 39282 9608
rect 39316 9605 39328 9639
rect 39270 9599 39328 9605
rect 38105 9571 38163 9577
rect 38105 9537 38117 9571
rect 38151 9537 38163 9571
rect 38105 9531 38163 9537
rect 38197 9571 38255 9577
rect 38197 9537 38209 9571
rect 38243 9537 38255 9571
rect 39022 9568 39028 9580
rect 38983 9540 39028 9568
rect 38197 9531 38255 9537
rect 34514 9460 34520 9512
rect 34572 9500 34578 9512
rect 35437 9503 35495 9509
rect 35437 9500 35449 9503
rect 34572 9472 35449 9500
rect 34572 9460 34578 9472
rect 35437 9469 35449 9472
rect 35483 9469 35495 9503
rect 35437 9463 35495 9469
rect 35618 9460 35624 9512
rect 35676 9500 35682 9512
rect 37182 9500 37188 9512
rect 35676 9472 37188 9500
rect 35676 9460 35682 9472
rect 37182 9460 37188 9472
rect 37240 9500 37246 9512
rect 38120 9500 38148 9531
rect 39022 9528 39028 9540
rect 39080 9528 39086 9580
rect 37240 9472 38148 9500
rect 37240 9460 37246 9472
rect 35526 9432 35532 9444
rect 33520 9404 35532 9432
rect 35526 9392 35532 9404
rect 35584 9392 35590 9444
rect 29086 9364 29092 9376
rect 28307 9336 28764 9364
rect 29047 9336 29092 9364
rect 28307 9333 28319 9336
rect 28261 9327 28319 9333
rect 29086 9324 29092 9336
rect 29144 9324 29150 9376
rect 29362 9364 29368 9376
rect 29323 9336 29368 9364
rect 29362 9324 29368 9336
rect 29420 9324 29426 9376
rect 31110 9324 31116 9376
rect 31168 9364 31174 9376
rect 31205 9367 31263 9373
rect 31205 9364 31217 9367
rect 31168 9336 31217 9364
rect 31168 9324 31174 9336
rect 31205 9333 31217 9336
rect 31251 9333 31263 9367
rect 31205 9327 31263 9333
rect 34793 9367 34851 9373
rect 34793 9333 34805 9367
rect 34839 9364 34851 9367
rect 35894 9364 35900 9376
rect 34839 9336 35900 9364
rect 34839 9333 34851 9336
rect 34793 9327 34851 9333
rect 35894 9324 35900 9336
rect 35952 9364 35958 9376
rect 37182 9364 37188 9376
rect 35952 9336 37188 9364
rect 35952 9324 35958 9336
rect 37182 9324 37188 9336
rect 37240 9324 37246 9376
rect 37826 9324 37832 9376
rect 37884 9364 37890 9376
rect 40405 9367 40463 9373
rect 40405 9364 40417 9367
rect 37884 9336 40417 9364
rect 37884 9324 37890 9336
rect 40405 9333 40417 9336
rect 40451 9333 40463 9367
rect 40405 9327 40463 9333
rect 1104 9274 68816 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 65654 9274
rect 65706 9222 65718 9274
rect 65770 9222 65782 9274
rect 65834 9222 65846 9274
rect 65898 9222 65910 9274
rect 65962 9222 68816 9274
rect 1104 9200 68816 9222
rect 3053 9163 3111 9169
rect 3053 9160 3065 9163
rect 2746 9132 3065 9160
rect 2314 9024 2320 9036
rect 2148 8996 2320 9024
rect 1762 8916 1768 8968
rect 1820 8956 1826 8968
rect 2148 8965 2176 8996
rect 2314 8984 2320 8996
rect 2372 8984 2378 9036
rect 1857 8959 1915 8965
rect 1857 8956 1869 8959
rect 1820 8928 1869 8956
rect 1820 8916 1826 8928
rect 1857 8925 1869 8928
rect 1903 8925 1915 8959
rect 1857 8919 1915 8925
rect 2041 8959 2099 8965
rect 2041 8925 2053 8959
rect 2087 8925 2099 8959
rect 2041 8919 2099 8925
rect 2133 8959 2191 8965
rect 2133 8925 2145 8959
rect 2179 8925 2191 8959
rect 2133 8919 2191 8925
rect 2225 8959 2283 8965
rect 2225 8925 2237 8959
rect 2271 8956 2283 8959
rect 2746 8956 2774 9132
rect 3053 9129 3065 9132
rect 3099 9160 3111 9163
rect 3234 9160 3240 9172
rect 3099 9132 3240 9160
rect 3099 9129 3111 9132
rect 3053 9123 3111 9129
rect 3234 9120 3240 9132
rect 3292 9120 3298 9172
rect 6914 9120 6920 9172
rect 6972 9160 6978 9172
rect 7009 9163 7067 9169
rect 7009 9160 7021 9163
rect 6972 9132 7021 9160
rect 6972 9120 6978 9132
rect 7009 9129 7021 9132
rect 7055 9160 7067 9163
rect 9950 9160 9956 9172
rect 7055 9132 9956 9160
rect 7055 9129 7067 9132
rect 7009 9123 7067 9129
rect 9950 9120 9956 9132
rect 10008 9120 10014 9172
rect 12526 9120 12532 9172
rect 12584 9160 12590 9172
rect 15286 9160 15292 9172
rect 12584 9132 15292 9160
rect 12584 9120 12590 9132
rect 15286 9120 15292 9132
rect 15344 9120 15350 9172
rect 15562 9160 15568 9172
rect 15523 9132 15568 9160
rect 15562 9120 15568 9132
rect 15620 9120 15626 9172
rect 17678 9160 17684 9172
rect 15672 9132 16988 9160
rect 17639 9132 17684 9160
rect 8110 9052 8116 9104
rect 8168 9092 8174 9104
rect 9858 9092 9864 9104
rect 8168 9064 9864 9092
rect 8168 9052 8174 9064
rect 9858 9052 9864 9064
rect 9916 9052 9922 9104
rect 12066 9052 12072 9104
rect 12124 9092 12130 9104
rect 12124 9064 12756 9092
rect 12124 9052 12130 9064
rect 11974 8984 11980 9036
rect 12032 9024 12038 9036
rect 12345 9027 12403 9033
rect 12345 9024 12357 9027
rect 12032 8996 12357 9024
rect 12032 8984 12038 8996
rect 12345 8993 12357 8996
rect 12391 8993 12403 9027
rect 12345 8987 12403 8993
rect 12434 8984 12440 9036
rect 12492 9024 12498 9036
rect 12492 8996 12537 9024
rect 12492 8984 12498 8996
rect 4157 8959 4215 8965
rect 4157 8956 4169 8959
rect 2271 8928 2774 8956
rect 3436 8928 4169 8956
rect 2271 8925 2283 8928
rect 2225 8919 2283 8925
rect 2056 8888 2084 8919
rect 3436 8888 3464 8928
rect 4157 8925 4169 8928
rect 4203 8925 4215 8959
rect 4157 8919 4215 8925
rect 4614 8916 4620 8968
rect 4672 8956 4678 8968
rect 5629 8959 5687 8965
rect 5629 8956 5641 8959
rect 4672 8928 5641 8956
rect 4672 8916 4678 8928
rect 5629 8925 5641 8928
rect 5675 8925 5687 8959
rect 5629 8919 5687 8925
rect 5896 8959 5954 8965
rect 5896 8925 5908 8959
rect 5942 8956 5954 8959
rect 6362 8956 6368 8968
rect 5942 8928 6368 8956
rect 5942 8925 5954 8928
rect 5896 8919 5954 8925
rect 6362 8916 6368 8928
rect 6420 8916 6426 8968
rect 10870 8916 10876 8968
rect 10928 8956 10934 8968
rect 12728 8965 12756 9064
rect 13630 9052 13636 9104
rect 13688 9092 13694 9104
rect 15105 9095 15163 9101
rect 15105 9092 15117 9095
rect 13688 9064 15117 9092
rect 13688 9052 13694 9064
rect 15105 9061 15117 9064
rect 15151 9061 15163 9095
rect 15105 9055 15163 9061
rect 13541 9027 13599 9033
rect 13541 8993 13553 9027
rect 13587 9024 13599 9027
rect 15010 9024 15016 9036
rect 13587 8996 15016 9024
rect 13587 8993 13599 8996
rect 13541 8987 13599 8993
rect 15010 8984 15016 8996
rect 15068 8984 15074 9036
rect 15672 9024 15700 9132
rect 16960 9033 16988 9132
rect 17678 9120 17684 9132
rect 17736 9120 17742 9172
rect 18616 9132 24532 9160
rect 18616 9101 18644 9132
rect 18601 9095 18659 9101
rect 18601 9061 18613 9095
rect 18647 9061 18659 9095
rect 19518 9092 19524 9104
rect 19479 9064 19524 9092
rect 18601 9055 18659 9061
rect 19518 9052 19524 9064
rect 19576 9092 19582 9104
rect 20346 9092 20352 9104
rect 19576 9064 20352 9092
rect 19576 9052 19582 9064
rect 20346 9052 20352 9064
rect 20404 9052 20410 9104
rect 15120 8996 15700 9024
rect 16945 9027 17003 9033
rect 11517 8959 11575 8965
rect 11517 8956 11529 8959
rect 10928 8928 11529 8956
rect 10928 8916 10934 8928
rect 11517 8925 11529 8928
rect 11563 8925 11575 8959
rect 11517 8919 11575 8925
rect 12161 8959 12219 8965
rect 12161 8925 12173 8959
rect 12207 8925 12219 8959
rect 12161 8919 12219 8925
rect 12529 8959 12587 8965
rect 12529 8925 12541 8959
rect 12575 8925 12587 8959
rect 12529 8919 12587 8925
rect 12713 8959 12771 8965
rect 12713 8925 12725 8959
rect 12759 8956 12771 8959
rect 14274 8956 14280 8968
rect 12759 8928 14280 8956
rect 12759 8925 12771 8928
rect 12713 8919 12771 8925
rect 3786 8888 3792 8900
rect 2056 8860 3464 8888
rect 3747 8860 3792 8888
rect 3786 8848 3792 8860
rect 3844 8848 3850 8900
rect 3973 8891 4031 8897
rect 3973 8857 3985 8891
rect 4019 8888 4031 8891
rect 5166 8888 5172 8900
rect 4019 8860 5172 8888
rect 4019 8857 4031 8860
rect 3973 8851 4031 8857
rect 5166 8848 5172 8860
rect 5224 8848 5230 8900
rect 5442 8848 5448 8900
rect 5500 8888 5506 8900
rect 10318 8888 10324 8900
rect 5500 8860 10324 8888
rect 5500 8848 5506 8860
rect 10318 8848 10324 8860
rect 10376 8848 10382 8900
rect 11272 8891 11330 8897
rect 11272 8857 11284 8891
rect 11318 8888 11330 8891
rect 11977 8891 12035 8897
rect 11977 8888 11989 8891
rect 11318 8860 11989 8888
rect 11318 8857 11330 8860
rect 11272 8851 11330 8857
rect 11977 8857 11989 8860
rect 12023 8857 12035 8891
rect 11977 8851 12035 8857
rect 2501 8823 2559 8829
rect 2501 8789 2513 8823
rect 2547 8820 2559 8823
rect 4062 8820 4068 8832
rect 2547 8792 4068 8820
rect 2547 8789 2559 8792
rect 2501 8783 2559 8789
rect 4062 8780 4068 8792
rect 4120 8780 4126 8832
rect 4709 8823 4767 8829
rect 4709 8789 4721 8823
rect 4755 8820 4767 8823
rect 5074 8820 5080 8832
rect 4755 8792 5080 8820
rect 4755 8789 4767 8792
rect 4709 8783 4767 8789
rect 5074 8780 5080 8792
rect 5132 8780 5138 8832
rect 7282 8780 7288 8832
rect 7340 8820 7346 8832
rect 7469 8823 7527 8829
rect 7469 8820 7481 8823
rect 7340 8792 7481 8820
rect 7340 8780 7346 8792
rect 7469 8789 7481 8792
rect 7515 8789 7527 8823
rect 7469 8783 7527 8789
rect 8478 8780 8484 8832
rect 8536 8820 8542 8832
rect 10137 8823 10195 8829
rect 10137 8820 10149 8823
rect 8536 8792 10149 8820
rect 8536 8780 8542 8792
rect 10137 8789 10149 8792
rect 10183 8820 10195 8823
rect 12176 8820 12204 8919
rect 10183 8792 12204 8820
rect 12544 8820 12572 8919
rect 14274 8916 14280 8928
rect 14332 8916 14338 8968
rect 14553 8959 14611 8965
rect 14553 8925 14565 8959
rect 14599 8925 14611 8959
rect 14553 8919 14611 8925
rect 14568 8888 14596 8919
rect 14734 8916 14740 8968
rect 14792 8956 14798 8968
rect 15120 8956 15148 8996
rect 16945 8993 16957 9027
rect 16991 9024 17003 9027
rect 19978 9024 19984 9036
rect 16991 8996 19984 9024
rect 16991 8993 17003 8996
rect 16945 8987 17003 8993
rect 19978 8984 19984 8996
rect 20036 8984 20042 9036
rect 20530 9024 20536 9036
rect 20088 8996 20536 9024
rect 14792 8928 15148 8956
rect 14792 8916 14798 8928
rect 15378 8916 15384 8968
rect 15436 8956 15442 8968
rect 16678 8959 16736 8965
rect 16678 8956 16690 8959
rect 15436 8928 16690 8956
rect 15436 8916 15442 8928
rect 16678 8925 16690 8928
rect 16724 8925 16736 8959
rect 17770 8956 17776 8968
rect 17731 8928 17776 8956
rect 16678 8919 16736 8925
rect 17770 8916 17776 8928
rect 17828 8916 17834 8968
rect 17865 8959 17923 8965
rect 17865 8925 17877 8959
rect 17911 8925 17923 8959
rect 17865 8919 17923 8925
rect 16758 8888 16764 8900
rect 14568 8860 16764 8888
rect 16758 8848 16764 8860
rect 16816 8848 16822 8900
rect 17218 8820 17224 8832
rect 12544 8792 17224 8820
rect 10183 8789 10195 8792
rect 10137 8783 10195 8789
rect 17218 8780 17224 8792
rect 17276 8780 17282 8832
rect 17494 8820 17500 8832
rect 17455 8792 17500 8820
rect 17494 8780 17500 8792
rect 17552 8780 17558 8832
rect 17880 8820 17908 8919
rect 18138 8916 18144 8968
rect 18196 8956 18202 8968
rect 18414 8956 18420 8968
rect 18196 8928 18420 8956
rect 18196 8916 18202 8928
rect 18414 8916 18420 8928
rect 18472 8916 18478 8968
rect 18509 8959 18567 8965
rect 18509 8925 18521 8959
rect 18555 8925 18567 8959
rect 18509 8919 18567 8925
rect 19337 8959 19395 8965
rect 19337 8925 19349 8959
rect 19383 8925 19395 8959
rect 19337 8919 19395 8925
rect 17954 8848 17960 8900
rect 18012 8888 18018 8900
rect 18524 8888 18552 8919
rect 18012 8860 18552 8888
rect 19352 8888 19380 8919
rect 19886 8916 19892 8968
rect 19944 8956 19950 8968
rect 20088 8956 20116 8996
rect 20530 8984 20536 8996
rect 20588 8984 20594 9036
rect 24504 9024 24532 9132
rect 24578 9120 24584 9172
rect 24636 9160 24642 9172
rect 24765 9163 24823 9169
rect 24765 9160 24777 9163
rect 24636 9132 24777 9160
rect 24636 9120 24642 9132
rect 24765 9129 24777 9132
rect 24811 9129 24823 9163
rect 25314 9160 25320 9172
rect 25227 9132 25320 9160
rect 24765 9123 24823 9129
rect 25314 9120 25320 9132
rect 25372 9160 25378 9172
rect 27430 9160 27436 9172
rect 25372 9132 27108 9160
rect 27391 9132 27436 9160
rect 25372 9120 25378 9132
rect 27080 9024 27108 9132
rect 27430 9120 27436 9132
rect 27488 9120 27494 9172
rect 28813 9163 28871 9169
rect 28813 9129 28825 9163
rect 28859 9160 28871 9163
rect 28902 9160 28908 9172
rect 28859 9132 28908 9160
rect 28859 9129 28871 9132
rect 28813 9123 28871 9129
rect 28902 9120 28908 9132
rect 28960 9120 28966 9172
rect 30834 9160 30840 9172
rect 30795 9132 30840 9160
rect 30834 9120 30840 9132
rect 30892 9120 30898 9172
rect 33137 9163 33195 9169
rect 33137 9129 33149 9163
rect 33183 9160 33195 9163
rect 33594 9160 33600 9172
rect 33183 9132 33600 9160
rect 33183 9129 33195 9132
rect 33137 9123 33195 9129
rect 33594 9120 33600 9132
rect 33652 9120 33658 9172
rect 34606 9120 34612 9172
rect 34664 9160 34670 9172
rect 35250 9160 35256 9172
rect 34664 9132 35256 9160
rect 34664 9120 34670 9132
rect 35250 9120 35256 9132
rect 35308 9120 35314 9172
rect 38010 9160 38016 9172
rect 37971 9132 38016 9160
rect 38010 9120 38016 9132
rect 38068 9120 38074 9172
rect 29730 9052 29736 9104
rect 29788 9092 29794 9104
rect 36633 9095 36691 9101
rect 36633 9092 36645 9095
rect 29788 9064 36645 9092
rect 29788 9052 29794 9064
rect 36633 9061 36645 9064
rect 36679 9061 36691 9095
rect 36633 9055 36691 9061
rect 33318 9024 33324 9036
rect 24504 8996 26188 9024
rect 27080 8996 33324 9024
rect 19944 8928 20116 8956
rect 20165 8959 20223 8965
rect 19944 8916 19950 8928
rect 20165 8925 20177 8959
rect 20211 8956 20223 8959
rect 21910 8956 21916 8968
rect 20211 8928 21916 8956
rect 20211 8925 20223 8928
rect 20165 8919 20223 8925
rect 21910 8916 21916 8928
rect 21968 8916 21974 8968
rect 22097 8959 22155 8965
rect 22097 8925 22109 8959
rect 22143 8956 22155 8959
rect 23382 8956 23388 8968
rect 22143 8928 23388 8956
rect 22143 8925 22155 8928
rect 22097 8919 22155 8925
rect 23382 8916 23388 8928
rect 23440 8956 23446 8968
rect 26053 8959 26111 8965
rect 26053 8956 26065 8959
rect 23440 8928 26065 8956
rect 23440 8916 23446 8928
rect 26053 8925 26065 8928
rect 26099 8925 26111 8959
rect 26053 8919 26111 8925
rect 20349 8891 20407 8897
rect 20349 8888 20361 8891
rect 19352 8860 20361 8888
rect 18012 8848 18018 8860
rect 20349 8857 20361 8860
rect 20395 8888 20407 8891
rect 20714 8888 20720 8900
rect 20395 8860 20720 8888
rect 20395 8857 20407 8860
rect 20349 8851 20407 8857
rect 20714 8848 20720 8860
rect 20772 8848 20778 8900
rect 22364 8891 22422 8897
rect 22364 8857 22376 8891
rect 22410 8888 22422 8891
rect 24118 8888 24124 8900
rect 22410 8860 24124 8888
rect 22410 8857 22422 8860
rect 22364 8851 22422 8857
rect 24118 8848 24124 8860
rect 24176 8848 24182 8900
rect 24394 8888 24400 8900
rect 24355 8860 24400 8888
rect 24394 8848 24400 8860
rect 24452 8848 24458 8900
rect 24581 8891 24639 8897
rect 24581 8857 24593 8891
rect 24627 8857 24639 8891
rect 24581 8851 24639 8857
rect 25409 8891 25467 8897
rect 25409 8857 25421 8891
rect 25455 8888 25467 8891
rect 25590 8888 25596 8900
rect 25455 8860 25596 8888
rect 25455 8857 25467 8860
rect 25409 8851 25467 8857
rect 19886 8820 19892 8832
rect 17880 8792 19892 8820
rect 19886 8780 19892 8792
rect 19944 8780 19950 8832
rect 19981 8823 20039 8829
rect 19981 8789 19993 8823
rect 20027 8820 20039 8823
rect 20438 8820 20444 8832
rect 20027 8792 20444 8820
rect 20027 8789 20039 8792
rect 19981 8783 20039 8789
rect 20438 8780 20444 8792
rect 20496 8780 20502 8832
rect 23198 8780 23204 8832
rect 23256 8820 23262 8832
rect 23477 8823 23535 8829
rect 23477 8820 23489 8823
rect 23256 8792 23489 8820
rect 23256 8780 23262 8792
rect 23477 8789 23489 8792
rect 23523 8820 23535 8823
rect 24596 8820 24624 8851
rect 25590 8848 25596 8860
rect 25648 8848 25654 8900
rect 26160 8888 26188 8996
rect 33318 8984 33324 8996
rect 33376 8984 33382 9036
rect 34790 8984 34796 9036
rect 34848 9024 34854 9036
rect 35345 9027 35403 9033
rect 35345 9024 35357 9027
rect 34848 8996 35357 9024
rect 34848 8984 34854 8996
rect 35345 8993 35357 8996
rect 35391 9024 35403 9027
rect 35710 9024 35716 9036
rect 35391 8996 35716 9024
rect 35391 8993 35403 8996
rect 35345 8987 35403 8993
rect 35710 8984 35716 8996
rect 35768 8984 35774 9036
rect 37090 9024 37096 9036
rect 36832 8996 37096 9024
rect 26320 8959 26378 8965
rect 26320 8925 26332 8959
rect 26366 8956 26378 8959
rect 26786 8956 26792 8968
rect 26366 8928 26792 8956
rect 26366 8925 26378 8928
rect 26320 8919 26378 8925
rect 26786 8916 26792 8928
rect 26844 8916 26850 8968
rect 30377 8959 30435 8965
rect 30377 8956 30389 8959
rect 27586 8928 30389 8956
rect 27586 8888 27614 8928
rect 30377 8925 30389 8928
rect 30423 8956 30435 8959
rect 31018 8956 31024 8968
rect 30423 8928 31024 8956
rect 30423 8925 30435 8928
rect 30377 8919 30435 8925
rect 31018 8916 31024 8928
rect 31076 8916 31082 8968
rect 31110 8916 31116 8968
rect 31168 8956 31174 8968
rect 31168 8928 31340 8956
rect 31168 8916 31174 8928
rect 31202 8888 31208 8900
rect 26160 8860 27614 8888
rect 31163 8860 31208 8888
rect 31202 8848 31208 8860
rect 31260 8848 31266 8900
rect 31312 8888 31340 8928
rect 31386 8916 31392 8968
rect 31444 8956 31450 8968
rect 33505 8959 33563 8965
rect 31444 8928 31489 8956
rect 31444 8916 31450 8928
rect 33505 8925 33517 8959
rect 33551 8956 33563 8959
rect 34606 8956 34612 8968
rect 33551 8928 34612 8956
rect 33551 8925 33563 8928
rect 33505 8919 33563 8925
rect 34606 8916 34612 8928
rect 34664 8956 34670 8968
rect 35434 8956 35440 8968
rect 34664 8928 35440 8956
rect 34664 8916 34670 8928
rect 35434 8916 35440 8928
rect 35492 8916 35498 8968
rect 35618 8956 35624 8968
rect 35579 8928 35624 8956
rect 35618 8916 35624 8928
rect 35676 8916 35682 8968
rect 36832 8965 36860 8996
rect 37090 8984 37096 8996
rect 37148 8984 37154 9036
rect 37200 8996 38700 9024
rect 36817 8959 36875 8965
rect 36817 8925 36829 8959
rect 36863 8925 36875 8959
rect 36998 8956 37004 8968
rect 36959 8928 37004 8956
rect 36817 8919 36875 8925
rect 36998 8916 37004 8928
rect 37056 8916 37062 8968
rect 37200 8965 37228 8996
rect 37185 8959 37243 8965
rect 37185 8925 37197 8959
rect 37231 8925 37243 8959
rect 37185 8919 37243 8925
rect 37274 8916 37280 8968
rect 37332 8956 37338 8968
rect 37645 8959 37703 8965
rect 37645 8956 37657 8959
rect 37332 8928 37657 8956
rect 37332 8916 37338 8928
rect 37645 8925 37657 8928
rect 37691 8925 37703 8959
rect 37826 8956 37832 8968
rect 37787 8928 37832 8956
rect 37645 8919 37703 8925
rect 37826 8916 37832 8928
rect 37884 8916 37890 8968
rect 33321 8891 33379 8897
rect 33321 8888 33333 8891
rect 31312 8860 33333 8888
rect 33321 8857 33333 8860
rect 33367 8857 33379 8891
rect 33321 8851 33379 8857
rect 36909 8891 36967 8897
rect 36909 8857 36921 8891
rect 36955 8857 36967 8891
rect 36909 8851 36967 8857
rect 38473 8891 38531 8897
rect 38473 8857 38485 8891
rect 38519 8888 38531 8891
rect 38562 8888 38568 8900
rect 38519 8860 38568 8888
rect 38519 8857 38531 8860
rect 38473 8851 38531 8857
rect 23523 8792 24624 8820
rect 31220 8820 31248 8848
rect 31849 8823 31907 8829
rect 31849 8820 31861 8823
rect 31220 8792 31861 8820
rect 23523 8789 23535 8792
rect 23477 8783 23535 8789
rect 31849 8789 31861 8792
rect 31895 8820 31907 8823
rect 32490 8820 32496 8832
rect 31895 8792 32496 8820
rect 31895 8789 31907 8792
rect 31849 8783 31907 8789
rect 32490 8780 32496 8792
rect 32548 8820 32554 8832
rect 33965 8823 34023 8829
rect 33965 8820 33977 8823
rect 32548 8792 33977 8820
rect 32548 8780 32554 8792
rect 33965 8789 33977 8792
rect 34011 8820 34023 8823
rect 34514 8820 34520 8832
rect 34011 8792 34520 8820
rect 34011 8789 34023 8792
rect 33965 8783 34023 8789
rect 34514 8780 34520 8792
rect 34572 8820 34578 8832
rect 34793 8823 34851 8829
rect 34793 8820 34805 8823
rect 34572 8792 34805 8820
rect 34572 8780 34578 8792
rect 34793 8789 34805 8792
rect 34839 8789 34851 8823
rect 36924 8820 36952 8851
rect 38562 8848 38568 8860
rect 38620 8848 38626 8900
rect 38672 8897 38700 8996
rect 68094 8956 68100 8968
rect 68055 8928 68100 8956
rect 68094 8916 68100 8928
rect 68152 8916 68158 8968
rect 38657 8891 38715 8897
rect 38657 8857 38669 8891
rect 38703 8888 38715 8891
rect 41230 8888 41236 8900
rect 38703 8860 41236 8888
rect 38703 8857 38715 8860
rect 38657 8851 38715 8857
rect 41230 8848 41236 8860
rect 41288 8848 41294 8900
rect 37458 8820 37464 8832
rect 36924 8792 37464 8820
rect 34793 8783 34851 8789
rect 37458 8780 37464 8792
rect 37516 8780 37522 8832
rect 38838 8820 38844 8832
rect 38799 8792 38844 8820
rect 38838 8780 38844 8792
rect 38896 8780 38902 8832
rect 1104 8730 68816 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 68816 8730
rect 1104 8656 68816 8678
rect 1581 8619 1639 8625
rect 1581 8585 1593 8619
rect 1627 8616 1639 8619
rect 3142 8616 3148 8628
rect 1627 8588 3148 8616
rect 1627 8585 1639 8588
rect 1581 8579 1639 8585
rect 3142 8576 3148 8588
rect 3200 8576 3206 8628
rect 3970 8616 3976 8628
rect 3931 8588 3976 8616
rect 3970 8576 3976 8588
rect 4028 8576 4034 8628
rect 6457 8619 6515 8625
rect 6457 8585 6469 8619
rect 6503 8616 6515 8619
rect 6730 8616 6736 8628
rect 6503 8588 6736 8616
rect 6503 8585 6515 8588
rect 6457 8579 6515 8585
rect 6730 8576 6736 8588
rect 6788 8576 6794 8628
rect 7374 8616 7380 8628
rect 6840 8588 7380 8616
rect 2682 8508 2688 8560
rect 2740 8548 2746 8560
rect 2838 8551 2896 8557
rect 2838 8548 2850 8551
rect 2740 8520 2850 8548
rect 2740 8508 2746 8520
rect 2838 8517 2850 8520
rect 2884 8517 2896 8551
rect 5718 8548 5724 8560
rect 5631 8520 5724 8548
rect 2838 8511 2896 8517
rect 5718 8508 5724 8520
rect 5776 8548 5782 8560
rect 6840 8548 6868 8588
rect 7374 8576 7380 8588
rect 7432 8576 7438 8628
rect 7469 8619 7527 8625
rect 7469 8585 7481 8619
rect 7515 8616 7527 8619
rect 12434 8616 12440 8628
rect 7515 8588 12440 8616
rect 7515 8585 7527 8588
rect 7469 8579 7527 8585
rect 12434 8576 12440 8588
rect 12492 8576 12498 8628
rect 14274 8576 14280 8628
rect 14332 8616 14338 8628
rect 19518 8616 19524 8628
rect 14332 8588 19524 8616
rect 14332 8576 14338 8588
rect 19518 8576 19524 8588
rect 19576 8576 19582 8628
rect 20070 8576 20076 8628
rect 20128 8616 20134 8628
rect 20128 8588 20199 8616
rect 20128 8576 20134 8588
rect 7101 8551 7159 8557
rect 7101 8548 7113 8551
rect 5776 8520 6868 8548
rect 6932 8520 7113 8548
rect 5776 8508 5782 8520
rect 2038 8440 2044 8492
rect 2096 8480 2102 8492
rect 2133 8483 2191 8489
rect 2133 8480 2145 8483
rect 2096 8452 2145 8480
rect 2096 8440 2102 8452
rect 2133 8449 2145 8452
rect 2179 8480 2191 8483
rect 3878 8480 3884 8492
rect 2179 8452 3884 8480
rect 2179 8449 2191 8452
rect 2133 8443 2191 8449
rect 3878 8440 3884 8452
rect 3936 8440 3942 8492
rect 4798 8480 4804 8492
rect 4759 8452 4804 8480
rect 4798 8440 4804 8452
rect 4856 8440 4862 8492
rect 2593 8415 2651 8421
rect 2593 8381 2605 8415
rect 2639 8381 2651 8415
rect 2593 8375 2651 8381
rect 2608 8276 2636 8375
rect 3970 8372 3976 8424
rect 4028 8412 4034 8424
rect 6932 8412 6960 8520
rect 7101 8517 7113 8520
rect 7147 8517 7159 8551
rect 8389 8551 8447 8557
rect 7101 8511 7159 8517
rect 7300 8520 8248 8548
rect 7300 8489 7328 8520
rect 8220 8492 8248 8520
rect 8389 8517 8401 8551
rect 8435 8548 8447 8551
rect 10410 8548 10416 8560
rect 8435 8520 10416 8548
rect 8435 8517 8447 8520
rect 8389 8511 8447 8517
rect 10410 8508 10416 8520
rect 10468 8508 10474 8560
rect 11146 8548 11152 8560
rect 10704 8520 11152 8548
rect 7009 8483 7067 8489
rect 7009 8449 7021 8483
rect 7055 8449 7067 8483
rect 7009 8443 7067 8449
rect 7285 8483 7343 8489
rect 7285 8449 7297 8483
rect 7331 8449 7343 8483
rect 7285 8443 7343 8449
rect 4028 8384 6960 8412
rect 7024 8412 7052 8443
rect 7650 8440 7656 8492
rect 7708 8480 7714 8492
rect 7929 8483 7987 8489
rect 7929 8480 7941 8483
rect 7708 8452 7941 8480
rect 7708 8440 7714 8452
rect 7929 8449 7941 8452
rect 7975 8449 7987 8483
rect 7929 8443 7987 8449
rect 8021 8483 8079 8489
rect 8021 8449 8033 8483
rect 8067 8449 8079 8483
rect 8202 8480 8208 8492
rect 8163 8452 8208 8480
rect 8021 8443 8079 8449
rect 7668 8412 7696 8440
rect 7024 8384 7696 8412
rect 4028 8372 4034 8384
rect 7834 8372 7840 8424
rect 7892 8412 7898 8424
rect 8036 8412 8064 8443
rect 8202 8440 8208 8452
rect 8260 8440 8266 8492
rect 9677 8483 9735 8489
rect 9677 8449 9689 8483
rect 9723 8480 9735 8483
rect 10137 8483 10195 8489
rect 10137 8480 10149 8483
rect 9723 8452 10149 8480
rect 9723 8449 9735 8452
rect 9677 8443 9735 8449
rect 10137 8449 10149 8452
rect 10183 8480 10195 8483
rect 10704 8480 10732 8520
rect 11146 8508 11152 8520
rect 11204 8508 11210 8560
rect 19426 8548 19432 8560
rect 12360 8520 19432 8548
rect 10183 8452 10732 8480
rect 10965 8483 11023 8489
rect 10183 8449 10195 8452
rect 10137 8443 10195 8449
rect 10965 8449 10977 8483
rect 11011 8480 11023 8483
rect 12066 8480 12072 8492
rect 11011 8452 11468 8480
rect 12027 8452 12072 8480
rect 11011 8449 11023 8452
rect 10965 8443 11023 8449
rect 7892 8384 8064 8412
rect 7892 8372 7898 8384
rect 8662 8372 8668 8424
rect 8720 8412 8726 8424
rect 8849 8415 8907 8421
rect 8849 8412 8861 8415
rect 8720 8384 8861 8412
rect 8720 8372 8726 8384
rect 8849 8381 8861 8384
rect 8895 8381 8907 8415
rect 11238 8412 11244 8424
rect 8849 8375 8907 8381
rect 10336 8384 11244 8412
rect 7742 8304 7748 8356
rect 7800 8344 7806 8356
rect 9674 8344 9680 8356
rect 7800 8316 9680 8344
rect 7800 8304 7806 8316
rect 9674 8304 9680 8316
rect 9732 8304 9738 8356
rect 10336 8353 10364 8384
rect 11238 8372 11244 8384
rect 11296 8372 11302 8424
rect 11440 8356 11468 8452
rect 12066 8440 12072 8452
rect 12124 8440 12130 8492
rect 12158 8440 12164 8492
rect 12216 8480 12222 8492
rect 12360 8489 12388 8520
rect 19426 8508 19432 8520
rect 19484 8508 19490 8560
rect 12253 8483 12311 8489
rect 12253 8480 12265 8483
rect 12216 8452 12265 8480
rect 12216 8440 12222 8452
rect 12253 8449 12265 8452
rect 12299 8449 12311 8483
rect 12253 8443 12311 8449
rect 12345 8483 12403 8489
rect 12345 8449 12357 8483
rect 12391 8449 12403 8483
rect 12345 8443 12403 8449
rect 12526 8440 12532 8492
rect 12584 8480 12590 8492
rect 12621 8483 12679 8489
rect 12621 8480 12633 8483
rect 12584 8452 12633 8480
rect 12584 8440 12590 8452
rect 12621 8449 12633 8452
rect 12667 8449 12679 8483
rect 12621 8443 12679 8449
rect 13909 8483 13967 8489
rect 13909 8449 13921 8483
rect 13955 8480 13967 8483
rect 16390 8480 16396 8492
rect 13955 8452 16396 8480
rect 13955 8449 13967 8452
rect 13909 8443 13967 8449
rect 16390 8440 16396 8452
rect 16448 8440 16454 8492
rect 18046 8440 18052 8492
rect 18104 8480 18110 8492
rect 18610 8483 18668 8489
rect 18610 8480 18622 8483
rect 18104 8452 18622 8480
rect 18104 8440 18110 8452
rect 18610 8449 18622 8452
rect 18656 8449 18668 8483
rect 18610 8443 18668 8449
rect 19610 8440 19616 8492
rect 19668 8480 19674 8492
rect 19889 8483 19947 8489
rect 19889 8480 19901 8483
rect 19668 8452 19901 8480
rect 19668 8440 19674 8452
rect 19889 8449 19901 8452
rect 19935 8449 19947 8483
rect 19889 8443 19947 8449
rect 20073 8486 20131 8492
rect 20171 8489 20199 8588
rect 20254 8576 20260 8628
rect 20312 8576 20318 8628
rect 23477 8619 23535 8625
rect 23477 8585 23489 8619
rect 23523 8616 23535 8619
rect 23658 8616 23664 8628
rect 23523 8588 23664 8616
rect 23523 8585 23535 8588
rect 23477 8579 23535 8585
rect 23658 8576 23664 8588
rect 23716 8576 23722 8628
rect 24302 8576 24308 8628
rect 24360 8616 24366 8628
rect 28626 8616 28632 8628
rect 24360 8588 28632 8616
rect 24360 8576 24366 8588
rect 28626 8576 28632 8588
rect 28684 8576 28690 8628
rect 28810 8616 28816 8628
rect 28771 8588 28816 8616
rect 28810 8576 28816 8588
rect 28868 8576 28874 8628
rect 32122 8616 32128 8628
rect 32083 8588 32128 8616
rect 32122 8576 32128 8588
rect 32180 8576 32186 8628
rect 32324 8588 33456 8616
rect 20272 8489 20300 8576
rect 20533 8551 20591 8557
rect 20533 8517 20545 8551
rect 20579 8548 20591 8551
rect 20806 8548 20812 8560
rect 20579 8520 20812 8548
rect 20579 8517 20591 8520
rect 20533 8511 20591 8517
rect 20806 8508 20812 8520
rect 20864 8508 20870 8560
rect 23198 8548 23204 8560
rect 23159 8520 23204 8548
rect 23198 8508 23204 8520
rect 23256 8508 23262 8560
rect 24854 8508 24860 8560
rect 24912 8508 24918 8560
rect 27798 8508 27804 8560
rect 27856 8548 27862 8560
rect 28445 8551 28503 8557
rect 28445 8548 28457 8551
rect 27856 8520 28457 8548
rect 27856 8508 27862 8520
rect 28445 8517 28457 8520
rect 28491 8517 28503 8551
rect 28445 8511 28503 8517
rect 28537 8551 28595 8557
rect 28537 8517 28549 8551
rect 28583 8548 28595 8551
rect 28583 8520 29500 8548
rect 28583 8517 28595 8520
rect 28537 8511 28595 8517
rect 20073 8452 20085 8486
rect 20119 8452 20131 8486
rect 20073 8446 20131 8452
rect 20165 8483 20223 8489
rect 20165 8449 20177 8483
rect 20211 8449 20223 8483
rect 11974 8372 11980 8424
rect 12032 8412 12038 8424
rect 12437 8415 12495 8421
rect 12437 8412 12449 8415
rect 12032 8384 12449 8412
rect 12032 8372 12038 8384
rect 12437 8381 12449 8384
rect 12483 8381 12495 8415
rect 13630 8412 13636 8424
rect 13591 8384 13636 8412
rect 12437 8375 12495 8381
rect 13630 8372 13636 8384
rect 13688 8372 13694 8424
rect 15286 8372 15292 8424
rect 15344 8412 15350 8424
rect 15381 8415 15439 8421
rect 15381 8412 15393 8415
rect 15344 8384 15393 8412
rect 15344 8372 15350 8384
rect 15381 8381 15393 8384
rect 15427 8381 15439 8415
rect 15381 8375 15439 8381
rect 15838 8372 15844 8424
rect 15896 8412 15902 8424
rect 16025 8415 16083 8421
rect 16025 8412 16037 8415
rect 15896 8384 16037 8412
rect 15896 8372 15902 8384
rect 16025 8381 16037 8384
rect 16071 8381 16083 8415
rect 16025 8375 16083 8381
rect 18877 8415 18935 8421
rect 18877 8381 18889 8415
rect 18923 8412 18935 8415
rect 20091 8412 20119 8446
rect 20165 8443 20223 8449
rect 20257 8483 20315 8489
rect 20257 8449 20269 8483
rect 20303 8449 20315 8483
rect 20257 8443 20315 8449
rect 21910 8440 21916 8492
rect 21968 8480 21974 8492
rect 22925 8483 22983 8489
rect 22925 8480 22937 8483
rect 21968 8452 22937 8480
rect 21968 8440 21974 8452
rect 22925 8449 22937 8452
rect 22971 8449 22983 8483
rect 23106 8480 23112 8492
rect 23067 8452 23112 8480
rect 22925 8443 22983 8449
rect 23106 8440 23112 8452
rect 23164 8440 23170 8492
rect 23293 8483 23351 8489
rect 23293 8449 23305 8483
rect 23339 8480 23351 8483
rect 23566 8480 23572 8492
rect 23339 8452 23572 8480
rect 23339 8449 23351 8452
rect 23293 8443 23351 8449
rect 23566 8440 23572 8452
rect 23624 8440 23630 8492
rect 24872 8480 24900 8508
rect 29472 8492 29500 8520
rect 31018 8508 31024 8560
rect 31076 8548 31082 8560
rect 31573 8551 31631 8557
rect 31573 8548 31585 8551
rect 31076 8520 31585 8548
rect 31076 8508 31082 8520
rect 31573 8517 31585 8520
rect 31619 8548 31631 8551
rect 32324 8548 32352 8588
rect 32490 8548 32496 8560
rect 31619 8520 32352 8548
rect 32451 8520 32496 8548
rect 31619 8517 31631 8520
rect 31573 8511 31631 8517
rect 25133 8483 25191 8489
rect 25133 8480 25145 8483
rect 24872 8452 25145 8480
rect 25133 8449 25145 8452
rect 25179 8449 25191 8483
rect 26142 8480 26148 8492
rect 26103 8452 26148 8480
rect 25133 8443 25191 8449
rect 26142 8440 26148 8452
rect 26200 8440 26206 8492
rect 27154 8440 27160 8492
rect 27212 8480 27218 8492
rect 28261 8483 28319 8489
rect 28261 8480 28273 8483
rect 27212 8452 28273 8480
rect 27212 8440 27218 8452
rect 28261 8449 28273 8452
rect 28307 8449 28319 8483
rect 28626 8480 28632 8492
rect 28261 8443 28319 8449
rect 28368 8452 28632 8480
rect 20438 8412 20444 8424
rect 18923 8384 20024 8412
rect 20091 8384 20444 8412
rect 18923 8381 18935 8384
rect 18877 8375 18935 8381
rect 19996 8356 20024 8384
rect 20438 8372 20444 8384
rect 20496 8372 20502 8424
rect 24857 8415 24915 8421
rect 24857 8381 24869 8415
rect 24903 8412 24915 8415
rect 25038 8412 25044 8424
rect 24903 8384 25044 8412
rect 24903 8381 24915 8384
rect 24857 8375 24915 8381
rect 25038 8372 25044 8384
rect 25096 8372 25102 8424
rect 26421 8415 26479 8421
rect 26421 8381 26433 8415
rect 26467 8412 26479 8415
rect 26694 8412 26700 8424
rect 26467 8384 26700 8412
rect 26467 8381 26479 8384
rect 26421 8375 26479 8381
rect 10321 8347 10379 8353
rect 10321 8313 10333 8347
rect 10367 8313 10379 8347
rect 10778 8344 10784 8356
rect 10739 8316 10784 8344
rect 10321 8307 10379 8313
rect 10778 8304 10784 8316
rect 10836 8304 10842 8356
rect 11422 8304 11428 8356
rect 11480 8344 11486 8356
rect 11517 8347 11575 8353
rect 11517 8344 11529 8347
rect 11480 8316 11529 8344
rect 11480 8304 11486 8316
rect 11517 8313 11529 8316
rect 11563 8313 11575 8347
rect 11517 8307 11575 8313
rect 11882 8304 11888 8356
rect 11940 8344 11946 8356
rect 12250 8344 12256 8356
rect 11940 8316 12256 8344
rect 11940 8304 11946 8316
rect 12250 8304 12256 8316
rect 12308 8344 12314 8356
rect 16853 8347 16911 8353
rect 16853 8344 16865 8347
rect 12308 8316 12388 8344
rect 12308 8304 12314 8316
rect 2958 8276 2964 8288
rect 2608 8248 2964 8276
rect 2958 8236 2964 8248
rect 3016 8236 3022 8288
rect 4985 8279 5043 8285
rect 4985 8245 4997 8279
rect 5031 8276 5043 8279
rect 5074 8276 5080 8288
rect 5031 8248 5080 8276
rect 5031 8245 5043 8248
rect 4985 8239 5043 8245
rect 5074 8236 5080 8248
rect 5132 8236 5138 8288
rect 12360 8276 12388 8316
rect 12452 8316 16865 8344
rect 12452 8276 12480 8316
rect 16853 8313 16865 8316
rect 16899 8344 16911 8347
rect 17034 8344 17040 8356
rect 16899 8316 17040 8344
rect 16899 8313 16911 8316
rect 16853 8307 16911 8313
rect 17034 8304 17040 8316
rect 17092 8304 17098 8356
rect 17218 8304 17224 8356
rect 17276 8344 17282 8356
rect 17276 8316 18000 8344
rect 17276 8304 17282 8316
rect 12802 8276 12808 8288
rect 12360 8248 12480 8276
rect 12763 8248 12808 8276
rect 12802 8236 12808 8248
rect 12860 8236 12866 8288
rect 13354 8236 13360 8288
rect 13412 8276 13418 8288
rect 16206 8276 16212 8288
rect 13412 8248 16212 8276
rect 13412 8236 13418 8248
rect 16206 8236 16212 8248
rect 16264 8236 16270 8288
rect 17402 8236 17408 8288
rect 17460 8276 17466 8288
rect 17497 8279 17555 8285
rect 17497 8276 17509 8279
rect 17460 8248 17509 8276
rect 17460 8236 17466 8248
rect 17497 8245 17509 8248
rect 17543 8245 17555 8279
rect 17972 8276 18000 8316
rect 18892 8316 19932 8344
rect 18892 8276 18920 8316
rect 17972 8248 18920 8276
rect 17497 8239 17555 8245
rect 19334 8236 19340 8288
rect 19392 8276 19398 8288
rect 19904 8276 19932 8316
rect 19978 8304 19984 8356
rect 20036 8344 20042 8356
rect 20530 8344 20536 8356
rect 20036 8316 20536 8344
rect 20036 8304 20042 8316
rect 20530 8304 20536 8316
rect 20588 8304 20594 8356
rect 23566 8304 23572 8356
rect 23624 8344 23630 8356
rect 26436 8344 26464 8375
rect 26694 8372 26700 8384
rect 26752 8412 26758 8424
rect 26973 8415 27031 8421
rect 26973 8412 26985 8415
rect 26752 8384 26985 8412
rect 26752 8372 26758 8384
rect 26973 8381 26985 8384
rect 27019 8381 27031 8415
rect 26973 8375 27031 8381
rect 27249 8415 27307 8421
rect 27249 8381 27261 8415
rect 27295 8412 27307 8415
rect 27706 8412 27712 8424
rect 27295 8384 27712 8412
rect 27295 8381 27307 8384
rect 27249 8375 27307 8381
rect 27706 8372 27712 8384
rect 27764 8412 27770 8424
rect 28368 8412 28396 8452
rect 28626 8440 28632 8452
rect 28684 8440 28690 8492
rect 29270 8480 29276 8492
rect 29231 8452 29276 8480
rect 29270 8440 29276 8452
rect 29328 8440 29334 8492
rect 29454 8480 29460 8492
rect 29415 8452 29460 8480
rect 29454 8440 29460 8452
rect 29512 8440 29518 8492
rect 32324 8489 32352 8520
rect 32490 8508 32496 8520
rect 32548 8508 32554 8560
rect 32309 8483 32367 8489
rect 32309 8449 32321 8483
rect 32355 8449 32367 8483
rect 32309 8443 32367 8449
rect 32398 8440 32404 8492
rect 32456 8480 32462 8492
rect 32456 8452 32501 8480
rect 32456 8440 32462 8452
rect 32582 8440 32588 8492
rect 32640 8480 32646 8492
rect 33428 8489 33456 8588
rect 39022 8576 39028 8628
rect 39080 8616 39086 8628
rect 39850 8616 39856 8628
rect 39080 8588 39856 8616
rect 39080 8576 39086 8588
rect 39850 8576 39856 8588
rect 39908 8616 39914 8628
rect 40037 8619 40095 8625
rect 40037 8616 40049 8619
rect 39908 8588 40049 8616
rect 39908 8576 39914 8588
rect 40037 8585 40049 8588
rect 40083 8585 40095 8619
rect 40037 8579 40095 8585
rect 34149 8551 34207 8557
rect 34149 8517 34161 8551
rect 34195 8548 34207 8551
rect 34790 8548 34796 8560
rect 34195 8520 34796 8548
rect 34195 8517 34207 8520
rect 34149 8511 34207 8517
rect 34790 8508 34796 8520
rect 34848 8508 34854 8560
rect 38746 8548 38752 8560
rect 38707 8520 38752 8548
rect 38746 8508 38752 8520
rect 38804 8508 38810 8560
rect 32677 8483 32735 8489
rect 32677 8480 32689 8483
rect 32640 8452 32689 8480
rect 32640 8440 32646 8452
rect 32677 8449 32689 8452
rect 32723 8449 32735 8483
rect 32677 8443 32735 8449
rect 33413 8483 33471 8489
rect 33413 8449 33425 8483
rect 33459 8480 33471 8483
rect 34054 8480 34060 8492
rect 33459 8452 34060 8480
rect 33459 8449 33471 8452
rect 33413 8443 33471 8449
rect 34054 8440 34060 8452
rect 34112 8440 34118 8492
rect 34241 8483 34299 8489
rect 34241 8449 34253 8483
rect 34287 8449 34299 8483
rect 34422 8480 34428 8492
rect 34383 8452 34428 8480
rect 34241 8443 34299 8449
rect 27764 8384 28396 8412
rect 27764 8372 27770 8384
rect 28718 8372 28724 8424
rect 28776 8412 28782 8424
rect 34256 8412 34284 8443
rect 34422 8440 34428 8452
rect 34480 8440 34486 8492
rect 34698 8440 34704 8492
rect 34756 8480 34762 8492
rect 34885 8483 34943 8489
rect 34885 8480 34897 8483
rect 34756 8452 34897 8480
rect 34756 8440 34762 8452
rect 34885 8449 34897 8452
rect 34931 8449 34943 8483
rect 35710 8480 35716 8492
rect 35671 8452 35716 8480
rect 34885 8443 34943 8449
rect 35710 8440 35716 8452
rect 35768 8440 35774 8492
rect 37090 8440 37096 8492
rect 37148 8480 37154 8492
rect 37553 8483 37611 8489
rect 37553 8480 37565 8483
rect 37148 8452 37565 8480
rect 37148 8440 37154 8452
rect 37553 8449 37565 8452
rect 37599 8449 37611 8483
rect 37553 8443 37611 8449
rect 34514 8412 34520 8424
rect 28776 8384 32720 8412
rect 34256 8384 34520 8412
rect 28776 8372 28782 8384
rect 32692 8356 32720 8384
rect 34514 8372 34520 8384
rect 34572 8372 34578 8424
rect 35986 8412 35992 8424
rect 35947 8384 35992 8412
rect 35986 8372 35992 8384
rect 36044 8372 36050 8424
rect 37274 8412 37280 8424
rect 37235 8384 37280 8412
rect 37274 8372 37280 8384
rect 37332 8372 37338 8424
rect 23624 8316 26464 8344
rect 23624 8304 23630 8316
rect 28166 8304 28172 8356
rect 28224 8344 28230 8356
rect 30469 8347 30527 8353
rect 30469 8344 30481 8347
rect 28224 8316 30481 8344
rect 28224 8304 28230 8316
rect 30469 8313 30481 8316
rect 30515 8344 30527 8347
rect 31202 8344 31208 8356
rect 30515 8316 31208 8344
rect 30515 8313 30527 8316
rect 30469 8307 30527 8313
rect 31202 8304 31208 8316
rect 31260 8304 31266 8356
rect 32674 8304 32680 8356
rect 32732 8304 32738 8356
rect 33870 8344 33876 8356
rect 33831 8316 33876 8344
rect 33870 8304 33876 8316
rect 33928 8304 33934 8356
rect 35069 8347 35127 8353
rect 35069 8313 35081 8347
rect 35115 8344 35127 8347
rect 35894 8344 35900 8356
rect 35115 8316 35900 8344
rect 35115 8313 35127 8316
rect 35069 8307 35127 8313
rect 35894 8304 35900 8316
rect 35952 8344 35958 8356
rect 38562 8344 38568 8356
rect 35952 8316 38568 8344
rect 35952 8304 35958 8316
rect 38562 8304 38568 8316
rect 38620 8304 38626 8356
rect 20898 8276 20904 8288
rect 19392 8248 19437 8276
rect 19904 8248 20904 8276
rect 19392 8236 19398 8248
rect 20898 8236 20904 8248
rect 20956 8236 20962 8288
rect 29641 8279 29699 8285
rect 29641 8245 29653 8279
rect 29687 8276 29699 8279
rect 29730 8276 29736 8288
rect 29687 8248 29736 8276
rect 29687 8245 29699 8248
rect 29641 8239 29699 8245
rect 29730 8236 29736 8248
rect 29788 8236 29794 8288
rect 1104 8186 68816 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 65654 8186
rect 65706 8134 65718 8186
rect 65770 8134 65782 8186
rect 65834 8134 65846 8186
rect 65898 8134 65910 8186
rect 65962 8134 68816 8186
rect 1104 8112 68816 8134
rect 2590 8032 2596 8084
rect 2648 8072 2654 8084
rect 2866 8072 2872 8084
rect 2648 8044 2872 8072
rect 2648 8032 2654 8044
rect 2866 8032 2872 8044
rect 2924 8032 2930 8084
rect 7742 8072 7748 8084
rect 7703 8044 7748 8072
rect 7742 8032 7748 8044
rect 7800 8032 7806 8084
rect 8389 8075 8447 8081
rect 8389 8041 8401 8075
rect 8435 8072 8447 8075
rect 9769 8075 9827 8081
rect 8435 8044 9720 8072
rect 8435 8041 8447 8044
rect 8389 8035 8447 8041
rect 2682 7964 2688 8016
rect 2740 8004 2746 8016
rect 3326 8004 3332 8016
rect 2740 7976 3332 8004
rect 2740 7964 2746 7976
rect 3326 7964 3332 7976
rect 3384 7964 3390 8016
rect 6181 8007 6239 8013
rect 6181 7973 6193 8007
rect 6227 8004 6239 8007
rect 6822 8004 6828 8016
rect 6227 7976 6828 8004
rect 6227 7973 6239 7976
rect 6181 7967 6239 7973
rect 6822 7964 6828 7976
rect 6880 8004 6886 8016
rect 6880 7976 9444 8004
rect 6880 7964 6886 7976
rect 2314 7936 2320 7948
rect 2275 7908 2320 7936
rect 2314 7896 2320 7908
rect 2372 7896 2378 7948
rect 2041 7871 2099 7877
rect 2041 7837 2053 7871
rect 2087 7868 2099 7871
rect 2590 7868 2596 7880
rect 2087 7840 2596 7868
rect 2087 7837 2099 7840
rect 2041 7831 2099 7837
rect 2590 7828 2596 7840
rect 2648 7828 2654 7880
rect 4614 7828 4620 7880
rect 4672 7868 4678 7880
rect 5074 7877 5080 7880
rect 4801 7871 4859 7877
rect 4801 7868 4813 7871
rect 4672 7840 4813 7868
rect 4672 7828 4678 7840
rect 4801 7837 4813 7840
rect 4847 7837 4859 7871
rect 5068 7868 5080 7877
rect 5035 7840 5080 7868
rect 4801 7831 4859 7837
rect 5068 7831 5080 7840
rect 5074 7828 5080 7831
rect 5132 7828 5138 7880
rect 7285 7871 7343 7877
rect 7285 7837 7297 7871
rect 7331 7868 7343 7871
rect 7561 7871 7619 7877
rect 7331 7840 7512 7868
rect 7331 7837 7343 7840
rect 7285 7831 7343 7837
rect 2133 7803 2191 7809
rect 2133 7769 2145 7803
rect 2179 7800 2191 7803
rect 4430 7800 4436 7812
rect 2179 7772 4436 7800
rect 2179 7769 2191 7772
rect 2133 7763 2191 7769
rect 4430 7760 4436 7772
rect 4488 7800 4494 7812
rect 7377 7803 7435 7809
rect 7377 7800 7389 7803
rect 4488 7772 7389 7800
rect 4488 7760 4494 7772
rect 7377 7769 7389 7772
rect 7423 7769 7435 7803
rect 7484 7800 7512 7840
rect 7561 7837 7573 7871
rect 7607 7868 7619 7871
rect 8202 7868 8208 7880
rect 7607 7840 8208 7868
rect 7607 7837 7619 7840
rect 7561 7831 7619 7837
rect 8202 7828 8208 7840
rect 8260 7828 8266 7880
rect 9416 7877 9444 7976
rect 9692 7936 9720 8044
rect 9769 8041 9781 8075
rect 9815 8072 9827 8075
rect 12158 8072 12164 8084
rect 9815 8044 12164 8072
rect 9815 8041 9827 8044
rect 9769 8035 9827 8041
rect 12158 8032 12164 8044
rect 12216 8032 12222 8084
rect 17494 8072 17500 8084
rect 17052 8044 17500 8072
rect 11701 8007 11759 8013
rect 11701 7973 11713 8007
rect 11747 8004 11759 8007
rect 12526 8004 12532 8016
rect 11747 7976 12532 8004
rect 11747 7973 11759 7976
rect 11701 7967 11759 7973
rect 12526 7964 12532 7976
rect 12584 7964 12590 8016
rect 12158 7936 12164 7948
rect 9692 7908 12164 7936
rect 12158 7896 12164 7908
rect 12216 7896 12222 7948
rect 9309 7871 9367 7877
rect 9309 7837 9321 7871
rect 9355 7837 9367 7871
rect 9309 7831 9367 7837
rect 9401 7871 9459 7877
rect 9401 7837 9413 7871
rect 9447 7837 9459 7871
rect 9401 7831 9459 7837
rect 7650 7800 7656 7812
rect 7484 7772 7656 7800
rect 7377 7763 7435 7769
rect 7650 7760 7656 7772
rect 7708 7760 7714 7812
rect 9324 7800 9352 7831
rect 9490 7828 9496 7880
rect 9548 7868 9554 7880
rect 9585 7871 9643 7877
rect 9585 7868 9597 7871
rect 9548 7840 9597 7868
rect 9548 7828 9554 7840
rect 9585 7837 9597 7840
rect 9631 7868 9643 7871
rect 10321 7871 10379 7877
rect 10321 7868 10333 7871
rect 9631 7840 10333 7868
rect 9631 7837 9643 7840
rect 9585 7831 9643 7837
rect 10321 7837 10333 7840
rect 10367 7837 10379 7871
rect 10321 7831 10379 7837
rect 11517 7871 11575 7877
rect 11517 7837 11529 7871
rect 11563 7868 11575 7871
rect 11790 7868 11796 7880
rect 11563 7840 11796 7868
rect 11563 7837 11575 7840
rect 11517 7831 11575 7837
rect 11790 7828 11796 7840
rect 11848 7828 11854 7880
rect 12802 7828 12808 7880
rect 12860 7868 12866 7880
rect 13274 7871 13332 7877
rect 13274 7868 13286 7871
rect 12860 7840 13286 7868
rect 12860 7828 12866 7840
rect 13274 7837 13286 7840
rect 13320 7837 13332 7871
rect 13274 7831 13332 7837
rect 13446 7828 13452 7880
rect 13504 7868 13510 7880
rect 13541 7871 13599 7877
rect 13541 7868 13553 7871
rect 13504 7840 13553 7868
rect 13504 7828 13510 7840
rect 13541 7837 13553 7840
rect 13587 7868 13599 7871
rect 15933 7871 15991 7877
rect 15933 7868 15945 7871
rect 13587 7840 15945 7868
rect 13587 7837 13599 7840
rect 13541 7831 13599 7837
rect 15933 7837 15945 7840
rect 15979 7868 15991 7871
rect 16298 7868 16304 7880
rect 15979 7840 16304 7868
rect 15979 7837 15991 7840
rect 15933 7831 15991 7837
rect 16298 7828 16304 7840
rect 16356 7828 16362 7880
rect 16390 7828 16396 7880
rect 16448 7868 16454 7880
rect 17052 7877 17080 8044
rect 17494 8032 17500 8044
rect 17552 8032 17558 8084
rect 17589 8075 17647 8081
rect 17589 8041 17601 8075
rect 17635 8072 17647 8075
rect 18046 8072 18052 8084
rect 17635 8044 18052 8072
rect 17635 8041 17647 8044
rect 17589 8035 17647 8041
rect 18046 8032 18052 8044
rect 18104 8032 18110 8084
rect 21910 8072 21916 8084
rect 21871 8044 21916 8072
rect 21910 8032 21916 8044
rect 21968 8032 21974 8084
rect 23750 8072 23756 8084
rect 23711 8044 23756 8072
rect 23750 8032 23756 8044
rect 23808 8032 23814 8084
rect 26881 8075 26939 8081
rect 26881 8041 26893 8075
rect 26927 8072 26939 8075
rect 27062 8072 27068 8084
rect 26927 8044 27068 8072
rect 26927 8041 26939 8044
rect 26881 8035 26939 8041
rect 27062 8032 27068 8044
rect 27120 8032 27126 8084
rect 28997 8075 29055 8081
rect 28997 8072 29009 8075
rect 27586 8044 29009 8072
rect 17862 8004 17868 8016
rect 17144 7976 17868 8004
rect 17144 7945 17172 7976
rect 17862 7964 17868 7976
rect 17920 7964 17926 8016
rect 25590 7964 25596 8016
rect 25648 7964 25654 8016
rect 26050 7964 26056 8016
rect 26108 8004 26114 8016
rect 27586 8004 27614 8044
rect 28997 8041 29009 8044
rect 29043 8072 29055 8075
rect 29043 8044 34376 8072
rect 29043 8041 29055 8044
rect 28997 8035 29055 8041
rect 29730 8004 29736 8016
rect 26108 7976 27614 8004
rect 29656 7976 29736 8004
rect 26108 7964 26114 7976
rect 17123 7939 17181 7945
rect 17123 7905 17135 7939
rect 17169 7905 17181 7939
rect 23474 7936 23480 7948
rect 17123 7899 17181 7905
rect 23216 7908 23480 7936
rect 16853 7871 16911 7877
rect 16853 7868 16865 7871
rect 16448 7840 16865 7868
rect 16448 7828 16454 7840
rect 16853 7837 16865 7840
rect 16899 7837 16911 7871
rect 16853 7831 16911 7837
rect 17037 7871 17095 7877
rect 17037 7837 17049 7871
rect 17083 7837 17095 7871
rect 17037 7831 17095 7837
rect 17221 7871 17279 7877
rect 17221 7837 17233 7871
rect 17267 7837 17279 7871
rect 17402 7868 17408 7880
rect 17363 7840 17408 7868
rect 17221 7831 17279 7837
rect 9674 7800 9680 7812
rect 9324 7772 9680 7800
rect 9674 7760 9680 7772
rect 9732 7760 9738 7812
rect 10505 7803 10563 7809
rect 10505 7769 10517 7803
rect 10551 7800 10563 7803
rect 10551 7772 14872 7800
rect 10551 7769 10563 7772
rect 10505 7763 10563 7769
rect 1673 7735 1731 7741
rect 1673 7701 1685 7735
rect 1719 7732 1731 7735
rect 1854 7732 1860 7744
rect 1719 7704 1860 7732
rect 1719 7701 1731 7704
rect 1673 7695 1731 7701
rect 1854 7692 1860 7704
rect 1912 7692 1918 7744
rect 2866 7692 2872 7744
rect 2924 7732 2930 7744
rect 2961 7735 3019 7741
rect 2961 7732 2973 7735
rect 2924 7704 2973 7732
rect 2924 7692 2930 7704
rect 2961 7701 2973 7704
rect 3007 7732 3019 7735
rect 3326 7732 3332 7744
rect 3007 7704 3332 7732
rect 3007 7701 3019 7704
rect 2961 7695 3019 7701
rect 3326 7692 3332 7704
rect 3384 7692 3390 7744
rect 4341 7735 4399 7741
rect 4341 7701 4353 7735
rect 4387 7732 4399 7735
rect 4890 7732 4896 7744
rect 4387 7704 4896 7732
rect 4387 7701 4399 7704
rect 4341 7695 4399 7701
rect 4890 7692 4896 7704
rect 4948 7692 4954 7744
rect 6825 7735 6883 7741
rect 6825 7701 6837 7735
rect 6871 7732 6883 7735
rect 7190 7732 7196 7744
rect 6871 7704 7196 7732
rect 6871 7701 6883 7704
rect 6825 7695 6883 7701
rect 7190 7692 7196 7704
rect 7248 7692 7254 7744
rect 8386 7692 8392 7744
rect 8444 7732 8450 7744
rect 10520 7732 10548 7763
rect 11054 7732 11060 7744
rect 8444 7704 10548 7732
rect 11015 7704 11060 7732
rect 8444 7692 8450 7704
rect 11054 7692 11060 7704
rect 11112 7692 11118 7744
rect 12161 7735 12219 7741
rect 12161 7701 12173 7735
rect 12207 7732 12219 7735
rect 12434 7732 12440 7744
rect 12207 7704 12440 7732
rect 12207 7701 12219 7704
rect 12161 7695 12219 7701
rect 12434 7692 12440 7704
rect 12492 7692 12498 7744
rect 14553 7735 14611 7741
rect 14553 7701 14565 7735
rect 14599 7732 14611 7735
rect 14734 7732 14740 7744
rect 14599 7704 14740 7732
rect 14599 7701 14611 7704
rect 14553 7695 14611 7701
rect 14734 7692 14740 7704
rect 14792 7692 14798 7744
rect 14844 7732 14872 7772
rect 14918 7760 14924 7812
rect 14976 7800 14982 7812
rect 15666 7803 15724 7809
rect 15666 7800 15678 7803
rect 14976 7772 15678 7800
rect 14976 7760 14982 7772
rect 15666 7769 15678 7772
rect 15712 7769 15724 7803
rect 15666 7763 15724 7769
rect 16942 7760 16948 7812
rect 17000 7800 17006 7812
rect 17236 7800 17264 7831
rect 17402 7828 17408 7840
rect 17460 7828 17466 7880
rect 18233 7871 18291 7877
rect 18233 7837 18245 7871
rect 18279 7868 18291 7871
rect 18322 7868 18328 7880
rect 18279 7840 18328 7868
rect 18279 7837 18291 7840
rect 18233 7831 18291 7837
rect 18322 7828 18328 7840
rect 18380 7828 18386 7880
rect 20530 7868 20536 7880
rect 20491 7840 20536 7868
rect 20530 7828 20536 7840
rect 20588 7828 20594 7880
rect 20806 7877 20812 7880
rect 20800 7868 20812 7877
rect 20767 7840 20812 7868
rect 20800 7831 20812 7840
rect 20806 7828 20812 7831
rect 20864 7828 20870 7880
rect 23216 7877 23244 7908
rect 23474 7896 23480 7908
rect 23532 7896 23538 7948
rect 24946 7896 24952 7948
rect 25004 7936 25010 7948
rect 25608 7936 25636 7964
rect 25869 7939 25927 7945
rect 25869 7936 25881 7939
rect 25004 7908 25881 7936
rect 25004 7896 25010 7908
rect 25869 7905 25881 7908
rect 25915 7905 25927 7939
rect 27341 7939 27399 7945
rect 27341 7936 27353 7939
rect 25869 7899 25927 7905
rect 26528 7908 27353 7936
rect 23201 7871 23259 7877
rect 23201 7837 23213 7871
rect 23247 7837 23259 7871
rect 23566 7868 23572 7880
rect 23527 7840 23572 7868
rect 23201 7831 23259 7837
rect 23566 7828 23572 7840
rect 23624 7828 23630 7880
rect 24394 7868 24400 7880
rect 24355 7840 24400 7868
rect 24394 7828 24400 7840
rect 24452 7828 24458 7880
rect 25593 7871 25651 7877
rect 25593 7837 25605 7871
rect 25639 7868 25651 7871
rect 25774 7868 25780 7880
rect 25639 7840 25780 7868
rect 25639 7837 25651 7840
rect 25593 7831 25651 7837
rect 25774 7828 25780 7840
rect 25832 7828 25838 7880
rect 25958 7828 25964 7880
rect 26016 7868 26022 7880
rect 26329 7871 26387 7877
rect 26329 7868 26341 7871
rect 26016 7840 26341 7868
rect 26016 7828 26022 7840
rect 26329 7837 26341 7840
rect 26375 7837 26387 7871
rect 26329 7831 26387 7837
rect 17000 7772 17264 7800
rect 17000 7760 17006 7772
rect 22646 7760 22652 7812
rect 22704 7800 22710 7812
rect 23106 7800 23112 7812
rect 22704 7772 23112 7800
rect 22704 7760 22710 7772
rect 23106 7760 23112 7772
rect 23164 7800 23170 7812
rect 23385 7803 23443 7809
rect 23385 7800 23397 7803
rect 23164 7772 23397 7800
rect 23164 7760 23170 7772
rect 23385 7769 23397 7772
rect 23431 7769 23443 7803
rect 23385 7763 23443 7769
rect 23477 7803 23535 7809
rect 23477 7769 23489 7803
rect 23523 7800 23535 7803
rect 23658 7800 23664 7812
rect 23523 7772 23664 7800
rect 23523 7769 23535 7772
rect 23477 7763 23535 7769
rect 18506 7732 18512 7744
rect 14844 7704 18512 7732
rect 18506 7692 18512 7704
rect 18564 7692 18570 7744
rect 19337 7735 19395 7741
rect 19337 7701 19349 7735
rect 19383 7732 19395 7735
rect 20438 7732 20444 7744
rect 19383 7704 20444 7732
rect 19383 7701 19395 7704
rect 19337 7695 19395 7701
rect 20438 7692 20444 7704
rect 20496 7692 20502 7744
rect 23400 7732 23428 7763
rect 23658 7760 23664 7772
rect 23716 7760 23722 7812
rect 26528 7809 26556 7908
rect 27341 7905 27353 7908
rect 27387 7936 27399 7939
rect 27522 7936 27528 7948
rect 27387 7908 27528 7936
rect 27387 7905 27399 7908
rect 27341 7899 27399 7905
rect 27522 7896 27528 7908
rect 27580 7896 27586 7948
rect 27617 7939 27675 7945
rect 27617 7905 27629 7939
rect 27663 7936 27675 7939
rect 27798 7936 27804 7948
rect 27663 7908 27804 7936
rect 27663 7905 27675 7908
rect 27617 7899 27675 7905
rect 27798 7896 27804 7908
rect 27856 7936 27862 7948
rect 28534 7936 28540 7948
rect 27856 7908 28540 7936
rect 27856 7896 27862 7908
rect 28534 7896 28540 7908
rect 28592 7896 28598 7948
rect 26694 7868 26700 7880
rect 26655 7840 26700 7868
rect 26694 7828 26700 7840
rect 26752 7828 26758 7880
rect 29086 7828 29092 7880
rect 29144 7868 29150 7880
rect 29549 7871 29607 7877
rect 29549 7868 29561 7871
rect 29144 7840 29561 7868
rect 29144 7828 29150 7840
rect 29549 7837 29561 7840
rect 29595 7837 29607 7871
rect 29656 7868 29684 7976
rect 29730 7964 29736 7976
rect 29788 7964 29794 8016
rect 29822 7964 29828 8016
rect 29880 7964 29886 8016
rect 29712 7871 29770 7877
rect 29840 7874 29868 7964
rect 29712 7868 29724 7871
rect 29656 7840 29724 7868
rect 29549 7831 29607 7837
rect 29712 7837 29724 7840
rect 29758 7837 29770 7871
rect 29712 7831 29770 7837
rect 29828 7868 29886 7874
rect 29937 7871 29995 7877
rect 29937 7868 29949 7871
rect 29828 7834 29840 7868
rect 29874 7834 29886 7868
rect 29932 7837 29949 7868
rect 29983 7862 29995 7871
rect 30116 7862 30144 8044
rect 33778 7964 33784 8016
rect 33836 8004 33842 8016
rect 33836 7976 34192 8004
rect 33836 7964 33842 7976
rect 33686 7896 33692 7948
rect 33744 7936 33750 7948
rect 33744 7908 33913 7936
rect 33744 7896 33750 7908
rect 31202 7868 31208 7880
rect 29983 7837 30144 7862
rect 31163 7840 31208 7868
rect 29932 7834 30144 7837
rect 29828 7828 29886 7834
rect 29937 7831 29995 7834
rect 31202 7828 31208 7840
rect 31260 7828 31266 7880
rect 32950 7828 32956 7880
rect 33008 7868 33014 7880
rect 33885 7877 33913 7908
rect 34164 7877 34192 7976
rect 33781 7871 33839 7877
rect 33781 7868 33793 7871
rect 33008 7840 33793 7868
rect 33008 7828 33014 7840
rect 33781 7837 33793 7840
rect 33827 7837 33839 7871
rect 33781 7831 33839 7837
rect 33870 7871 33928 7877
rect 33870 7837 33882 7871
rect 33916 7837 33928 7871
rect 33870 7831 33928 7837
rect 26513 7803 26571 7809
rect 26513 7800 26525 7803
rect 24504 7772 26525 7800
rect 24504 7732 24532 7772
rect 26513 7769 26525 7772
rect 26559 7769 26571 7803
rect 26513 7763 26571 7769
rect 26605 7803 26663 7809
rect 26605 7769 26617 7803
rect 26651 7769 26663 7803
rect 26605 7763 26663 7769
rect 31472 7803 31530 7809
rect 31472 7769 31484 7803
rect 31518 7800 31530 7803
rect 33505 7803 33563 7809
rect 33505 7800 33517 7803
rect 31518 7772 33517 7800
rect 31518 7769 31530 7772
rect 31472 7763 31530 7769
rect 33505 7769 33517 7772
rect 33551 7769 33563 7803
rect 33505 7763 33563 7769
rect 23400 7704 24532 7732
rect 24581 7735 24639 7741
rect 24581 7701 24593 7735
rect 24627 7732 24639 7735
rect 24854 7732 24860 7744
rect 24627 7704 24860 7732
rect 24627 7701 24639 7704
rect 24581 7695 24639 7701
rect 24854 7692 24860 7704
rect 24912 7732 24918 7744
rect 25590 7732 25596 7744
rect 24912 7704 25596 7732
rect 24912 7692 24918 7704
rect 25590 7692 25596 7704
rect 25648 7692 25654 7744
rect 26234 7692 26240 7744
rect 26292 7732 26298 7744
rect 26620 7732 26648 7763
rect 30190 7732 30196 7744
rect 26292 7704 26648 7732
rect 30151 7704 30196 7732
rect 26292 7692 26298 7704
rect 30190 7692 30196 7704
rect 30248 7692 30254 7744
rect 32582 7732 32588 7744
rect 32543 7704 32588 7732
rect 32582 7692 32588 7704
rect 32640 7692 32646 7744
rect 33796 7732 33824 7831
rect 33962 7822 33968 7874
rect 34020 7862 34026 7874
rect 34149 7871 34207 7877
rect 34020 7834 34065 7862
rect 34149 7837 34161 7871
rect 34195 7868 34207 7871
rect 34238 7868 34244 7880
rect 34195 7840 34244 7868
rect 34195 7837 34207 7840
rect 34020 7822 34026 7834
rect 34149 7831 34207 7837
rect 34238 7828 34244 7840
rect 34296 7828 34302 7880
rect 34348 7868 34376 8044
rect 34514 8032 34520 8084
rect 34572 8072 34578 8084
rect 35253 8075 35311 8081
rect 35253 8072 35265 8075
rect 34572 8044 35265 8072
rect 34572 8032 34578 8044
rect 35253 8041 35265 8044
rect 35299 8041 35311 8075
rect 35253 8035 35311 8041
rect 37185 8075 37243 8081
rect 37185 8041 37197 8075
rect 37231 8072 37243 8075
rect 37274 8072 37280 8084
rect 37231 8044 37280 8072
rect 37231 8041 37243 8044
rect 37185 8035 37243 8041
rect 35268 7936 35296 8035
rect 37274 8032 37280 8044
rect 37332 8032 37338 8084
rect 41230 8072 41236 8084
rect 41191 8044 41236 8072
rect 41230 8032 41236 8044
rect 41288 8032 41294 8084
rect 35805 7939 35863 7945
rect 35805 7936 35817 7939
rect 35268 7908 35817 7936
rect 35805 7905 35817 7908
rect 35851 7905 35863 7939
rect 35805 7899 35863 7905
rect 36081 7939 36139 7945
rect 36081 7905 36093 7939
rect 36127 7936 36139 7939
rect 36170 7936 36176 7948
rect 36127 7908 36176 7936
rect 36127 7905 36139 7908
rect 36081 7899 36139 7905
rect 36170 7896 36176 7908
rect 36228 7936 36234 7948
rect 36998 7936 37004 7948
rect 36228 7908 37004 7936
rect 36228 7896 36234 7908
rect 36998 7896 37004 7908
rect 37056 7896 37062 7948
rect 38838 7936 38844 7948
rect 38120 7908 38844 7936
rect 37366 7868 37372 7880
rect 34348 7840 37372 7868
rect 37366 7828 37372 7840
rect 37424 7828 37430 7880
rect 37550 7828 37556 7880
rect 37608 7868 37614 7880
rect 37918 7868 37924 7880
rect 37608 7840 37924 7868
rect 37608 7828 37614 7840
rect 37918 7828 37924 7840
rect 37976 7828 37982 7880
rect 38120 7877 38148 7908
rect 38838 7896 38844 7908
rect 38896 7896 38902 7948
rect 39850 7936 39856 7948
rect 39811 7908 39856 7936
rect 39850 7896 39856 7908
rect 39908 7896 39914 7948
rect 38084 7871 38148 7877
rect 38084 7837 38096 7871
rect 38130 7840 38148 7871
rect 38200 7871 38258 7877
rect 38200 7868 38212 7871
rect 38130 7837 38142 7840
rect 38084 7831 38142 7837
rect 38199 7837 38212 7868
rect 38246 7837 38258 7871
rect 38199 7831 38258 7837
rect 35986 7760 35992 7812
rect 36044 7800 36050 7812
rect 38199 7800 38227 7831
rect 38286 7828 38292 7880
rect 38344 7868 38350 7880
rect 39025 7871 39083 7877
rect 39025 7868 39037 7871
rect 38344 7840 39037 7868
rect 38344 7828 38350 7840
rect 39025 7837 39037 7840
rect 39071 7837 39083 7871
rect 68094 7868 68100 7880
rect 68055 7840 68100 7868
rect 39025 7831 39083 7837
rect 68094 7828 68100 7840
rect 68152 7828 68158 7880
rect 36044 7772 38227 7800
rect 36044 7760 36050 7772
rect 34701 7735 34759 7741
rect 34701 7732 34713 7735
rect 33796 7704 34713 7732
rect 34701 7701 34713 7704
rect 34747 7701 34759 7735
rect 38199 7732 38227 7772
rect 38565 7803 38623 7809
rect 38565 7769 38577 7803
rect 38611 7800 38623 7803
rect 40098 7803 40156 7809
rect 40098 7800 40110 7803
rect 38611 7772 40110 7800
rect 38611 7769 38623 7772
rect 38565 7763 38623 7769
rect 40098 7769 40110 7772
rect 40144 7769 40156 7803
rect 40098 7763 40156 7769
rect 38378 7732 38384 7744
rect 38199 7704 38384 7732
rect 34701 7695 34759 7701
rect 38378 7692 38384 7704
rect 38436 7692 38442 7744
rect 1104 7642 68816 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 68816 7642
rect 1104 7568 68816 7590
rect 2317 7531 2375 7537
rect 2317 7497 2329 7531
rect 2363 7497 2375 7531
rect 2317 7491 2375 7497
rect 4341 7531 4399 7537
rect 4341 7497 4353 7531
rect 4387 7528 4399 7531
rect 4430 7528 4436 7540
rect 4387 7500 4436 7528
rect 4387 7497 4399 7500
rect 4341 7491 4399 7497
rect 2332 7460 2360 7491
rect 4430 7488 4436 7500
rect 4488 7488 4494 7540
rect 4798 7488 4804 7540
rect 4856 7528 4862 7540
rect 5261 7531 5319 7537
rect 5261 7528 5273 7531
rect 4856 7500 5273 7528
rect 4856 7488 4862 7500
rect 5261 7497 5273 7500
rect 5307 7497 5319 7531
rect 8573 7531 8631 7537
rect 5261 7491 5319 7497
rect 6932 7500 8340 7528
rect 3206 7463 3264 7469
rect 3206 7460 3218 7463
rect 2332 7432 3218 7460
rect 3206 7429 3218 7432
rect 3252 7429 3264 7463
rect 3206 7423 3264 7429
rect 2130 7392 2136 7404
rect 2091 7364 2136 7392
rect 2130 7352 2136 7364
rect 2188 7352 2194 7404
rect 5445 7395 5503 7401
rect 5445 7361 5457 7395
rect 5491 7392 5503 7395
rect 6362 7392 6368 7404
rect 5491 7364 6368 7392
rect 5491 7361 5503 7364
rect 5445 7355 5503 7361
rect 6362 7352 6368 7364
rect 6420 7352 6426 7404
rect 6932 7392 6960 7500
rect 8312 7472 8340 7500
rect 8573 7497 8585 7531
rect 8619 7528 8631 7531
rect 10686 7528 10692 7540
rect 8619 7500 10692 7528
rect 8619 7497 8631 7500
rect 8573 7491 8631 7497
rect 10686 7488 10692 7500
rect 10744 7488 10750 7540
rect 14918 7528 14924 7540
rect 12176 7500 14596 7528
rect 14879 7500 14924 7528
rect 8205 7463 8263 7469
rect 8205 7460 8217 7463
rect 7116 7432 8217 7460
rect 7009 7395 7067 7401
rect 7009 7392 7021 7395
rect 6932 7364 7021 7392
rect 7009 7361 7021 7364
rect 7055 7361 7067 7395
rect 7009 7355 7067 7361
rect 1673 7327 1731 7333
rect 1673 7293 1685 7327
rect 1719 7324 1731 7327
rect 2682 7324 2688 7336
rect 1719 7296 2688 7324
rect 1719 7293 1731 7296
rect 1673 7287 1731 7293
rect 2682 7284 2688 7296
rect 2740 7284 2746 7336
rect 2958 7324 2964 7336
rect 2919 7296 2964 7324
rect 2958 7284 2964 7296
rect 3016 7284 3022 7336
rect 5629 7327 5687 7333
rect 5629 7293 5641 7327
rect 5675 7324 5687 7327
rect 6914 7324 6920 7336
rect 5675 7296 6920 7324
rect 5675 7293 5687 7296
rect 5629 7287 5687 7293
rect 6914 7284 6920 7296
rect 6972 7284 6978 7336
rect 5810 7216 5816 7268
rect 5868 7256 5874 7268
rect 5868 7228 6592 7256
rect 5868 7216 5874 7228
rect 6086 7148 6092 7200
rect 6144 7188 6150 7200
rect 6454 7188 6460 7200
rect 6144 7160 6460 7188
rect 6144 7148 6150 7160
rect 6454 7148 6460 7160
rect 6512 7148 6518 7200
rect 6564 7188 6592 7228
rect 7116 7188 7144 7432
rect 8205 7429 8217 7432
rect 8251 7429 8263 7463
rect 8205 7423 8263 7429
rect 8294 7420 8300 7472
rect 8352 7460 8358 7472
rect 9214 7460 9220 7472
rect 8352 7432 9220 7460
rect 8352 7420 8358 7432
rect 9214 7420 9220 7432
rect 9272 7420 9278 7472
rect 10965 7463 11023 7469
rect 10965 7429 10977 7463
rect 11011 7460 11023 7463
rect 12066 7460 12072 7472
rect 11011 7432 12072 7460
rect 11011 7429 11023 7432
rect 10965 7423 11023 7429
rect 12066 7420 12072 7432
rect 12124 7420 12130 7472
rect 8113 7395 8171 7401
rect 8113 7361 8125 7395
rect 8159 7361 8171 7395
rect 8386 7392 8392 7404
rect 8347 7364 8392 7392
rect 8113 7355 8171 7361
rect 7650 7284 7656 7336
rect 7708 7324 7714 7336
rect 8128 7324 8156 7355
rect 8386 7352 8392 7364
rect 8444 7352 8450 7404
rect 9033 7395 9091 7401
rect 9033 7361 9045 7395
rect 9079 7392 9091 7395
rect 9674 7392 9680 7404
rect 9079 7364 9680 7392
rect 9079 7361 9091 7364
rect 9033 7355 9091 7361
rect 9674 7352 9680 7364
rect 9732 7392 9738 7404
rect 10134 7392 10140 7404
rect 9732 7364 10140 7392
rect 9732 7352 9738 7364
rect 10134 7352 10140 7364
rect 10192 7352 10198 7404
rect 10781 7395 10839 7401
rect 10781 7361 10793 7395
rect 10827 7392 10839 7395
rect 11054 7392 11060 7404
rect 10827 7364 11060 7392
rect 10827 7361 10839 7364
rect 10781 7355 10839 7361
rect 9309 7327 9367 7333
rect 9309 7324 9321 7327
rect 7708 7296 9321 7324
rect 7708 7284 7714 7296
rect 9309 7293 9321 7296
rect 9355 7293 9367 7327
rect 9309 7287 9367 7293
rect 7190 7216 7196 7268
rect 7248 7256 7254 7268
rect 10796 7256 10824 7355
rect 11054 7352 11060 7364
rect 11112 7392 11118 7404
rect 11793 7395 11851 7401
rect 11112 7364 11744 7392
rect 11112 7352 11118 7364
rect 11517 7327 11575 7333
rect 11517 7293 11529 7327
rect 11563 7324 11575 7327
rect 11606 7324 11612 7336
rect 11563 7296 11612 7324
rect 11563 7293 11575 7296
rect 11517 7287 11575 7293
rect 11606 7284 11612 7296
rect 11664 7284 11670 7336
rect 11716 7324 11744 7364
rect 11793 7361 11805 7395
rect 11839 7392 11851 7395
rect 11974 7392 11980 7404
rect 11839 7364 11980 7392
rect 11839 7361 11851 7364
rect 11793 7355 11851 7361
rect 11974 7352 11980 7364
rect 12032 7392 12038 7404
rect 12176 7392 12204 7500
rect 13814 7460 13820 7472
rect 12032 7364 12204 7392
rect 12406 7432 12756 7460
rect 12032 7352 12038 7364
rect 12406 7324 12434 7432
rect 11716 7296 12434 7324
rect 12728 7324 12756 7432
rect 13004 7432 13820 7460
rect 13004 7401 13032 7432
rect 13814 7420 13820 7432
rect 13872 7420 13878 7472
rect 12989 7395 13047 7401
rect 12989 7361 13001 7395
rect 13035 7361 13047 7395
rect 12989 7355 13047 7361
rect 13633 7395 13691 7401
rect 13633 7361 13645 7395
rect 13679 7392 13691 7395
rect 13998 7392 14004 7404
rect 13679 7364 14004 7392
rect 13679 7361 13691 7364
rect 13633 7355 13691 7361
rect 13998 7352 14004 7364
rect 14056 7352 14062 7404
rect 14274 7392 14280 7404
rect 14235 7364 14280 7392
rect 14274 7352 14280 7364
rect 14332 7352 14338 7404
rect 14568 7401 14596 7500
rect 14918 7488 14924 7500
rect 14976 7488 14982 7540
rect 16945 7531 17003 7537
rect 16945 7497 16957 7531
rect 16991 7528 17003 7531
rect 23566 7528 23572 7540
rect 16991 7500 23572 7528
rect 16991 7497 17003 7500
rect 16945 7491 17003 7497
rect 23566 7488 23572 7500
rect 23624 7488 23630 7540
rect 23845 7531 23903 7537
rect 23845 7497 23857 7531
rect 23891 7528 23903 7531
rect 24946 7528 24952 7540
rect 23891 7500 24952 7528
rect 23891 7497 23903 7500
rect 23845 7491 23903 7497
rect 24946 7488 24952 7500
rect 25004 7488 25010 7540
rect 27893 7531 27951 7537
rect 27893 7497 27905 7531
rect 27939 7528 27951 7531
rect 28074 7528 28080 7540
rect 27939 7500 28080 7528
rect 27939 7497 27951 7500
rect 27893 7491 27951 7497
rect 28074 7488 28080 7500
rect 28132 7488 28138 7540
rect 28905 7531 28963 7537
rect 28905 7497 28917 7531
rect 28951 7528 28963 7531
rect 28994 7528 29000 7540
rect 28951 7500 29000 7528
rect 28951 7497 28963 7500
rect 28905 7491 28963 7497
rect 28994 7488 29000 7500
rect 29052 7488 29058 7540
rect 29454 7488 29460 7540
rect 29512 7528 29518 7540
rect 29733 7531 29791 7537
rect 29733 7528 29745 7531
rect 29512 7500 29745 7528
rect 29512 7488 29518 7500
rect 29733 7497 29745 7500
rect 29779 7497 29791 7531
rect 29733 7491 29791 7497
rect 33597 7531 33655 7537
rect 33597 7497 33609 7531
rect 33643 7528 33655 7531
rect 33962 7528 33968 7540
rect 33643 7500 33968 7528
rect 33643 7497 33655 7500
rect 33597 7491 33655 7497
rect 33962 7488 33968 7500
rect 34020 7488 34026 7540
rect 37366 7528 37372 7540
rect 37327 7500 37372 7528
rect 37366 7488 37372 7500
rect 37424 7528 37430 7540
rect 38470 7528 38476 7540
rect 37424 7500 38476 7528
rect 37424 7488 37430 7500
rect 38470 7488 38476 7500
rect 38528 7488 38534 7540
rect 38746 7488 38752 7540
rect 38804 7528 38810 7540
rect 39025 7531 39083 7537
rect 39025 7528 39037 7531
rect 38804 7500 39037 7528
rect 38804 7488 38810 7500
rect 39025 7497 39037 7500
rect 39071 7497 39083 7531
rect 39025 7491 39083 7497
rect 15102 7420 15108 7472
rect 15160 7460 15166 7472
rect 18693 7463 18751 7469
rect 15160 7432 16896 7460
rect 15160 7420 15166 7432
rect 14461 7395 14519 7401
rect 14461 7361 14473 7395
rect 14507 7361 14519 7395
rect 14461 7355 14519 7361
rect 14553 7395 14611 7401
rect 14553 7361 14565 7395
rect 14599 7361 14611 7395
rect 14553 7355 14611 7361
rect 14645 7395 14703 7401
rect 14645 7361 14657 7395
rect 14691 7392 14703 7395
rect 14826 7392 14832 7404
rect 14691 7364 14832 7392
rect 14691 7361 14703 7364
rect 14645 7355 14703 7361
rect 13538 7324 13544 7336
rect 12728 7296 13544 7324
rect 13538 7284 13544 7296
rect 13596 7284 13602 7336
rect 14476 7324 14504 7355
rect 14826 7352 14832 7364
rect 14884 7352 14890 7404
rect 16666 7392 16672 7404
rect 16627 7364 16672 7392
rect 16666 7352 16672 7364
rect 16724 7352 16730 7404
rect 16868 7401 16896 7432
rect 18693 7429 18705 7463
rect 18739 7460 18751 7463
rect 19978 7460 19984 7472
rect 18739 7432 19984 7460
rect 18739 7429 18751 7432
rect 18693 7423 18751 7429
rect 19978 7420 19984 7432
rect 20036 7420 20042 7472
rect 23658 7420 23664 7472
rect 23716 7460 23722 7472
rect 24489 7463 24547 7469
rect 24489 7460 24501 7463
rect 23716 7432 24501 7460
rect 23716 7420 23722 7432
rect 24489 7429 24501 7432
rect 24535 7429 24547 7463
rect 27522 7460 27528 7472
rect 27483 7432 27528 7460
rect 24489 7423 24547 7429
rect 27522 7420 27528 7432
rect 27580 7420 27586 7472
rect 27617 7463 27675 7469
rect 27617 7429 27629 7463
rect 27663 7460 27675 7463
rect 28442 7460 28448 7472
rect 27663 7432 28448 7460
rect 27663 7429 27675 7432
rect 27617 7423 27675 7429
rect 28442 7420 28448 7432
rect 28500 7420 28506 7472
rect 28629 7463 28687 7469
rect 28629 7429 28641 7463
rect 28675 7460 28687 7463
rect 29638 7460 29644 7472
rect 28675 7432 29644 7460
rect 28675 7429 28687 7432
rect 28629 7423 28687 7429
rect 29638 7420 29644 7432
rect 29696 7420 29702 7472
rect 30190 7420 30196 7472
rect 30248 7460 30254 7472
rect 30846 7463 30904 7469
rect 30846 7460 30858 7463
rect 30248 7432 30858 7460
rect 30248 7420 30254 7432
rect 30846 7429 30858 7432
rect 30892 7429 30904 7463
rect 30846 7423 30904 7429
rect 32582 7420 32588 7472
rect 32640 7460 32646 7472
rect 33781 7463 33839 7469
rect 33781 7460 33793 7463
rect 32640 7432 33793 7460
rect 32640 7420 32646 7432
rect 33781 7429 33793 7432
rect 33827 7429 33839 7463
rect 34793 7463 34851 7469
rect 34793 7460 34805 7463
rect 33781 7423 33839 7429
rect 33980 7432 34805 7460
rect 16853 7395 16911 7401
rect 16853 7361 16865 7395
rect 16899 7361 16911 7395
rect 18506 7392 18512 7404
rect 18467 7364 18512 7392
rect 16853 7355 16911 7361
rect 18506 7352 18512 7364
rect 18564 7352 18570 7404
rect 18785 7395 18843 7401
rect 18785 7361 18797 7395
rect 18831 7392 18843 7395
rect 21542 7392 21548 7404
rect 18831 7364 21548 7392
rect 18831 7361 18843 7364
rect 18785 7355 18843 7361
rect 21542 7352 21548 7364
rect 21600 7352 21606 7404
rect 22646 7392 22652 7404
rect 22607 7364 22652 7392
rect 22646 7352 22652 7364
rect 22704 7352 22710 7404
rect 24305 7395 24363 7401
rect 24305 7361 24317 7395
rect 24351 7392 24363 7395
rect 24854 7392 24860 7404
rect 24351 7364 24860 7392
rect 24351 7361 24363 7364
rect 24305 7355 24363 7361
rect 24854 7352 24860 7364
rect 24912 7352 24918 7404
rect 25314 7352 25320 7404
rect 25372 7401 25378 7404
rect 25372 7395 25421 7401
rect 25372 7361 25375 7395
rect 25409 7361 25421 7395
rect 25372 7355 25421 7361
rect 25498 7395 25556 7401
rect 25498 7361 25510 7395
rect 25544 7361 25556 7395
rect 25614 7395 25672 7401
rect 25614 7392 25626 7395
rect 25498 7355 25556 7361
rect 25608 7361 25626 7392
rect 25660 7361 25672 7395
rect 25608 7355 25672 7361
rect 25372 7352 25378 7355
rect 18325 7327 18383 7333
rect 18325 7324 18337 7327
rect 14476 7296 18337 7324
rect 18325 7293 18337 7296
rect 18371 7293 18383 7327
rect 18325 7287 18383 7293
rect 18414 7284 18420 7336
rect 18472 7324 18478 7336
rect 19797 7327 19855 7333
rect 19797 7324 19809 7327
rect 18472 7296 19809 7324
rect 18472 7284 18478 7296
rect 19797 7293 19809 7296
rect 19843 7293 19855 7327
rect 22370 7324 22376 7336
rect 22331 7296 22376 7324
rect 19797 7287 19855 7293
rect 22370 7284 22376 7296
rect 22428 7284 22434 7336
rect 25038 7284 25044 7336
rect 25096 7324 25102 7336
rect 25516 7324 25544 7355
rect 25096 7296 25544 7324
rect 25096 7284 25102 7296
rect 7248 7228 10824 7256
rect 13817 7259 13875 7265
rect 7248 7216 7254 7228
rect 13817 7225 13829 7259
rect 13863 7256 13875 7259
rect 19702 7256 19708 7268
rect 13863 7228 19708 7256
rect 13863 7225 13875 7228
rect 13817 7219 13875 7225
rect 19702 7216 19708 7228
rect 19760 7216 19766 7268
rect 24673 7259 24731 7265
rect 24673 7225 24685 7259
rect 24719 7256 24731 7259
rect 25608 7256 25636 7355
rect 25774 7352 25780 7404
rect 25832 7392 25838 7404
rect 27338 7392 27344 7404
rect 25832 7364 26464 7392
rect 27299 7364 27344 7392
rect 25832 7352 25838 7364
rect 24719 7228 25636 7256
rect 24719 7225 24731 7228
rect 24673 7219 24731 7225
rect 26436 7200 26464 7364
rect 27338 7352 27344 7364
rect 27396 7352 27402 7404
rect 27706 7392 27712 7404
rect 27667 7364 27712 7392
rect 27706 7352 27712 7364
rect 27764 7352 27770 7404
rect 27798 7352 27804 7404
rect 27856 7392 27862 7404
rect 28353 7395 28411 7401
rect 28353 7392 28365 7395
rect 27856 7364 28365 7392
rect 27856 7352 27862 7364
rect 28353 7361 28365 7364
rect 28399 7361 28411 7395
rect 28534 7392 28540 7404
rect 28495 7364 28540 7392
rect 28353 7355 28411 7361
rect 28534 7352 28540 7364
rect 28592 7352 28598 7404
rect 28721 7395 28779 7401
rect 28721 7361 28733 7395
rect 28767 7361 28779 7395
rect 28721 7355 28779 7361
rect 27724 7324 27752 7352
rect 28736 7324 28764 7355
rect 29546 7352 29552 7404
rect 29604 7392 29610 7404
rect 33980 7401 34008 7432
rect 34793 7429 34805 7432
rect 34839 7460 34851 7463
rect 35894 7460 35900 7472
rect 34839 7432 35900 7460
rect 34839 7429 34851 7432
rect 34793 7423 34851 7429
rect 35894 7420 35900 7432
rect 35952 7420 35958 7472
rect 36170 7460 36176 7472
rect 36131 7432 36176 7460
rect 36170 7420 36176 7432
rect 36228 7420 36234 7472
rect 33965 7395 34023 7401
rect 29604 7364 31800 7392
rect 29604 7352 29610 7364
rect 27724 7296 28764 7324
rect 31113 7327 31171 7333
rect 31113 7293 31125 7327
rect 31159 7324 31171 7327
rect 31202 7324 31208 7336
rect 31159 7296 31208 7324
rect 31159 7293 31171 7296
rect 31113 7287 31171 7293
rect 31202 7284 31208 7296
rect 31260 7324 31266 7336
rect 31570 7324 31576 7336
rect 31260 7296 31576 7324
rect 31260 7284 31266 7296
rect 31570 7284 31576 7296
rect 31628 7284 31634 7336
rect 31772 7256 31800 7364
rect 33965 7361 33977 7395
rect 34011 7361 34023 7395
rect 33965 7355 34023 7361
rect 34422 7352 34428 7404
rect 34480 7392 34486 7404
rect 34609 7395 34667 7401
rect 34609 7392 34621 7395
rect 34480 7364 34621 7392
rect 34480 7352 34486 7364
rect 34609 7361 34621 7364
rect 34655 7361 34667 7395
rect 34609 7355 34667 7361
rect 35989 7395 36047 7401
rect 35989 7361 36001 7395
rect 36035 7361 36047 7395
rect 35989 7355 36047 7361
rect 36004 7324 36032 7355
rect 36078 7352 36084 7404
rect 36136 7392 36142 7404
rect 36354 7392 36360 7404
rect 36136 7364 36181 7392
rect 36315 7364 36360 7392
rect 36136 7352 36142 7364
rect 36354 7352 36360 7364
rect 36412 7352 36418 7404
rect 37918 7392 37924 7404
rect 37879 7364 37924 7392
rect 37918 7352 37924 7364
rect 37976 7352 37982 7404
rect 38105 7395 38163 7401
rect 38028 7367 38117 7395
rect 37090 7324 37096 7336
rect 36004 7296 37096 7324
rect 37090 7284 37096 7296
rect 37148 7284 37154 7336
rect 35805 7259 35863 7265
rect 35805 7256 35817 7259
rect 31772 7228 35817 7256
rect 35805 7225 35817 7228
rect 35851 7225 35863 7259
rect 38028 7256 38056 7367
rect 38105 7361 38117 7367
rect 38151 7361 38163 7395
rect 38105 7355 38163 7361
rect 38200 7395 38258 7401
rect 38200 7361 38212 7395
rect 38246 7361 38258 7395
rect 38200 7355 38258 7361
rect 38289 7398 38347 7401
rect 38470 7398 38476 7404
rect 38289 7395 38476 7398
rect 38289 7361 38301 7395
rect 38335 7370 38476 7395
rect 38335 7361 38347 7370
rect 38289 7355 38347 7361
rect 38212 7324 38240 7355
rect 38470 7352 38476 7370
rect 38528 7352 38534 7404
rect 38378 7324 38384 7336
rect 38212 7296 38384 7324
rect 38378 7284 38384 7296
rect 38436 7284 38442 7336
rect 38194 7256 38200 7268
rect 38028 7228 38200 7256
rect 35805 7219 35863 7225
rect 38194 7216 38200 7228
rect 38252 7216 38258 7268
rect 6564 7160 7144 7188
rect 13173 7191 13231 7197
rect 13173 7157 13185 7191
rect 13219 7188 13231 7191
rect 13906 7188 13912 7200
rect 13219 7160 13912 7188
rect 13219 7157 13231 7160
rect 13173 7151 13231 7157
rect 13906 7148 13912 7160
rect 13964 7148 13970 7200
rect 13998 7148 14004 7200
rect 14056 7188 14062 7200
rect 14734 7188 14740 7200
rect 14056 7160 14740 7188
rect 14056 7148 14062 7160
rect 14734 7148 14740 7160
rect 14792 7188 14798 7200
rect 15381 7191 15439 7197
rect 15381 7188 15393 7191
rect 14792 7160 15393 7188
rect 14792 7148 14798 7160
rect 15381 7157 15393 7160
rect 15427 7157 15439 7191
rect 16114 7188 16120 7200
rect 16075 7160 16120 7188
rect 15381 7151 15439 7157
rect 16114 7148 16120 7160
rect 16172 7148 16178 7200
rect 17494 7148 17500 7200
rect 17552 7188 17558 7200
rect 17589 7191 17647 7197
rect 17589 7188 17601 7191
rect 17552 7160 17601 7188
rect 17552 7148 17558 7160
rect 17589 7157 17601 7160
rect 17635 7157 17647 7191
rect 17589 7151 17647 7157
rect 19337 7191 19395 7197
rect 19337 7157 19349 7191
rect 19383 7188 19395 7191
rect 20254 7188 20260 7200
rect 19383 7160 20260 7188
rect 19383 7157 19395 7160
rect 19337 7151 19395 7157
rect 20254 7148 20260 7160
rect 20312 7148 20318 7200
rect 23842 7148 23848 7200
rect 23900 7188 23906 7200
rect 25133 7191 25191 7197
rect 25133 7188 25145 7191
rect 23900 7160 25145 7188
rect 23900 7148 23906 7160
rect 25133 7157 25145 7160
rect 25179 7157 25191 7191
rect 25133 7151 25191 7157
rect 25314 7148 25320 7200
rect 25372 7188 25378 7200
rect 26326 7188 26332 7200
rect 25372 7160 26332 7188
rect 25372 7148 25378 7160
rect 26326 7148 26332 7160
rect 26384 7148 26390 7200
rect 26418 7148 26424 7200
rect 26476 7188 26482 7200
rect 29086 7188 29092 7200
rect 26476 7160 29092 7188
rect 26476 7148 26482 7160
rect 29086 7148 29092 7160
rect 29144 7148 29150 7200
rect 34054 7148 34060 7200
rect 34112 7188 34118 7200
rect 34425 7191 34483 7197
rect 34425 7188 34437 7191
rect 34112 7160 34437 7188
rect 34112 7148 34118 7160
rect 34425 7157 34437 7160
rect 34471 7157 34483 7191
rect 34425 7151 34483 7157
rect 38565 7191 38623 7197
rect 38565 7157 38577 7191
rect 38611 7188 38623 7191
rect 39942 7188 39948 7200
rect 38611 7160 39948 7188
rect 38611 7157 38623 7160
rect 38565 7151 38623 7157
rect 39942 7148 39948 7160
rect 40000 7148 40006 7200
rect 1104 7098 68816 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 65654 7098
rect 65706 7046 65718 7098
rect 65770 7046 65782 7098
rect 65834 7046 65846 7098
rect 65898 7046 65910 7098
rect 65962 7046 68816 7098
rect 1104 7024 68816 7046
rect 2041 6987 2099 6993
rect 2041 6953 2053 6987
rect 2087 6984 2099 6987
rect 2130 6984 2136 6996
rect 2087 6956 2136 6984
rect 2087 6953 2099 6956
rect 2041 6947 2099 6953
rect 2130 6944 2136 6956
rect 2188 6944 2194 6996
rect 6362 6984 6368 6996
rect 6323 6956 6368 6984
rect 6362 6944 6368 6956
rect 6420 6944 6426 6996
rect 12802 6944 12808 6996
rect 12860 6984 12866 6996
rect 13170 6984 13176 6996
rect 12860 6956 13176 6984
rect 12860 6944 12866 6956
rect 13170 6944 13176 6956
rect 13228 6984 13234 6996
rect 16666 6984 16672 6996
rect 13228 6956 16672 6984
rect 13228 6944 13234 6956
rect 16666 6944 16672 6956
rect 16724 6944 16730 6996
rect 33413 6987 33471 6993
rect 33413 6953 33425 6987
rect 33459 6984 33471 6987
rect 34422 6984 34428 6996
rect 33459 6956 34428 6984
rect 33459 6953 33471 6956
rect 33413 6947 33471 6953
rect 34422 6944 34428 6956
rect 34480 6944 34486 6996
rect 36354 6944 36360 6996
rect 36412 6984 36418 6996
rect 36725 6987 36783 6993
rect 36725 6984 36737 6987
rect 36412 6956 36737 6984
rect 36412 6944 36418 6956
rect 36725 6953 36737 6956
rect 36771 6953 36783 6987
rect 38194 6984 38200 6996
rect 38155 6956 38200 6984
rect 36725 6947 36783 6953
rect 38194 6944 38200 6956
rect 38252 6944 38258 6996
rect 9858 6876 9864 6928
rect 9916 6916 9922 6928
rect 9916 6888 9961 6916
rect 10428 6888 10732 6916
rect 9916 6876 9922 6888
rect 1673 6851 1731 6857
rect 1673 6817 1685 6851
rect 1719 6848 1731 6851
rect 1762 6848 1768 6860
rect 1719 6820 1768 6848
rect 1719 6817 1731 6820
rect 1673 6811 1731 6817
rect 1762 6808 1768 6820
rect 1820 6808 1826 6860
rect 3237 6851 3295 6857
rect 3237 6817 3249 6851
rect 3283 6848 3295 6851
rect 5902 6848 5908 6860
rect 3283 6820 5908 6848
rect 3283 6817 3295 6820
rect 3237 6811 3295 6817
rect 5902 6808 5908 6820
rect 5960 6808 5966 6860
rect 6822 6848 6828 6860
rect 6783 6820 6828 6848
rect 6822 6808 6828 6820
rect 6880 6808 6886 6860
rect 6917 6851 6975 6857
rect 6917 6817 6929 6851
rect 6963 6817 6975 6851
rect 8110 6848 8116 6860
rect 8071 6820 8116 6848
rect 6917 6811 6975 6817
rect 1854 6780 1860 6792
rect 1815 6752 1860 6780
rect 1854 6740 1860 6752
rect 1912 6740 1918 6792
rect 2685 6783 2743 6789
rect 2685 6749 2697 6783
rect 2731 6780 2743 6783
rect 5074 6780 5080 6792
rect 2731 6752 5080 6780
rect 2731 6749 2743 6752
rect 2685 6743 2743 6749
rect 5074 6740 5080 6752
rect 5132 6740 5138 6792
rect 6638 6740 6644 6792
rect 6696 6780 6702 6792
rect 6932 6780 6960 6811
rect 8110 6808 8116 6820
rect 8168 6808 8174 6860
rect 9766 6848 9772 6860
rect 9324 6820 9772 6848
rect 7650 6780 7656 6792
rect 6696 6752 6960 6780
rect 7611 6752 7656 6780
rect 6696 6740 6702 6752
rect 7650 6740 7656 6752
rect 7708 6740 7714 6792
rect 7926 6780 7932 6792
rect 7887 6752 7932 6780
rect 7926 6740 7932 6752
rect 7984 6740 7990 6792
rect 9324 6789 9352 6820
rect 9766 6808 9772 6820
rect 9824 6808 9830 6860
rect 10428 6848 10456 6888
rect 10594 6848 10600 6860
rect 10336 6820 10456 6848
rect 10555 6820 10600 6848
rect 9125 6783 9183 6789
rect 9125 6749 9137 6783
rect 9171 6749 9183 6783
rect 9125 6743 9183 6749
rect 9309 6783 9367 6789
rect 9309 6749 9321 6783
rect 9355 6749 9367 6783
rect 9309 6743 9367 6749
rect 9401 6783 9459 6789
rect 9401 6749 9413 6783
rect 9447 6749 9459 6783
rect 9401 6743 9459 6749
rect 4157 6715 4215 6721
rect 4157 6681 4169 6715
rect 4203 6712 4215 6715
rect 5534 6712 5540 6724
rect 4203 6684 5540 6712
rect 4203 6681 4215 6684
rect 4157 6675 4215 6681
rect 5534 6672 5540 6684
rect 5592 6672 5598 6724
rect 6914 6672 6920 6724
rect 6972 6712 6978 6724
rect 9140 6712 9168 6743
rect 6972 6684 9168 6712
rect 6972 6672 6978 6684
rect 4614 6604 4620 6656
rect 4672 6644 4678 6656
rect 5445 6647 5503 6653
rect 5445 6644 5457 6647
rect 4672 6616 5457 6644
rect 4672 6604 4678 6616
rect 5445 6613 5457 6616
rect 5491 6613 5503 6647
rect 5445 6607 5503 6613
rect 6454 6604 6460 6656
rect 6512 6644 6518 6656
rect 6733 6647 6791 6653
rect 6733 6644 6745 6647
rect 6512 6616 6745 6644
rect 6512 6604 6518 6616
rect 6733 6613 6745 6616
rect 6779 6644 6791 6647
rect 6822 6644 6828 6656
rect 6779 6616 6828 6644
rect 6779 6613 6791 6616
rect 6733 6607 6791 6613
rect 6822 6604 6828 6616
rect 6880 6604 6886 6656
rect 7006 6604 7012 6656
rect 7064 6644 7070 6656
rect 7745 6647 7803 6653
rect 7745 6644 7757 6647
rect 7064 6616 7757 6644
rect 7064 6604 7070 6616
rect 7745 6613 7757 6616
rect 7791 6613 7803 6647
rect 9140 6644 9168 6684
rect 9214 6672 9220 6724
rect 9272 6712 9278 6724
rect 9416 6712 9444 6743
rect 9490 6740 9496 6792
rect 9548 6780 9554 6792
rect 9674 6780 9680 6792
rect 9548 6752 9593 6780
rect 9635 6752 9680 6780
rect 9548 6740 9554 6752
rect 9674 6740 9680 6752
rect 9732 6740 9738 6792
rect 10336 6789 10364 6820
rect 10594 6808 10600 6820
rect 10652 6808 10658 6860
rect 10704 6848 10732 6888
rect 25038 6876 25044 6928
rect 25096 6916 25102 6928
rect 29822 6916 29828 6928
rect 25096 6888 29828 6916
rect 25096 6876 25102 6888
rect 12161 6851 12219 6857
rect 10704 6820 12112 6848
rect 10321 6783 10379 6789
rect 10321 6780 10333 6783
rect 9784 6752 10333 6780
rect 9272 6684 9444 6712
rect 9272 6672 9278 6684
rect 9784 6644 9812 6752
rect 10321 6749 10333 6752
rect 10367 6749 10379 6783
rect 10321 6743 10379 6749
rect 10505 6783 10563 6789
rect 10505 6749 10517 6783
rect 10551 6749 10563 6783
rect 10686 6780 10692 6792
rect 10647 6752 10692 6780
rect 10505 6743 10563 6749
rect 10042 6672 10048 6724
rect 10100 6712 10106 6724
rect 10520 6712 10548 6743
rect 10686 6740 10692 6752
rect 10744 6740 10750 6792
rect 10873 6783 10931 6789
rect 10873 6749 10885 6783
rect 10919 6780 10931 6783
rect 11698 6780 11704 6792
rect 10919 6752 11704 6780
rect 10919 6749 10931 6752
rect 10873 6743 10931 6749
rect 11698 6740 11704 6752
rect 11756 6740 11762 6792
rect 10100 6684 10548 6712
rect 10704 6712 10732 6740
rect 11606 6712 11612 6724
rect 10704 6684 11612 6712
rect 10100 6672 10106 6684
rect 11606 6672 11612 6684
rect 11664 6712 11670 6724
rect 11977 6715 12035 6721
rect 11977 6712 11989 6715
rect 11664 6684 11989 6712
rect 11664 6672 11670 6684
rect 11977 6681 11989 6684
rect 12023 6681 12035 6715
rect 12084 6712 12112 6820
rect 12161 6817 12173 6851
rect 12207 6848 12219 6851
rect 12618 6848 12624 6860
rect 12207 6820 12624 6848
rect 12207 6817 12219 6820
rect 12161 6811 12219 6817
rect 12618 6808 12624 6820
rect 12676 6808 12682 6860
rect 14553 6851 14611 6857
rect 14553 6817 14565 6851
rect 14599 6848 14611 6851
rect 15470 6848 15476 6860
rect 14599 6820 15476 6848
rect 14599 6817 14611 6820
rect 14553 6811 14611 6817
rect 15470 6808 15476 6820
rect 15528 6808 15534 6860
rect 16298 6848 16304 6860
rect 16259 6820 16304 6848
rect 16298 6808 16304 6820
rect 16356 6808 16362 6860
rect 18601 6851 18659 6857
rect 18601 6817 18613 6851
rect 18647 6848 18659 6851
rect 20530 6848 20536 6860
rect 18647 6820 20392 6848
rect 20491 6820 20536 6848
rect 18647 6817 18659 6820
rect 18601 6811 18659 6817
rect 12897 6783 12955 6789
rect 12897 6749 12909 6783
rect 12943 6780 12955 6783
rect 13354 6780 13360 6792
rect 12943 6752 13360 6780
rect 12943 6749 12955 6752
rect 12897 6743 12955 6749
rect 13354 6740 13360 6752
rect 13412 6740 13418 6792
rect 13541 6783 13599 6789
rect 13541 6749 13553 6783
rect 13587 6780 13599 6783
rect 13722 6780 13728 6792
rect 13587 6752 13728 6780
rect 13587 6749 13599 6752
rect 13541 6743 13599 6749
rect 13722 6740 13728 6752
rect 13780 6740 13786 6792
rect 15197 6783 15255 6789
rect 15197 6749 15209 6783
rect 15243 6780 15255 6783
rect 15746 6780 15752 6792
rect 15243 6752 15752 6780
rect 15243 6749 15255 6752
rect 15197 6743 15255 6749
rect 15746 6740 15752 6752
rect 15804 6740 15810 6792
rect 15841 6783 15899 6789
rect 15841 6749 15853 6783
rect 15887 6780 15899 6783
rect 16390 6780 16396 6792
rect 15887 6752 16396 6780
rect 15887 6749 15899 6752
rect 15841 6743 15899 6749
rect 16390 6740 16396 6752
rect 16448 6740 16454 6792
rect 18506 6780 18512 6792
rect 18467 6752 18512 6780
rect 18506 6740 18512 6752
rect 18564 6740 18570 6792
rect 18693 6783 18751 6789
rect 18693 6749 18705 6783
rect 18739 6749 18751 6783
rect 19426 6780 19432 6792
rect 19387 6752 19432 6780
rect 18693 6743 18751 6749
rect 15930 6712 15936 6724
rect 12084 6684 15936 6712
rect 11977 6675 12035 6681
rect 15930 6672 15936 6684
rect 15988 6672 15994 6724
rect 16568 6715 16626 6721
rect 16568 6681 16580 6715
rect 16614 6712 16626 6715
rect 16666 6712 16672 6724
rect 16614 6684 16672 6712
rect 16614 6681 16626 6684
rect 16568 6675 16626 6681
rect 16666 6672 16672 6684
rect 16724 6672 16730 6724
rect 17218 6672 17224 6724
rect 17276 6712 17282 6724
rect 18708 6712 18736 6743
rect 19426 6740 19432 6752
rect 19484 6740 19490 6792
rect 19613 6783 19671 6789
rect 19613 6749 19625 6783
rect 19659 6749 19671 6783
rect 19613 6743 19671 6749
rect 19705 6783 19763 6789
rect 19705 6749 19717 6783
rect 19751 6749 19763 6783
rect 19705 6743 19763 6749
rect 17276 6684 18736 6712
rect 17276 6672 17282 6684
rect 11054 6644 11060 6656
rect 9140 6616 9812 6644
rect 11015 6616 11060 6644
rect 7745 6607 7803 6613
rect 11054 6604 11060 6616
rect 11112 6604 11118 6656
rect 11146 6604 11152 6656
rect 11204 6644 11210 6656
rect 12342 6644 12348 6656
rect 11204 6616 12348 6644
rect 11204 6604 11210 6616
rect 12342 6604 12348 6616
rect 12400 6604 12406 6656
rect 16850 6604 16856 6656
rect 16908 6644 16914 6656
rect 17681 6647 17739 6653
rect 17681 6644 17693 6647
rect 16908 6616 17693 6644
rect 16908 6604 16914 6616
rect 17681 6613 17693 6616
rect 17727 6613 17739 6647
rect 17681 6607 17739 6613
rect 19426 6604 19432 6656
rect 19484 6644 19490 6656
rect 19628 6644 19656 6743
rect 19720 6712 19748 6743
rect 19794 6740 19800 6792
rect 19852 6780 19858 6792
rect 20162 6780 20168 6792
rect 19852 6752 19897 6780
rect 19996 6752 20168 6780
rect 19852 6740 19858 6752
rect 19996 6712 20024 6752
rect 20162 6740 20168 6752
rect 20220 6740 20226 6792
rect 20364 6780 20392 6820
rect 20530 6808 20536 6820
rect 20588 6808 20594 6860
rect 21542 6808 21548 6860
rect 21600 6848 21606 6860
rect 22649 6851 22707 6857
rect 22649 6848 22661 6851
rect 21600 6820 22661 6848
rect 21600 6808 21606 6820
rect 22649 6817 22661 6820
rect 22695 6817 22707 6851
rect 22649 6811 22707 6817
rect 22370 6780 22376 6792
rect 20364 6752 22376 6780
rect 22370 6740 22376 6752
rect 22428 6740 22434 6792
rect 25777 6783 25835 6789
rect 25777 6749 25789 6783
rect 25823 6780 25835 6783
rect 26234 6780 26240 6792
rect 25823 6752 26240 6780
rect 25823 6749 25835 6752
rect 25777 6743 25835 6749
rect 26234 6740 26240 6752
rect 26292 6740 26298 6792
rect 26418 6780 26424 6792
rect 26379 6752 26424 6780
rect 26418 6740 26424 6752
rect 26476 6740 26482 6792
rect 26712 6789 26740 6888
rect 29822 6876 29828 6888
rect 29880 6916 29886 6928
rect 30190 6916 30196 6928
rect 29880 6888 30196 6916
rect 29880 6876 29886 6888
rect 30190 6876 30196 6888
rect 30248 6876 30254 6928
rect 26804 6820 29868 6848
rect 26804 6792 26832 6820
rect 26605 6783 26663 6789
rect 26605 6749 26617 6783
rect 26651 6749 26663 6783
rect 26605 6743 26663 6749
rect 26697 6783 26755 6789
rect 26697 6749 26709 6783
rect 26743 6749 26755 6783
rect 26697 6743 26755 6749
rect 19720 6684 20024 6712
rect 20073 6715 20131 6721
rect 20073 6681 20085 6715
rect 20119 6712 20131 6715
rect 20778 6715 20836 6721
rect 20778 6712 20790 6715
rect 20119 6684 20790 6712
rect 20119 6681 20131 6684
rect 20073 6675 20131 6681
rect 20778 6681 20790 6684
rect 20824 6681 20836 6715
rect 24949 6715 25007 6721
rect 24949 6712 24961 6715
rect 20778 6675 20836 6681
rect 23768 6684 24961 6712
rect 23768 6656 23796 6684
rect 24949 6681 24961 6684
rect 24995 6681 25007 6715
rect 25590 6712 25596 6724
rect 25503 6684 25596 6712
rect 24949 6675 25007 6681
rect 25590 6672 25596 6684
rect 25648 6672 25654 6724
rect 25961 6715 26019 6721
rect 25961 6681 25973 6715
rect 26007 6712 26019 6715
rect 26620 6712 26648 6743
rect 26786 6740 26792 6792
rect 26844 6780 26850 6792
rect 26844 6752 26937 6780
rect 26844 6740 26850 6752
rect 29270 6740 29276 6792
rect 29328 6780 29334 6792
rect 29549 6783 29607 6789
rect 29549 6780 29561 6783
rect 29328 6752 29561 6780
rect 29328 6740 29334 6752
rect 29549 6749 29561 6752
rect 29595 6749 29607 6783
rect 29549 6743 29607 6749
rect 29638 6740 29644 6792
rect 29696 6780 29702 6792
rect 29733 6783 29791 6789
rect 29733 6780 29745 6783
rect 29696 6752 29745 6780
rect 29696 6740 29702 6752
rect 29733 6749 29745 6752
rect 29779 6749 29791 6783
rect 29840 6780 29868 6820
rect 31570 6808 31576 6860
rect 31628 6848 31634 6860
rect 32033 6851 32091 6857
rect 32033 6848 32045 6851
rect 31628 6820 32045 6848
rect 31628 6808 31634 6820
rect 32033 6817 32045 6820
rect 32079 6817 32091 6851
rect 32033 6811 32091 6817
rect 36998 6808 37004 6860
rect 37056 6848 37062 6860
rect 39850 6848 39856 6860
rect 37056 6820 37596 6848
rect 39811 6820 39856 6848
rect 37056 6808 37062 6820
rect 32858 6780 32864 6792
rect 29840 6752 32864 6780
rect 29733 6743 29791 6749
rect 32858 6740 32864 6752
rect 32916 6740 32922 6792
rect 34606 6740 34612 6792
rect 34664 6780 34670 6792
rect 34701 6783 34759 6789
rect 34701 6780 34713 6783
rect 34664 6752 34713 6780
rect 34664 6740 34670 6752
rect 34701 6749 34713 6752
rect 34747 6749 34759 6783
rect 34701 6743 34759 6749
rect 35345 6783 35403 6789
rect 35345 6749 35357 6783
rect 35391 6780 35403 6783
rect 35391 6752 35848 6780
rect 35391 6749 35403 6752
rect 35345 6743 35403 6749
rect 29288 6712 29316 6740
rect 35820 6724 35848 6752
rect 37090 6740 37096 6792
rect 37148 6780 37154 6792
rect 37568 6789 37596 6820
rect 39850 6808 39856 6820
rect 39908 6808 39914 6860
rect 37369 6783 37427 6789
rect 37369 6780 37381 6783
rect 37148 6752 37381 6780
rect 37148 6740 37154 6752
rect 37369 6749 37381 6752
rect 37415 6749 37427 6783
rect 37369 6743 37427 6749
rect 37553 6783 37611 6789
rect 37553 6749 37565 6783
rect 37599 6749 37611 6783
rect 37553 6743 37611 6749
rect 37737 6783 37795 6789
rect 37737 6749 37749 6783
rect 37783 6749 37795 6783
rect 38562 6780 38568 6792
rect 38523 6752 38568 6780
rect 37737 6743 37795 6749
rect 32122 6712 32128 6724
rect 26007 6684 26648 6712
rect 26712 6684 29316 6712
rect 29840 6684 32128 6712
rect 26007 6681 26019 6684
rect 25961 6675 26019 6681
rect 19484 6616 19656 6644
rect 19484 6604 19490 6616
rect 19978 6604 19984 6656
rect 20036 6644 20042 6656
rect 21913 6647 21971 6653
rect 21913 6644 21925 6647
rect 20036 6616 21925 6644
rect 20036 6604 20042 6616
rect 21913 6613 21925 6616
rect 21959 6613 21971 6647
rect 23750 6644 23756 6656
rect 23711 6616 23756 6644
rect 21913 6607 21971 6613
rect 23750 6604 23756 6616
rect 23808 6604 23814 6656
rect 25038 6604 25044 6656
rect 25096 6644 25102 6656
rect 25608 6644 25636 6672
rect 26712 6644 26740 6684
rect 27062 6644 27068 6656
rect 25096 6616 25141 6644
rect 25608 6616 26740 6644
rect 27023 6616 27068 6644
rect 25096 6604 25102 6616
rect 27062 6604 27068 6616
rect 27120 6604 27126 6656
rect 28902 6644 28908 6656
rect 28863 6616 28908 6644
rect 28902 6604 28908 6616
rect 28960 6644 28966 6656
rect 29546 6644 29552 6656
rect 28960 6616 29552 6644
rect 28960 6604 28966 6616
rect 29546 6604 29552 6616
rect 29604 6644 29610 6656
rect 29840 6644 29868 6684
rect 32122 6672 32128 6684
rect 32180 6672 32186 6724
rect 32300 6715 32358 6721
rect 32300 6681 32312 6715
rect 32346 6712 32358 6715
rect 33594 6712 33600 6724
rect 32346 6684 33600 6712
rect 32346 6681 32358 6684
rect 32300 6675 32358 6681
rect 33594 6672 33600 6684
rect 33652 6672 33658 6724
rect 35158 6672 35164 6724
rect 35216 6712 35222 6724
rect 35590 6715 35648 6721
rect 35590 6712 35602 6715
rect 35216 6684 35602 6712
rect 35216 6672 35222 6684
rect 35590 6681 35602 6684
rect 35636 6681 35648 6715
rect 35590 6675 35648 6681
rect 35802 6672 35808 6724
rect 35860 6672 35866 6724
rect 37461 6715 37519 6721
rect 37461 6681 37473 6715
rect 37507 6681 37519 6715
rect 37752 6712 37780 6743
rect 38562 6740 38568 6752
rect 38620 6740 38626 6792
rect 39942 6740 39948 6792
rect 40000 6780 40006 6792
rect 40109 6783 40167 6789
rect 40109 6780 40121 6783
rect 40000 6752 40121 6780
rect 40000 6740 40006 6752
rect 40109 6749 40121 6752
rect 40155 6749 40167 6783
rect 40109 6743 40167 6749
rect 38381 6715 38439 6721
rect 38381 6712 38393 6715
rect 37752 6684 38393 6712
rect 37461 6675 37519 6681
rect 38381 6681 38393 6684
rect 38427 6681 38439 6715
rect 38381 6675 38439 6681
rect 29604 6616 29868 6644
rect 29604 6604 29610 6616
rect 29914 6604 29920 6656
rect 29972 6644 29978 6656
rect 32140 6644 32168 6672
rect 34606 6644 34612 6656
rect 29972 6616 30017 6644
rect 32140 6616 34612 6644
rect 29972 6604 29978 6616
rect 34606 6604 34612 6616
rect 34664 6604 34670 6656
rect 34698 6604 34704 6656
rect 34756 6644 34762 6656
rect 34885 6647 34943 6653
rect 34885 6644 34897 6647
rect 34756 6616 34897 6644
rect 34756 6604 34762 6616
rect 34885 6613 34897 6616
rect 34931 6613 34943 6647
rect 34885 6607 34943 6613
rect 36814 6604 36820 6656
rect 36872 6644 36878 6656
rect 37185 6647 37243 6653
rect 37185 6644 37197 6647
rect 36872 6616 37197 6644
rect 36872 6604 36878 6616
rect 37185 6613 37197 6616
rect 37231 6613 37243 6647
rect 37476 6644 37504 6675
rect 37642 6644 37648 6656
rect 37476 6616 37648 6644
rect 37185 6607 37243 6613
rect 37642 6604 37648 6616
rect 37700 6604 37706 6656
rect 38396 6644 38424 6675
rect 41233 6647 41291 6653
rect 41233 6644 41245 6647
rect 38396 6616 41245 6644
rect 41233 6613 41245 6616
rect 41279 6613 41291 6647
rect 41233 6607 41291 6613
rect 1104 6554 68816 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 68816 6554
rect 1104 6480 68816 6502
rect 4062 6440 4068 6452
rect 2746 6412 4068 6440
rect 2314 6332 2320 6384
rect 2372 6372 2378 6384
rect 2746 6372 2774 6412
rect 4062 6400 4068 6412
rect 4120 6400 4126 6452
rect 4157 6443 4215 6449
rect 4157 6409 4169 6443
rect 4203 6440 4215 6443
rect 5261 6443 5319 6449
rect 5261 6440 5273 6443
rect 4203 6412 5273 6440
rect 4203 6409 4215 6412
rect 4157 6403 4215 6409
rect 5261 6409 5273 6412
rect 5307 6440 5319 6443
rect 5810 6440 5816 6452
rect 5307 6412 5816 6440
rect 5307 6409 5319 6412
rect 5261 6403 5319 6409
rect 5810 6400 5816 6412
rect 5868 6400 5874 6452
rect 5902 6400 5908 6452
rect 5960 6440 5966 6452
rect 7190 6440 7196 6452
rect 5960 6412 7196 6440
rect 5960 6400 5966 6412
rect 7190 6400 7196 6412
rect 7248 6400 7254 6452
rect 8389 6443 8447 6449
rect 8389 6409 8401 6443
rect 8435 6440 8447 6443
rect 9214 6440 9220 6452
rect 8435 6412 9220 6440
rect 8435 6409 8447 6412
rect 8389 6403 8447 6409
rect 9214 6400 9220 6412
rect 9272 6400 9278 6452
rect 9490 6400 9496 6452
rect 9548 6440 9554 6452
rect 10686 6440 10692 6452
rect 9548 6412 10692 6440
rect 9548 6400 9554 6412
rect 10686 6400 10692 6412
rect 10744 6400 10750 6452
rect 16298 6400 16304 6452
rect 16356 6440 16362 6452
rect 18046 6440 18052 6452
rect 16356 6412 18052 6440
rect 16356 6400 16362 6412
rect 18046 6400 18052 6412
rect 18104 6440 18110 6452
rect 18325 6443 18383 6449
rect 18325 6440 18337 6443
rect 18104 6412 18337 6440
rect 18104 6400 18110 6412
rect 18325 6409 18337 6412
rect 18371 6409 18383 6443
rect 18325 6403 18383 6409
rect 19426 6400 19432 6452
rect 19484 6440 19490 6452
rect 19613 6443 19671 6449
rect 19613 6440 19625 6443
rect 19484 6412 19625 6440
rect 19484 6400 19490 6412
rect 19613 6409 19625 6412
rect 19659 6409 19671 6443
rect 23658 6440 23664 6452
rect 23619 6412 23664 6440
rect 19613 6403 19671 6409
rect 23658 6400 23664 6412
rect 23716 6400 23722 6452
rect 25038 6400 25044 6452
rect 25096 6440 25102 6452
rect 26421 6443 26479 6449
rect 26421 6440 26433 6443
rect 25096 6412 26433 6440
rect 25096 6400 25102 6412
rect 26421 6409 26433 6412
rect 26467 6440 26479 6443
rect 26786 6440 26792 6452
rect 26467 6412 26792 6440
rect 26467 6409 26479 6412
rect 26421 6403 26479 6409
rect 26786 6400 26792 6412
rect 26844 6400 26850 6452
rect 26896 6412 29592 6440
rect 2958 6372 2964 6384
rect 2372 6344 2774 6372
rect 2871 6344 2964 6372
rect 2372 6332 2378 6344
rect 2958 6332 2964 6344
rect 3016 6372 3022 6384
rect 4614 6372 4620 6384
rect 3016 6344 4620 6372
rect 3016 6332 3022 6344
rect 4614 6332 4620 6344
rect 4672 6332 4678 6384
rect 5169 6375 5227 6381
rect 5169 6341 5181 6375
rect 5215 6372 5227 6375
rect 5442 6372 5448 6384
rect 5215 6344 5448 6372
rect 5215 6341 5227 6344
rect 5169 6335 5227 6341
rect 5442 6332 5448 6344
rect 5500 6372 5506 6384
rect 5718 6372 5724 6384
rect 5500 6344 5724 6372
rect 5500 6332 5506 6344
rect 5718 6332 5724 6344
rect 5776 6332 5782 6384
rect 6454 6332 6460 6384
rect 6512 6372 6518 6384
rect 8294 6372 8300 6384
rect 6512 6344 8300 6372
rect 6512 6332 6518 6344
rect 1762 6304 1768 6316
rect 1723 6276 1768 6304
rect 1762 6264 1768 6276
rect 1820 6264 1826 6316
rect 1857 6307 1915 6313
rect 1857 6273 1869 6307
rect 1903 6304 1915 6307
rect 2777 6307 2835 6313
rect 1903 6276 2728 6304
rect 1903 6273 1915 6276
rect 1857 6267 1915 6273
rect 1946 6060 1952 6112
rect 2004 6100 2010 6112
rect 2041 6103 2099 6109
rect 2041 6100 2053 6103
rect 2004 6072 2053 6100
rect 2004 6060 2010 6072
rect 2041 6069 2053 6072
rect 2087 6069 2099 6103
rect 2700 6100 2728 6276
rect 2777 6273 2789 6307
rect 2823 6304 2835 6307
rect 2976 6304 3004 6332
rect 3050 6313 3056 6316
rect 2823 6276 3004 6304
rect 2823 6273 2835 6276
rect 2777 6267 2835 6273
rect 3044 6267 3056 6313
rect 3108 6304 3114 6316
rect 3108 6276 3144 6304
rect 3050 6264 3056 6267
rect 3108 6264 3114 6276
rect 6914 6264 6920 6316
rect 6972 6304 6978 6316
rect 7300 6313 7328 6344
rect 8294 6332 8300 6344
rect 8352 6372 8358 6384
rect 9122 6372 9128 6384
rect 8352 6344 9128 6372
rect 8352 6332 8358 6344
rect 9122 6332 9128 6344
rect 9180 6332 9186 6384
rect 11054 6332 11060 6384
rect 11112 6372 11118 6384
rect 11762 6375 11820 6381
rect 11762 6372 11774 6375
rect 11112 6344 11774 6372
rect 11112 6332 11118 6344
rect 11762 6341 11774 6344
rect 11808 6341 11820 6375
rect 12434 6372 12440 6384
rect 11762 6335 11820 6341
rect 11900 6344 12440 6372
rect 7009 6307 7067 6313
rect 7009 6304 7021 6307
rect 6972 6276 7021 6304
rect 6972 6264 6978 6276
rect 7009 6273 7021 6276
rect 7055 6273 7067 6307
rect 7009 6267 7067 6273
rect 7285 6307 7343 6313
rect 7285 6273 7297 6307
rect 7331 6273 7343 6307
rect 7285 6267 7343 6273
rect 7929 6307 7987 6313
rect 7929 6273 7941 6307
rect 7975 6273 7987 6307
rect 7929 6267 7987 6273
rect 4062 6196 4068 6248
rect 4120 6236 4126 6248
rect 5353 6239 5411 6245
rect 5353 6236 5365 6239
rect 4120 6208 5365 6236
rect 4120 6196 4126 6208
rect 5353 6205 5365 6208
rect 5399 6236 5411 6239
rect 6638 6236 6644 6248
rect 5399 6208 6644 6236
rect 5399 6205 5411 6208
rect 5353 6199 5411 6205
rect 6638 6196 6644 6208
rect 6696 6196 6702 6248
rect 6822 6196 6828 6248
rect 6880 6196 6886 6248
rect 7650 6196 7656 6248
rect 7708 6236 7714 6248
rect 7944 6236 7972 6267
rect 8018 6264 8024 6316
rect 8076 6304 8082 6316
rect 8205 6307 8263 6313
rect 8076 6276 8121 6304
rect 8076 6264 8082 6276
rect 8205 6273 8217 6307
rect 8251 6304 8263 6307
rect 9306 6304 9312 6316
rect 8251 6276 9312 6304
rect 8251 6273 8263 6276
rect 8205 6267 8263 6273
rect 9306 6264 9312 6276
rect 9364 6264 9370 6316
rect 9861 6307 9919 6313
rect 9861 6273 9873 6307
rect 9907 6304 9919 6307
rect 10134 6304 10140 6316
rect 9907 6276 10140 6304
rect 9907 6273 9919 6276
rect 9861 6267 9919 6273
rect 10134 6264 10140 6276
rect 10192 6264 10198 6316
rect 10965 6307 11023 6313
rect 10965 6273 10977 6307
rect 11011 6304 11023 6307
rect 11900 6304 11928 6344
rect 12434 6332 12440 6344
rect 12492 6332 12498 6384
rect 12618 6332 12624 6384
rect 12676 6372 12682 6384
rect 17034 6372 17040 6384
rect 12676 6344 15608 6372
rect 12676 6332 12682 6344
rect 11011 6276 11928 6304
rect 13357 6307 13415 6313
rect 11011 6273 11023 6276
rect 10965 6267 11023 6273
rect 13357 6273 13369 6307
rect 13403 6304 13415 6307
rect 13446 6304 13452 6316
rect 13403 6276 13452 6304
rect 13403 6273 13415 6276
rect 13357 6267 13415 6273
rect 13446 6264 13452 6276
rect 13504 6264 13510 6316
rect 15580 6313 15608 6344
rect 15764 6344 16896 6372
rect 16995 6344 17040 6372
rect 15764 6313 15792 6344
rect 13624 6307 13682 6313
rect 13624 6273 13636 6307
rect 13670 6304 13682 6307
rect 15197 6307 15255 6313
rect 15197 6304 15209 6307
rect 13670 6276 15209 6304
rect 13670 6273 13682 6276
rect 13624 6267 13682 6273
rect 15197 6273 15209 6276
rect 15243 6273 15255 6307
rect 15197 6267 15255 6273
rect 15381 6307 15439 6313
rect 15381 6273 15393 6307
rect 15427 6273 15439 6307
rect 15381 6267 15439 6273
rect 15565 6307 15623 6313
rect 15565 6273 15577 6307
rect 15611 6273 15623 6307
rect 15565 6267 15623 6273
rect 15749 6307 15807 6313
rect 15749 6273 15761 6307
rect 15795 6273 15807 6307
rect 15930 6304 15936 6316
rect 15891 6276 15936 6304
rect 15749 6267 15807 6273
rect 9582 6236 9588 6248
rect 7708 6208 9588 6236
rect 7708 6196 7714 6208
rect 9582 6196 9588 6208
rect 9640 6196 9646 6248
rect 9950 6196 9956 6248
rect 10008 6236 10014 6248
rect 10870 6236 10876 6248
rect 10008 6208 10876 6236
rect 10008 6196 10014 6208
rect 10870 6196 10876 6208
rect 10928 6236 10934 6248
rect 11517 6239 11575 6245
rect 11517 6236 11529 6239
rect 10928 6208 11529 6236
rect 10928 6196 10934 6208
rect 11517 6205 11529 6208
rect 11563 6205 11575 6239
rect 15396 6236 15424 6267
rect 15930 6264 15936 6276
rect 15988 6264 15994 6316
rect 16868 6304 16896 6344
rect 17034 6332 17040 6344
rect 17092 6332 17098 6384
rect 19245 6375 19303 6381
rect 19245 6341 19257 6375
rect 19291 6372 19303 6375
rect 23382 6372 23388 6384
rect 19291 6344 20760 6372
rect 19291 6341 19303 6344
rect 19245 6335 19303 6341
rect 20732 6316 20760 6344
rect 22296 6344 23388 6372
rect 19150 6304 19156 6316
rect 16868 6276 19156 6304
rect 19150 6264 19156 6276
rect 19208 6264 19214 6316
rect 19429 6307 19487 6313
rect 19429 6273 19441 6307
rect 19475 6304 19487 6307
rect 19978 6304 19984 6316
rect 19475 6276 19984 6304
rect 19475 6273 19487 6276
rect 19429 6267 19487 6273
rect 19978 6264 19984 6276
rect 20036 6264 20042 6316
rect 20714 6304 20720 6316
rect 20675 6276 20720 6304
rect 20714 6264 20720 6276
rect 20772 6264 20778 6316
rect 22094 6264 22100 6316
rect 22152 6304 22158 6316
rect 22296 6313 22324 6344
rect 23382 6332 23388 6344
rect 23440 6372 23446 6384
rect 24121 6375 24179 6381
rect 24121 6372 24133 6375
rect 23440 6344 24133 6372
rect 23440 6332 23446 6344
rect 24121 6341 24133 6344
rect 24167 6341 24179 6375
rect 24121 6335 24179 6341
rect 26326 6332 26332 6384
rect 26384 6372 26390 6384
rect 26896 6372 26924 6412
rect 26384 6344 26924 6372
rect 26384 6332 26390 6344
rect 27062 6332 27068 6384
rect 27120 6372 27126 6384
rect 28178 6375 28236 6381
rect 28178 6372 28190 6375
rect 27120 6344 28190 6372
rect 27120 6332 27126 6344
rect 28178 6341 28190 6344
rect 28224 6341 28236 6375
rect 29564 6372 29592 6412
rect 29638 6400 29644 6452
rect 29696 6440 29702 6452
rect 30193 6443 30251 6449
rect 30193 6440 30205 6443
rect 29696 6412 30205 6440
rect 29696 6400 29702 6412
rect 30193 6409 30205 6412
rect 30239 6409 30251 6443
rect 33594 6440 33600 6452
rect 33555 6412 33600 6440
rect 30193 6403 30251 6409
rect 33594 6400 33600 6412
rect 33652 6400 33658 6452
rect 33686 6400 33692 6452
rect 33744 6440 33750 6452
rect 35158 6440 35164 6452
rect 33744 6412 34008 6440
rect 35119 6412 35164 6440
rect 33744 6400 33750 6412
rect 29730 6372 29736 6384
rect 29564 6344 29736 6372
rect 28178 6335 28236 6341
rect 29730 6332 29736 6344
rect 29788 6372 29794 6384
rect 33137 6375 33195 6381
rect 33137 6372 33149 6375
rect 29788 6344 33149 6372
rect 29788 6332 29794 6344
rect 33137 6341 33149 6344
rect 33183 6372 33195 6375
rect 33980 6372 34008 6412
rect 35158 6400 35164 6412
rect 35216 6400 35222 6452
rect 35986 6440 35992 6452
rect 35544 6412 35992 6440
rect 35544 6372 35572 6412
rect 35986 6400 35992 6412
rect 36044 6400 36050 6452
rect 38562 6440 38568 6452
rect 36648 6412 38568 6440
rect 36265 6375 36323 6381
rect 36265 6372 36277 6375
rect 33183 6344 33916 6372
rect 33183 6341 33195 6344
rect 33137 6335 33195 6341
rect 33888 6316 33916 6344
rect 33980 6344 35572 6372
rect 22281 6307 22339 6313
rect 22281 6304 22293 6307
rect 22152 6276 22293 6304
rect 22152 6264 22158 6276
rect 22281 6273 22293 6276
rect 22327 6273 22339 6307
rect 22281 6267 22339 6273
rect 22548 6307 22606 6313
rect 22548 6273 22560 6307
rect 22594 6304 22606 6307
rect 23842 6304 23848 6316
rect 22594 6276 23848 6304
rect 22594 6273 22606 6276
rect 22548 6267 22606 6273
rect 23842 6264 23848 6276
rect 23900 6264 23906 6316
rect 25869 6307 25927 6313
rect 25869 6273 25881 6307
rect 25915 6304 25927 6307
rect 27614 6304 27620 6316
rect 25915 6276 27620 6304
rect 25915 6273 25927 6276
rect 25869 6267 25927 6273
rect 27614 6264 27620 6276
rect 27672 6264 27678 6316
rect 29086 6304 29092 6316
rect 29047 6276 29092 6304
rect 29086 6264 29092 6276
rect 29144 6264 29150 6316
rect 29252 6307 29310 6313
rect 29252 6304 29264 6307
rect 29196 6276 29264 6304
rect 11517 6199 11575 6205
rect 14752 6208 15424 6236
rect 4801 6171 4859 6177
rect 4801 6168 4813 6171
rect 3804 6140 4813 6168
rect 3804 6100 3832 6140
rect 4801 6137 4813 6140
rect 4847 6137 4859 6171
rect 6840 6168 6868 6196
rect 10502 6168 10508 6180
rect 6840 6140 10508 6168
rect 4801 6131 4859 6137
rect 10502 6128 10508 6140
rect 10560 6128 10566 6180
rect 14752 6177 14780 6208
rect 15212 6180 15240 6208
rect 15654 6196 15660 6248
rect 15712 6236 15718 6248
rect 15948 6236 15976 6264
rect 17678 6236 17684 6248
rect 15712 6208 15757 6236
rect 15948 6208 17684 6236
rect 15712 6196 15718 6208
rect 17678 6196 17684 6208
rect 17736 6196 17742 6248
rect 28445 6239 28503 6245
rect 28445 6205 28457 6239
rect 28491 6236 28503 6239
rect 28994 6236 29000 6248
rect 28491 6208 29000 6236
rect 28491 6205 28503 6208
rect 28445 6199 28503 6205
rect 28994 6196 29000 6208
rect 29052 6196 29058 6248
rect 14737 6171 14795 6177
rect 14737 6137 14749 6171
rect 14783 6137 14795 6171
rect 14737 6131 14795 6137
rect 15194 6128 15200 6180
rect 15252 6128 15258 6180
rect 26234 6128 26240 6180
rect 26292 6168 26298 6180
rect 27065 6171 27123 6177
rect 27065 6168 27077 6171
rect 26292 6140 27077 6168
rect 26292 6128 26298 6140
rect 27065 6137 27077 6140
rect 27111 6137 27123 6171
rect 29196 6168 29224 6276
rect 29252 6273 29264 6276
rect 29298 6273 29310 6307
rect 29252 6267 29310 6273
rect 29365 6307 29423 6313
rect 29365 6273 29377 6307
rect 29411 6273 29423 6307
rect 29365 6267 29423 6273
rect 29457 6307 29515 6313
rect 29546 6307 29552 6316
rect 29457 6273 29469 6307
rect 29503 6279 29552 6307
rect 29503 6273 29515 6279
rect 29457 6267 29515 6273
rect 29380 6236 29408 6267
rect 29546 6264 29552 6279
rect 29604 6264 29610 6316
rect 30466 6264 30472 6316
rect 30524 6304 30530 6316
rect 31306 6307 31364 6313
rect 31306 6304 31318 6307
rect 30524 6276 31318 6304
rect 30524 6264 30530 6276
rect 31306 6273 31318 6276
rect 31352 6273 31364 6307
rect 33870 6304 33876 6316
rect 33783 6276 33876 6304
rect 31306 6267 31364 6273
rect 33870 6264 33876 6276
rect 33928 6264 33934 6316
rect 33980 6313 34008 6344
rect 33965 6307 34023 6313
rect 33965 6273 33977 6307
rect 34011 6273 34023 6307
rect 33965 6267 34023 6273
rect 34054 6264 34060 6316
rect 34112 6304 34118 6316
rect 34112 6276 34157 6304
rect 34112 6264 34118 6276
rect 34238 6264 34244 6316
rect 34296 6304 34302 6316
rect 34296 6276 34341 6304
rect 34296 6264 34302 6276
rect 34606 6264 34612 6316
rect 34664 6304 34670 6316
rect 35434 6304 35440 6316
rect 34664 6276 35440 6304
rect 34664 6264 34670 6276
rect 35434 6264 35440 6276
rect 35492 6264 35498 6316
rect 35544 6313 35572 6344
rect 35636 6344 36277 6372
rect 35636 6313 35664 6344
rect 36265 6341 36277 6344
rect 36311 6341 36323 6375
rect 36265 6335 36323 6341
rect 36354 6332 36360 6384
rect 36412 6372 36418 6384
rect 36648 6381 36676 6412
rect 38562 6400 38568 6412
rect 38620 6400 38626 6452
rect 36449 6375 36507 6381
rect 36449 6372 36461 6375
rect 36412 6344 36461 6372
rect 36412 6332 36418 6344
rect 36449 6341 36461 6344
rect 36495 6341 36507 6375
rect 36449 6335 36507 6341
rect 36633 6375 36691 6381
rect 36633 6341 36645 6375
rect 36679 6341 36691 6375
rect 36633 6335 36691 6341
rect 37461 6375 37519 6381
rect 37461 6341 37473 6375
rect 37507 6372 37519 6375
rect 37642 6372 37648 6384
rect 37507 6344 37648 6372
rect 37507 6341 37519 6344
rect 37461 6335 37519 6341
rect 37642 6332 37648 6344
rect 37700 6372 37706 6384
rect 38654 6372 38660 6384
rect 37700 6344 38660 6372
rect 37700 6332 37706 6344
rect 38654 6332 38660 6344
rect 38712 6332 38718 6384
rect 35529 6307 35587 6313
rect 35529 6273 35541 6307
rect 35575 6273 35587 6307
rect 35529 6267 35587 6273
rect 35621 6307 35679 6313
rect 35621 6273 35633 6307
rect 35667 6273 35679 6307
rect 35621 6267 35679 6273
rect 35805 6307 35863 6313
rect 35805 6273 35817 6307
rect 35851 6273 35863 6307
rect 35805 6267 35863 6273
rect 37277 6307 37335 6313
rect 37277 6273 37289 6307
rect 37323 6304 37335 6307
rect 37366 6304 37372 6316
rect 37323 6276 37372 6304
rect 37323 6273 37335 6276
rect 37277 6267 37335 6273
rect 30190 6236 30196 6248
rect 29380 6208 30196 6236
rect 30190 6196 30196 6208
rect 30248 6196 30254 6248
rect 31570 6236 31576 6248
rect 31531 6208 31576 6236
rect 31570 6196 31576 6208
rect 31628 6196 31634 6248
rect 29270 6168 29276 6180
rect 29196 6140 29276 6168
rect 27065 6131 27123 6137
rect 29270 6128 29276 6140
rect 29328 6128 29334 6180
rect 29733 6171 29791 6177
rect 29733 6137 29745 6171
rect 29779 6168 29791 6171
rect 30558 6168 30564 6180
rect 29779 6140 30564 6168
rect 29779 6137 29791 6140
rect 29733 6131 29791 6137
rect 30558 6128 30564 6140
rect 30616 6128 30622 6180
rect 34256 6168 34284 6264
rect 35820 6168 35848 6267
rect 37366 6264 37372 6276
rect 37424 6264 37430 6316
rect 38102 6304 38108 6316
rect 38063 6276 38108 6304
rect 38102 6264 38108 6276
rect 38160 6264 38166 6316
rect 38289 6307 38347 6313
rect 38289 6273 38301 6307
rect 38335 6273 38347 6307
rect 38289 6267 38347 6273
rect 38381 6307 38439 6313
rect 38381 6273 38393 6307
rect 38427 6273 38439 6307
rect 38381 6267 38439 6273
rect 37645 6239 37703 6245
rect 37645 6205 37657 6239
rect 37691 6236 37703 6239
rect 38304 6236 38332 6267
rect 37691 6208 38332 6236
rect 37691 6205 37703 6208
rect 37645 6199 37703 6205
rect 34256 6140 35848 6168
rect 37182 6128 37188 6180
rect 37240 6168 37246 6180
rect 38396 6168 38424 6267
rect 38470 6264 38476 6316
rect 38528 6304 38534 6316
rect 38528 6276 38573 6304
rect 38528 6264 38534 6276
rect 67634 6168 67640 6180
rect 37240 6140 38424 6168
rect 67595 6140 67640 6168
rect 37240 6128 37246 6140
rect 67634 6128 67640 6140
rect 67692 6128 67698 6180
rect 2700 6072 3832 6100
rect 2041 6063 2099 6069
rect 8110 6060 8116 6112
rect 8168 6100 8174 6112
rect 10594 6100 10600 6112
rect 8168 6072 10600 6100
rect 8168 6060 8174 6072
rect 10594 6060 10600 6072
rect 10652 6060 10658 6112
rect 10781 6103 10839 6109
rect 10781 6069 10793 6103
rect 10827 6100 10839 6103
rect 11330 6100 11336 6112
rect 10827 6072 11336 6100
rect 10827 6069 10839 6072
rect 10781 6063 10839 6069
rect 11330 6060 11336 6072
rect 11388 6060 11394 6112
rect 11698 6060 11704 6112
rect 11756 6100 11762 6112
rect 12897 6103 12955 6109
rect 12897 6100 12909 6103
rect 11756 6072 12909 6100
rect 11756 6060 11762 6072
rect 12897 6069 12909 6072
rect 12943 6100 12955 6103
rect 14550 6100 14556 6112
rect 12943 6072 14556 6100
rect 12943 6069 12955 6072
rect 12897 6063 12955 6069
rect 14550 6060 14556 6072
rect 14608 6060 14614 6112
rect 20070 6100 20076 6112
rect 20031 6072 20076 6100
rect 20070 6060 20076 6072
rect 20128 6060 20134 6112
rect 20901 6103 20959 6109
rect 20901 6069 20913 6103
rect 20947 6100 20959 6103
rect 23014 6100 23020 6112
rect 20947 6072 23020 6100
rect 20947 6069 20959 6072
rect 20901 6063 20959 6069
rect 23014 6060 23020 6072
rect 23072 6060 23078 6112
rect 28258 6060 28264 6112
rect 28316 6100 28322 6112
rect 30282 6100 30288 6112
rect 28316 6072 30288 6100
rect 28316 6060 28322 6072
rect 30282 6060 30288 6072
rect 30340 6100 30346 6112
rect 30926 6100 30932 6112
rect 30340 6072 30932 6100
rect 30340 6060 30346 6072
rect 30926 6060 30932 6072
rect 30984 6060 30990 6112
rect 38746 6100 38752 6112
rect 38707 6072 38752 6100
rect 38746 6060 38752 6072
rect 38804 6060 38810 6112
rect 1104 6010 68816 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 65654 6010
rect 65706 5958 65718 6010
rect 65770 5958 65782 6010
rect 65834 5958 65846 6010
rect 65898 5958 65910 6010
rect 65962 5958 68816 6010
rect 1104 5936 68816 5958
rect 2133 5899 2191 5905
rect 2133 5865 2145 5899
rect 2179 5896 2191 5899
rect 3050 5896 3056 5908
rect 2179 5868 3056 5896
rect 2179 5865 2191 5868
rect 2133 5859 2191 5865
rect 3050 5856 3056 5868
rect 3108 5856 3114 5908
rect 3234 5896 3240 5908
rect 3195 5868 3240 5896
rect 3234 5856 3240 5868
rect 3292 5856 3298 5908
rect 5445 5899 5503 5905
rect 5445 5865 5457 5899
rect 5491 5896 5503 5899
rect 5534 5896 5540 5908
rect 5491 5868 5540 5896
rect 5491 5865 5503 5868
rect 5445 5859 5503 5865
rect 5534 5856 5540 5868
rect 5592 5896 5598 5908
rect 6730 5896 6736 5908
rect 5592 5868 6736 5896
rect 5592 5856 5598 5868
rect 6730 5856 6736 5868
rect 6788 5856 6794 5908
rect 9582 5856 9588 5908
rect 9640 5896 9646 5908
rect 15654 5896 15660 5908
rect 9640 5868 15148 5896
rect 15615 5868 15660 5896
rect 9640 5856 9646 5868
rect 1489 5831 1547 5837
rect 1489 5797 1501 5831
rect 1535 5828 1547 5831
rect 5258 5828 5264 5840
rect 1535 5800 5264 5828
rect 1535 5797 1547 5800
rect 1489 5791 1547 5797
rect 5258 5788 5264 5800
rect 5316 5788 5322 5840
rect 6089 5831 6147 5837
rect 6089 5797 6101 5831
rect 6135 5828 6147 5831
rect 9214 5828 9220 5840
rect 6135 5800 9220 5828
rect 6135 5797 6147 5800
rect 6089 5791 6147 5797
rect 9214 5788 9220 5800
rect 9272 5788 9278 5840
rect 13630 5788 13636 5840
rect 13688 5828 13694 5840
rect 13814 5828 13820 5840
rect 13688 5800 13820 5828
rect 13688 5788 13694 5800
rect 13814 5788 13820 5800
rect 13872 5788 13878 5840
rect 4893 5763 4951 5769
rect 4893 5729 4905 5763
rect 4939 5760 4951 5763
rect 8202 5760 8208 5772
rect 4939 5732 8208 5760
rect 4939 5729 4951 5732
rect 4893 5723 4951 5729
rect 8202 5720 8208 5732
rect 8260 5720 8266 5772
rect 9858 5720 9864 5772
rect 9916 5760 9922 5772
rect 15120 5760 15148 5868
rect 15654 5856 15660 5868
rect 15712 5856 15718 5908
rect 16666 5896 16672 5908
rect 16627 5868 16672 5896
rect 16666 5856 16672 5868
rect 16724 5856 16730 5908
rect 17862 5896 17868 5908
rect 17823 5868 17868 5896
rect 17862 5856 17868 5868
rect 17920 5856 17926 5908
rect 18874 5856 18880 5908
rect 18932 5896 18938 5908
rect 23474 5896 23480 5908
rect 18932 5868 23336 5896
rect 23435 5868 23480 5896
rect 18932 5856 18938 5868
rect 15197 5831 15255 5837
rect 15197 5797 15209 5831
rect 15243 5828 15255 5831
rect 17770 5828 17776 5840
rect 15243 5800 17776 5828
rect 15243 5797 15255 5800
rect 15197 5791 15255 5797
rect 17770 5788 17776 5800
rect 17828 5788 17834 5840
rect 23308 5828 23336 5868
rect 23474 5856 23480 5868
rect 23532 5856 23538 5908
rect 25685 5899 25743 5905
rect 25685 5865 25697 5899
rect 25731 5896 25743 5899
rect 26326 5896 26332 5908
rect 25731 5868 26332 5896
rect 25731 5865 25743 5868
rect 25685 5859 25743 5865
rect 26326 5856 26332 5868
rect 26384 5856 26390 5908
rect 26513 5899 26571 5905
rect 26513 5865 26525 5899
rect 26559 5896 26571 5899
rect 28902 5896 28908 5908
rect 26559 5868 28908 5896
rect 26559 5865 26571 5868
rect 26513 5859 26571 5865
rect 28902 5856 28908 5868
rect 28960 5856 28966 5908
rect 28997 5899 29055 5905
rect 28997 5865 29009 5899
rect 29043 5896 29055 5899
rect 29270 5896 29276 5908
rect 29043 5868 29276 5896
rect 29043 5865 29055 5868
rect 28997 5859 29055 5865
rect 29270 5856 29276 5868
rect 29328 5856 29334 5908
rect 30466 5896 30472 5908
rect 30427 5868 30472 5896
rect 30466 5856 30472 5868
rect 30524 5856 30530 5908
rect 35434 5856 35440 5908
rect 35492 5896 35498 5908
rect 35986 5896 35992 5908
rect 35492 5868 35992 5896
rect 35492 5856 35498 5868
rect 35986 5856 35992 5868
rect 36044 5856 36050 5908
rect 38289 5899 38347 5905
rect 38289 5865 38301 5899
rect 38335 5896 38347 5899
rect 38470 5896 38476 5908
rect 38335 5868 38476 5896
rect 38335 5865 38347 5868
rect 38289 5859 38347 5865
rect 38470 5856 38476 5868
rect 38528 5856 38534 5908
rect 26418 5828 26424 5840
rect 23308 5800 26424 5828
rect 26418 5788 26424 5800
rect 26476 5828 26482 5840
rect 27617 5831 27675 5837
rect 27617 5828 27629 5831
rect 26476 5800 27629 5828
rect 26476 5788 26482 5800
rect 27617 5797 27629 5800
rect 27663 5797 27675 5831
rect 30926 5828 30932 5840
rect 30887 5800 30932 5828
rect 27617 5791 27675 5797
rect 30926 5788 30932 5800
rect 30984 5828 30990 5840
rect 36541 5831 36599 5837
rect 36541 5828 36553 5831
rect 30984 5800 36553 5828
rect 30984 5788 30990 5800
rect 36541 5797 36553 5800
rect 36587 5828 36599 5831
rect 36587 5800 37504 5828
rect 36587 5797 36599 5800
rect 36541 5791 36599 5797
rect 17037 5763 17095 5769
rect 9916 5732 12296 5760
rect 15120 5732 16160 5760
rect 9916 5720 9922 5732
rect 1946 5692 1952 5704
rect 1907 5664 1952 5692
rect 1946 5652 1952 5664
rect 2004 5652 2010 5704
rect 3973 5695 4031 5701
rect 3973 5661 3985 5695
rect 4019 5692 4031 5695
rect 5810 5692 5816 5704
rect 4019 5664 5816 5692
rect 4019 5661 4031 5664
rect 3973 5655 4031 5661
rect 5810 5652 5816 5664
rect 5868 5652 5874 5704
rect 5905 5695 5963 5701
rect 5905 5661 5917 5695
rect 5951 5692 5963 5695
rect 7742 5692 7748 5704
rect 5951 5664 7748 5692
rect 5951 5661 5963 5664
rect 5905 5655 5963 5661
rect 7742 5652 7748 5664
rect 7800 5652 7806 5704
rect 7834 5652 7840 5704
rect 7892 5692 7898 5704
rect 8113 5695 8171 5701
rect 7892 5664 7937 5692
rect 7892 5652 7898 5664
rect 8113 5661 8125 5695
rect 8159 5661 8171 5695
rect 8113 5655 8171 5661
rect 9033 5695 9091 5701
rect 9033 5661 9045 5695
rect 9079 5692 9091 5695
rect 9306 5692 9312 5704
rect 9079 5664 9312 5692
rect 9079 5661 9091 5664
rect 9033 5655 9091 5661
rect 2685 5627 2743 5633
rect 2685 5593 2697 5627
rect 2731 5624 2743 5627
rect 6641 5627 6699 5633
rect 2731 5596 3924 5624
rect 2731 5593 2743 5596
rect 2685 5587 2743 5593
rect 3786 5556 3792 5568
rect 3747 5528 3792 5556
rect 3786 5516 3792 5528
rect 3844 5516 3850 5568
rect 3896 5556 3924 5596
rect 6641 5593 6653 5627
rect 6687 5593 6699 5627
rect 6641 5587 6699 5593
rect 6362 5556 6368 5568
rect 3896 5528 6368 5556
rect 6362 5516 6368 5528
rect 6420 5516 6426 5568
rect 6454 5516 6460 5568
rect 6512 5556 6518 5568
rect 6656 5556 6684 5587
rect 7190 5584 7196 5636
rect 7248 5624 7254 5636
rect 8128 5624 8156 5655
rect 9306 5652 9312 5664
rect 9364 5652 9370 5704
rect 12161 5695 12219 5701
rect 12161 5692 12173 5695
rect 9968 5664 12173 5692
rect 9968 5636 9996 5664
rect 12161 5661 12173 5664
rect 12207 5661 12219 5695
rect 12268 5692 12296 5732
rect 12417 5695 12475 5701
rect 12417 5692 12429 5695
rect 12268 5664 12429 5692
rect 12161 5655 12219 5661
rect 12417 5661 12429 5664
rect 12463 5661 12475 5695
rect 12417 5655 12475 5661
rect 13170 5652 13176 5704
rect 13228 5692 13234 5704
rect 14093 5695 14151 5701
rect 14093 5692 14105 5695
rect 13228 5664 14105 5692
rect 13228 5652 13234 5664
rect 14093 5661 14105 5664
rect 14139 5692 14151 5695
rect 14182 5692 14188 5704
rect 14139 5664 14188 5692
rect 14139 5661 14151 5664
rect 14093 5655 14151 5661
rect 14182 5652 14188 5664
rect 14240 5652 14246 5704
rect 15013 5695 15071 5701
rect 15013 5661 15025 5695
rect 15059 5692 15071 5695
rect 15378 5692 15384 5704
rect 15059 5664 15384 5692
rect 15059 5661 15071 5664
rect 15013 5655 15071 5661
rect 15378 5652 15384 5664
rect 15436 5652 15442 5704
rect 16132 5701 16160 5732
rect 17037 5729 17049 5763
rect 17083 5729 17095 5763
rect 17037 5723 17095 5729
rect 15841 5695 15899 5701
rect 15841 5661 15853 5695
rect 15887 5661 15899 5695
rect 15841 5655 15899 5661
rect 16117 5695 16175 5701
rect 16117 5661 16129 5695
rect 16163 5692 16175 5695
rect 16666 5692 16672 5704
rect 16163 5664 16672 5692
rect 16163 5661 16175 5664
rect 16117 5655 16175 5661
rect 9950 5624 9956 5636
rect 7248 5596 8156 5624
rect 9911 5596 9956 5624
rect 7248 5584 7254 5596
rect 9950 5584 9956 5596
rect 10008 5584 10014 5636
rect 11701 5627 11759 5633
rect 11701 5593 11713 5627
rect 11747 5624 11759 5627
rect 11882 5624 11888 5636
rect 11747 5596 11888 5624
rect 11747 5593 11759 5596
rect 11701 5587 11759 5593
rect 11882 5584 11888 5596
rect 11940 5584 11946 5636
rect 15856 5624 15884 5655
rect 16666 5652 16672 5664
rect 16724 5652 16730 5704
rect 16850 5692 16856 5704
rect 16811 5664 16856 5692
rect 16850 5652 16856 5664
rect 16908 5652 16914 5704
rect 17052 5636 17080 5723
rect 17586 5720 17592 5772
rect 17644 5760 17650 5772
rect 17644 5732 18368 5760
rect 17644 5720 17650 5732
rect 17129 5695 17187 5701
rect 17129 5661 17141 5695
rect 17175 5661 17187 5695
rect 17129 5655 17187 5661
rect 17221 5695 17279 5701
rect 17221 5661 17233 5695
rect 17267 5692 17279 5695
rect 17310 5692 17316 5704
rect 17267 5664 17316 5692
rect 17267 5661 17279 5664
rect 17221 5655 17279 5661
rect 16942 5624 16948 5636
rect 11992 5596 16948 5624
rect 6512 5528 6684 5556
rect 6512 5516 6518 5528
rect 6730 5516 6736 5568
rect 6788 5556 6794 5568
rect 7558 5556 7564 5568
rect 6788 5528 7564 5556
rect 6788 5516 6794 5528
rect 7558 5516 7564 5528
rect 7616 5516 7622 5568
rect 7926 5516 7932 5568
rect 7984 5556 7990 5568
rect 9125 5559 9183 5565
rect 9125 5556 9137 5559
rect 7984 5528 9137 5556
rect 7984 5516 7990 5528
rect 9125 5525 9137 5528
rect 9171 5556 9183 5559
rect 11992 5556 12020 5596
rect 16942 5584 16948 5596
rect 17000 5584 17006 5636
rect 17034 5584 17040 5636
rect 17092 5584 17098 5636
rect 17144 5568 17172 5655
rect 17310 5652 17316 5664
rect 17368 5652 17374 5704
rect 17405 5695 17463 5701
rect 17405 5661 17417 5695
rect 17451 5692 17463 5695
rect 17678 5692 17684 5704
rect 17451 5664 17684 5692
rect 17451 5661 17463 5664
rect 17405 5655 17463 5661
rect 17678 5652 17684 5664
rect 17736 5652 17742 5704
rect 18340 5701 18368 5732
rect 19426 5720 19432 5772
rect 19484 5760 19490 5772
rect 19797 5763 19855 5769
rect 19797 5760 19809 5763
rect 19484 5732 19809 5760
rect 19484 5720 19490 5732
rect 19797 5729 19809 5732
rect 19843 5729 19855 5763
rect 20254 5760 20260 5772
rect 19797 5723 19855 5729
rect 19904 5732 20260 5760
rect 18049 5695 18107 5701
rect 18049 5661 18061 5695
rect 18095 5661 18107 5695
rect 18049 5655 18107 5661
rect 18325 5695 18383 5701
rect 18325 5661 18337 5695
rect 18371 5661 18383 5695
rect 19610 5692 19616 5704
rect 19523 5664 19616 5692
rect 18325 5655 18383 5661
rect 18064 5624 18092 5655
rect 19610 5652 19616 5664
rect 19668 5692 19674 5704
rect 19904 5692 19932 5732
rect 20254 5720 20260 5732
rect 20312 5720 20318 5772
rect 21361 5763 21419 5769
rect 21361 5729 21373 5763
rect 21407 5760 21419 5763
rect 21407 5732 22048 5760
rect 21407 5729 21419 5732
rect 21361 5723 21419 5729
rect 19668 5664 19932 5692
rect 19668 5652 19674 5664
rect 20162 5652 20168 5704
rect 20220 5692 20226 5704
rect 21637 5695 21695 5701
rect 21637 5692 21649 5695
rect 20220 5664 21649 5692
rect 20220 5652 20226 5664
rect 21637 5661 21649 5664
rect 21683 5661 21695 5695
rect 22020 5692 22048 5732
rect 22094 5720 22100 5772
rect 22152 5760 22158 5772
rect 35253 5763 35311 5769
rect 22152 5732 22197 5760
rect 22152 5720 22158 5732
rect 35253 5729 35265 5763
rect 35299 5760 35311 5763
rect 37182 5760 37188 5772
rect 35299 5732 37188 5760
rect 35299 5729 35311 5732
rect 35253 5723 35311 5729
rect 37182 5720 37188 5732
rect 37240 5760 37246 5772
rect 37476 5760 37504 5800
rect 38286 5760 38292 5772
rect 37240 5732 37412 5760
rect 37240 5720 37246 5732
rect 23382 5692 23388 5704
rect 22020 5664 23388 5692
rect 21637 5655 21695 5661
rect 23382 5652 23388 5664
rect 23440 5692 23446 5704
rect 24670 5692 24676 5704
rect 23440 5664 24676 5692
rect 23440 5652 23446 5664
rect 24670 5652 24676 5664
rect 24728 5652 24734 5704
rect 24857 5695 24915 5701
rect 24857 5661 24869 5695
rect 24903 5692 24915 5695
rect 24903 5664 27200 5692
rect 24903 5661 24915 5664
rect 24857 5655 24915 5661
rect 27172 5636 27200 5664
rect 28442 5652 28448 5704
rect 28500 5692 28506 5704
rect 28813 5695 28871 5701
rect 28813 5692 28825 5695
rect 28500 5664 28825 5692
rect 28500 5652 28506 5664
rect 28813 5661 28825 5664
rect 28859 5661 28871 5695
rect 28813 5655 28871 5661
rect 29086 5652 29092 5704
rect 29144 5692 29150 5704
rect 29825 5695 29883 5701
rect 29825 5692 29837 5695
rect 29144 5664 29837 5692
rect 29144 5652 29150 5664
rect 29825 5661 29837 5664
rect 29871 5661 29883 5695
rect 29825 5655 29883 5661
rect 29914 5652 29920 5704
rect 29972 5692 29978 5704
rect 30009 5692 30067 5698
rect 29972 5664 30021 5692
rect 29972 5652 29978 5664
rect 30009 5658 30021 5664
rect 30055 5658 30067 5692
rect 30009 5652 30067 5658
rect 30098 5652 30104 5704
rect 30156 5692 30162 5704
rect 30282 5701 30288 5704
rect 30239 5695 30288 5701
rect 30156 5664 30201 5692
rect 30156 5652 30162 5664
rect 30239 5661 30251 5695
rect 30285 5661 30288 5695
rect 30239 5655 30288 5661
rect 30282 5652 30288 5655
rect 30340 5652 30346 5704
rect 31941 5695 31999 5701
rect 31941 5692 31953 5695
rect 30484 5664 31953 5692
rect 17328 5596 18092 5624
rect 18233 5627 18291 5633
rect 17328 5568 17356 5596
rect 18233 5593 18245 5627
rect 18279 5624 18291 5627
rect 22364 5627 22422 5633
rect 18279 5596 19748 5624
rect 18279 5593 18291 5596
rect 18233 5587 18291 5593
rect 9171 5528 12020 5556
rect 9171 5525 9183 5528
rect 9125 5519 9183 5525
rect 12342 5516 12348 5568
rect 12400 5556 12406 5568
rect 12618 5556 12624 5568
rect 12400 5528 12624 5556
rect 12400 5516 12406 5528
rect 12618 5516 12624 5528
rect 12676 5516 12682 5568
rect 13538 5556 13544 5568
rect 13499 5528 13544 5556
rect 13538 5516 13544 5528
rect 13596 5516 13602 5568
rect 14277 5559 14335 5565
rect 14277 5525 14289 5559
rect 14323 5556 14335 5559
rect 14366 5556 14372 5568
rect 14323 5528 14372 5556
rect 14323 5525 14335 5528
rect 14277 5519 14335 5525
rect 14366 5516 14372 5528
rect 14424 5516 14430 5568
rect 15930 5516 15936 5568
rect 15988 5556 15994 5568
rect 16025 5559 16083 5565
rect 16025 5556 16037 5559
rect 15988 5528 16037 5556
rect 15988 5516 15994 5528
rect 16025 5525 16037 5528
rect 16071 5525 16083 5559
rect 16025 5519 16083 5525
rect 17126 5516 17132 5568
rect 17184 5516 17190 5568
rect 17310 5516 17316 5568
rect 17368 5516 17374 5568
rect 19150 5516 19156 5568
rect 19208 5556 19214 5568
rect 19720 5565 19748 5596
rect 22364 5593 22376 5627
rect 22410 5624 22422 5627
rect 23290 5624 23296 5636
rect 22410 5596 23296 5624
rect 22410 5593 22422 5596
rect 22364 5587 22422 5593
rect 23290 5584 23296 5596
rect 23348 5584 23354 5636
rect 25038 5624 25044 5636
rect 24504 5596 25044 5624
rect 19245 5559 19303 5565
rect 19245 5556 19257 5559
rect 19208 5528 19257 5556
rect 19208 5516 19214 5528
rect 19245 5525 19257 5528
rect 19291 5525 19303 5559
rect 19245 5519 19303 5525
rect 19705 5559 19763 5565
rect 19705 5525 19717 5559
rect 19751 5556 19763 5559
rect 20254 5556 20260 5568
rect 19751 5528 20260 5556
rect 19751 5525 19763 5528
rect 19705 5519 19763 5525
rect 20254 5516 20260 5528
rect 20312 5516 20318 5568
rect 23014 5516 23020 5568
rect 23072 5556 23078 5568
rect 24504 5556 24532 5596
rect 25038 5584 25044 5596
rect 25096 5584 25102 5636
rect 25590 5624 25596 5636
rect 25551 5596 25596 5624
rect 25590 5584 25596 5596
rect 25648 5584 25654 5636
rect 26418 5624 26424 5636
rect 26379 5596 26424 5624
rect 26418 5584 26424 5596
rect 26476 5584 26482 5636
rect 27154 5584 27160 5636
rect 27212 5584 27218 5636
rect 28629 5627 28687 5633
rect 28629 5593 28641 5627
rect 28675 5624 28687 5627
rect 29178 5624 29184 5636
rect 28675 5596 29184 5624
rect 28675 5593 28687 5596
rect 28629 5587 28687 5593
rect 29178 5584 29184 5596
rect 29236 5584 29242 5636
rect 23072 5528 24532 5556
rect 24673 5559 24731 5565
rect 23072 5516 23078 5528
rect 24673 5525 24685 5559
rect 24719 5556 24731 5559
rect 24762 5556 24768 5568
rect 24719 5528 24768 5556
rect 24719 5525 24731 5528
rect 24673 5519 24731 5525
rect 24762 5516 24768 5528
rect 24820 5516 24826 5568
rect 27065 5559 27123 5565
rect 27065 5525 27077 5559
rect 27111 5556 27123 5559
rect 27614 5556 27620 5568
rect 27111 5528 27620 5556
rect 27111 5525 27123 5528
rect 27065 5519 27123 5525
rect 27614 5516 27620 5528
rect 27672 5556 27678 5568
rect 30484 5556 30512 5664
rect 31941 5661 31953 5664
rect 31987 5692 31999 5695
rect 34149 5695 34207 5701
rect 34149 5692 34161 5695
rect 31987 5664 34161 5692
rect 31987 5661 31999 5664
rect 31941 5655 31999 5661
rect 34149 5661 34161 5664
rect 34195 5661 34207 5695
rect 35526 5692 35532 5704
rect 35487 5664 35532 5692
rect 34149 5655 34207 5661
rect 35526 5652 35532 5664
rect 35584 5652 35590 5704
rect 36446 5652 36452 5704
rect 36504 5692 36510 5704
rect 37093 5695 37151 5701
rect 37093 5692 37105 5695
rect 36504 5664 37105 5692
rect 36504 5652 36510 5664
rect 37093 5661 37105 5664
rect 37139 5661 37151 5695
rect 37274 5692 37280 5704
rect 37235 5664 37280 5692
rect 37093 5655 37151 5661
rect 31570 5584 31576 5636
rect 31628 5624 31634 5636
rect 32401 5627 32459 5633
rect 32401 5624 32413 5627
rect 31628 5596 32413 5624
rect 31628 5584 31634 5596
rect 32401 5593 32413 5596
rect 32447 5593 32459 5627
rect 37108 5624 37136 5655
rect 37274 5652 37280 5664
rect 37332 5652 37338 5704
rect 37384 5701 37412 5732
rect 37476 5732 38292 5760
rect 37476 5701 37504 5732
rect 38286 5720 38292 5732
rect 38344 5720 38350 5772
rect 37369 5695 37427 5701
rect 37369 5661 37381 5695
rect 37415 5661 37427 5695
rect 37369 5655 37427 5661
rect 37461 5695 37519 5701
rect 37461 5661 37473 5695
rect 37507 5661 37519 5695
rect 37461 5655 37519 5661
rect 38102 5624 38108 5636
rect 37108 5596 38108 5624
rect 32401 5587 32459 5593
rect 38102 5584 38108 5596
rect 38160 5584 38166 5636
rect 27672 5528 30512 5556
rect 27672 5516 27678 5528
rect 34698 5516 34704 5568
rect 34756 5556 34762 5568
rect 37366 5556 37372 5568
rect 34756 5528 37372 5556
rect 34756 5516 34762 5528
rect 37366 5516 37372 5528
rect 37424 5516 37430 5568
rect 37734 5556 37740 5568
rect 37695 5528 37740 5556
rect 37734 5516 37740 5528
rect 37792 5516 37798 5568
rect 1104 5466 68816 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 68816 5466
rect 1104 5392 68816 5414
rect 3789 5355 3847 5361
rect 3789 5321 3801 5355
rect 3835 5352 3847 5355
rect 8110 5352 8116 5364
rect 3835 5324 7972 5352
rect 8071 5324 8116 5352
rect 3835 5321 3847 5324
rect 3789 5315 3847 5321
rect 3237 5287 3295 5293
rect 3237 5253 3249 5287
rect 3283 5284 3295 5287
rect 6822 5284 6828 5296
rect 3283 5256 6828 5284
rect 3283 5253 3295 5256
rect 3237 5247 3295 5253
rect 6822 5244 6828 5256
rect 6880 5244 6886 5296
rect 7745 5287 7803 5293
rect 7745 5284 7757 5287
rect 6932 5256 7757 5284
rect 2222 5216 2228 5228
rect 2183 5188 2228 5216
rect 2222 5176 2228 5188
rect 2280 5176 2286 5228
rect 4985 5219 5043 5225
rect 4985 5185 4997 5219
rect 5031 5216 5043 5219
rect 5445 5219 5503 5225
rect 5445 5216 5457 5219
rect 5031 5188 5457 5216
rect 5031 5185 5043 5188
rect 4985 5179 5043 5185
rect 5445 5185 5457 5188
rect 5491 5185 5503 5219
rect 5445 5179 5503 5185
rect 5629 5219 5687 5225
rect 5629 5185 5641 5219
rect 5675 5185 5687 5219
rect 5629 5179 5687 5185
rect 5534 5148 5540 5160
rect 2746 5120 5540 5148
rect 1765 5083 1823 5089
rect 1765 5049 1777 5083
rect 1811 5080 1823 5083
rect 2746 5080 2774 5120
rect 5534 5108 5540 5120
rect 5592 5108 5598 5160
rect 1811 5052 2774 5080
rect 4341 5083 4399 5089
rect 1811 5049 1823 5052
rect 1765 5043 1823 5049
rect 4341 5049 4353 5083
rect 4387 5080 4399 5083
rect 5644 5080 5672 5179
rect 6932 5160 6960 5256
rect 7745 5253 7757 5256
rect 7791 5253 7803 5287
rect 7944 5284 7972 5324
rect 8110 5312 8116 5324
rect 8168 5312 8174 5364
rect 9490 5352 9496 5364
rect 9451 5324 9496 5352
rect 9490 5312 9496 5324
rect 9548 5312 9554 5364
rect 11238 5312 11244 5364
rect 11296 5352 11302 5364
rect 13078 5352 13084 5364
rect 11296 5324 13084 5352
rect 11296 5312 11302 5324
rect 13078 5312 13084 5324
rect 13136 5352 13142 5364
rect 14461 5355 14519 5361
rect 13136 5324 13768 5352
rect 13136 5312 13142 5324
rect 8846 5284 8852 5296
rect 7944 5256 8852 5284
rect 7745 5247 7803 5253
rect 8846 5244 8852 5256
rect 8904 5244 8910 5296
rect 11054 5284 11060 5296
rect 10796 5256 11060 5284
rect 7650 5216 7656 5228
rect 7611 5188 7656 5216
rect 7650 5176 7656 5188
rect 7708 5176 7714 5228
rect 7926 5216 7932 5228
rect 7887 5188 7932 5216
rect 7926 5176 7932 5188
rect 7984 5176 7990 5228
rect 9490 5216 9496 5228
rect 9451 5188 9496 5216
rect 9490 5176 9496 5188
rect 9548 5176 9554 5228
rect 9766 5216 9772 5228
rect 9727 5188 9772 5216
rect 9766 5176 9772 5188
rect 9824 5176 9830 5228
rect 10042 5216 10048 5228
rect 10003 5188 10048 5216
rect 10042 5176 10048 5188
rect 10100 5176 10106 5228
rect 5813 5151 5871 5157
rect 5813 5117 5825 5151
rect 5859 5148 5871 5151
rect 6914 5148 6920 5160
rect 5859 5120 6776 5148
rect 6875 5120 6920 5148
rect 5859 5117 5871 5120
rect 5813 5111 5871 5117
rect 6457 5083 6515 5089
rect 6457 5080 6469 5083
rect 4387 5052 5580 5080
rect 5644 5052 6469 5080
rect 4387 5049 4399 5052
rect 4341 5043 4399 5049
rect 2409 5015 2467 5021
rect 2409 4981 2421 5015
rect 2455 5012 2467 5015
rect 2958 5012 2964 5024
rect 2455 4984 2964 5012
rect 2455 4981 2467 4984
rect 2409 4975 2467 4981
rect 2958 4972 2964 4984
rect 3016 4972 3022 5024
rect 4706 4972 4712 5024
rect 4764 5012 4770 5024
rect 4801 5015 4859 5021
rect 4801 5012 4813 5015
rect 4764 4984 4813 5012
rect 4764 4972 4770 4984
rect 4801 4981 4813 4984
rect 4847 4981 4859 5015
rect 5552 5012 5580 5052
rect 6457 5049 6469 5052
rect 6503 5049 6515 5083
rect 6748 5080 6776 5120
rect 6914 5108 6920 5120
rect 6972 5108 6978 5160
rect 7101 5151 7159 5157
rect 7101 5117 7113 5151
rect 7147 5148 7159 5151
rect 7466 5148 7472 5160
rect 7147 5120 7472 5148
rect 7147 5117 7159 5120
rect 7101 5111 7159 5117
rect 7466 5108 7472 5120
rect 7524 5108 7530 5160
rect 10796 5148 10824 5256
rect 11054 5244 11060 5256
rect 11112 5244 11118 5296
rect 13262 5284 13268 5296
rect 12176 5256 13268 5284
rect 10962 5216 10968 5228
rect 10923 5188 10968 5216
rect 10962 5176 10968 5188
rect 11020 5176 11026 5228
rect 12176 5225 12204 5256
rect 13262 5244 13268 5256
rect 13320 5244 13326 5296
rect 13740 5293 13768 5324
rect 14461 5321 14473 5355
rect 14507 5352 14519 5355
rect 14642 5352 14648 5364
rect 14507 5324 14648 5352
rect 14507 5321 14519 5324
rect 14461 5315 14519 5321
rect 14642 5312 14648 5324
rect 14700 5312 14706 5364
rect 17126 5352 17132 5364
rect 17087 5324 17132 5352
rect 17126 5312 17132 5324
rect 17184 5312 17190 5364
rect 17497 5355 17555 5361
rect 17497 5321 17509 5355
rect 17543 5352 17555 5355
rect 18230 5352 18236 5364
rect 17543 5324 18236 5352
rect 17543 5321 17555 5324
rect 17497 5315 17555 5321
rect 18230 5312 18236 5324
rect 18288 5312 18294 5364
rect 23290 5352 23296 5364
rect 23251 5324 23296 5352
rect 23290 5312 23296 5324
rect 23348 5312 23354 5364
rect 28442 5312 28448 5364
rect 28500 5352 28506 5364
rect 29825 5355 29883 5361
rect 29825 5352 29837 5355
rect 28500 5324 29837 5352
rect 28500 5312 28506 5324
rect 29825 5321 29837 5324
rect 29871 5321 29883 5355
rect 29825 5315 29883 5321
rect 32401 5355 32459 5361
rect 32401 5321 32413 5355
rect 32447 5352 32459 5355
rect 32858 5352 32864 5364
rect 32447 5324 32864 5352
rect 32447 5321 32459 5324
rect 32401 5315 32459 5321
rect 32858 5312 32864 5324
rect 32916 5312 32922 5364
rect 34606 5312 34612 5364
rect 34664 5352 34670 5364
rect 35069 5355 35127 5361
rect 35069 5352 35081 5355
rect 34664 5324 35081 5352
rect 34664 5312 34670 5324
rect 35069 5321 35081 5324
rect 35115 5321 35127 5355
rect 35069 5315 35127 5321
rect 37274 5312 37280 5364
rect 37332 5352 37338 5364
rect 37645 5355 37703 5361
rect 37645 5352 37657 5355
rect 37332 5324 37657 5352
rect 37332 5312 37338 5324
rect 37645 5321 37657 5324
rect 37691 5321 37703 5355
rect 37645 5315 37703 5321
rect 38654 5312 38660 5364
rect 38712 5352 38718 5364
rect 40313 5355 40371 5361
rect 40313 5352 40325 5355
rect 38712 5324 40325 5352
rect 38712 5312 38718 5324
rect 40313 5321 40325 5324
rect 40359 5321 40371 5355
rect 40313 5315 40371 5321
rect 13725 5287 13783 5293
rect 13725 5253 13737 5287
rect 13771 5253 13783 5287
rect 13725 5247 13783 5253
rect 13906 5244 13912 5296
rect 13964 5244 13970 5296
rect 16666 5244 16672 5296
rect 16724 5284 16730 5296
rect 21266 5284 21272 5296
rect 16724 5256 17448 5284
rect 16724 5244 16730 5256
rect 12161 5219 12219 5225
rect 12161 5216 12173 5219
rect 11808 5188 12173 5216
rect 7760 5120 10824 5148
rect 7190 5080 7196 5092
rect 6748 5052 7196 5080
rect 6457 5043 6515 5049
rect 7190 5040 7196 5052
rect 7248 5040 7254 5092
rect 7760 5012 7788 5120
rect 10870 5108 10876 5160
rect 10928 5148 10934 5160
rect 11808 5148 11836 5188
rect 12161 5185 12173 5188
rect 12207 5185 12219 5219
rect 12161 5179 12219 5185
rect 12342 5176 12348 5228
rect 12400 5216 12406 5228
rect 12621 5219 12679 5225
rect 12621 5216 12633 5219
rect 12400 5188 12633 5216
rect 12400 5176 12406 5188
rect 12621 5185 12633 5188
rect 12667 5185 12679 5219
rect 12621 5179 12679 5185
rect 12897 5219 12955 5225
rect 12897 5185 12909 5219
rect 12943 5216 12955 5219
rect 13924 5216 13952 5244
rect 14090 5216 14096 5228
rect 12943 5188 14096 5216
rect 12943 5185 12955 5188
rect 12897 5179 12955 5185
rect 14090 5176 14096 5188
rect 14148 5216 14154 5228
rect 14185 5219 14243 5225
rect 14185 5216 14197 5219
rect 14148 5188 14197 5216
rect 14148 5176 14154 5188
rect 14185 5185 14197 5188
rect 14231 5185 14243 5219
rect 15194 5216 15200 5228
rect 15155 5188 15200 5216
rect 14185 5179 14243 5185
rect 15194 5176 15200 5188
rect 15252 5176 15258 5228
rect 16942 5176 16948 5228
rect 17000 5216 17006 5228
rect 17310 5216 17316 5228
rect 17000 5188 17316 5216
rect 17000 5176 17006 5188
rect 17310 5176 17316 5188
rect 17368 5176 17374 5228
rect 17420 5216 17448 5256
rect 17696 5256 21272 5284
rect 17586 5225 17592 5228
rect 17573 5219 17592 5225
rect 17573 5216 17585 5219
rect 17420 5188 17585 5216
rect 17573 5185 17585 5188
rect 17573 5179 17592 5185
rect 17586 5176 17592 5179
rect 17644 5176 17650 5228
rect 10928 5120 11836 5148
rect 11885 5151 11943 5157
rect 10928 5108 10934 5120
rect 11885 5117 11897 5151
rect 11931 5148 11943 5151
rect 11974 5148 11980 5160
rect 11931 5120 11980 5148
rect 11931 5117 11943 5120
rect 11885 5111 11943 5117
rect 11974 5108 11980 5120
rect 12032 5108 12038 5160
rect 12805 5151 12863 5157
rect 12805 5117 12817 5151
rect 12851 5148 12863 5151
rect 13906 5148 13912 5160
rect 12851 5120 13912 5148
rect 12851 5117 12863 5120
rect 12805 5111 12863 5117
rect 13906 5108 13912 5120
rect 13964 5108 13970 5160
rect 14277 5151 14335 5157
rect 14277 5117 14289 5151
rect 14323 5117 14335 5151
rect 14277 5111 14335 5117
rect 8938 5040 8944 5092
rect 8996 5080 9002 5092
rect 9033 5083 9091 5089
rect 9033 5080 9045 5083
rect 8996 5052 9045 5080
rect 8996 5040 9002 5052
rect 9033 5049 9045 5052
rect 9079 5049 9091 5083
rect 11609 5083 11667 5089
rect 11609 5080 11621 5083
rect 9033 5043 9091 5049
rect 9140 5052 11621 5080
rect 5552 4984 7788 5012
rect 4801 4975 4859 4981
rect 7834 4972 7840 5024
rect 7892 5012 7898 5024
rect 9140 5012 9168 5052
rect 11609 5049 11621 5052
rect 11655 5049 11667 5083
rect 12894 5080 12900 5092
rect 11609 5043 11667 5049
rect 12084 5052 12900 5080
rect 7892 4984 9168 5012
rect 10781 5015 10839 5021
rect 7892 4972 7898 4984
rect 10781 4981 10793 5015
rect 10827 5012 10839 5015
rect 10962 5012 10968 5024
rect 10827 4984 10968 5012
rect 10827 4981 10839 4984
rect 10781 4975 10839 4981
rect 10962 4972 10968 4984
rect 11020 4972 11026 5024
rect 12084 5021 12112 5052
rect 12894 5040 12900 5052
rect 12952 5080 12958 5092
rect 12952 5052 13124 5080
rect 12952 5040 12958 5052
rect 12069 5015 12127 5021
rect 12069 4981 12081 5015
rect 12115 4981 12127 5015
rect 12069 4975 12127 4981
rect 12526 4972 12532 5024
rect 12584 5012 12590 5024
rect 13096 5021 13124 5052
rect 13630 5040 13636 5092
rect 13688 5080 13694 5092
rect 13725 5083 13783 5089
rect 13725 5080 13737 5083
rect 13688 5052 13737 5080
rect 13688 5040 13694 5052
rect 13725 5049 13737 5052
rect 13771 5049 13783 5083
rect 13725 5043 13783 5049
rect 13814 5040 13820 5092
rect 13872 5080 13878 5092
rect 14292 5080 14320 5111
rect 14366 5108 14372 5160
rect 14424 5148 14430 5160
rect 14424 5120 14872 5148
rect 14424 5108 14430 5120
rect 14734 5080 14740 5092
rect 13872 5052 14740 5080
rect 13872 5040 13878 5052
rect 14734 5040 14740 5052
rect 14792 5040 14798 5092
rect 14844 5080 14872 5120
rect 17696 5080 17724 5256
rect 21266 5244 21272 5256
rect 21324 5244 21330 5296
rect 24670 5244 24676 5296
rect 24728 5284 24734 5296
rect 24728 5256 24900 5284
rect 24728 5244 24734 5256
rect 18325 5219 18383 5225
rect 18325 5185 18337 5219
rect 18371 5216 18383 5219
rect 18782 5216 18788 5228
rect 18371 5188 18788 5216
rect 18371 5185 18383 5188
rect 18325 5179 18383 5185
rect 18782 5176 18788 5188
rect 18840 5176 18846 5228
rect 19150 5216 19156 5228
rect 19111 5188 19156 5216
rect 19150 5176 19156 5188
rect 19208 5176 19214 5228
rect 19337 5219 19395 5225
rect 19337 5185 19349 5219
rect 19383 5216 19395 5219
rect 19797 5219 19855 5225
rect 19797 5216 19809 5219
rect 19383 5188 19809 5216
rect 19383 5185 19395 5188
rect 19337 5179 19395 5185
rect 19797 5185 19809 5188
rect 19843 5185 19855 5219
rect 22002 5216 22008 5228
rect 21963 5188 22008 5216
rect 19797 5179 19855 5185
rect 22002 5176 22008 5188
rect 22060 5176 22066 5228
rect 22738 5176 22744 5228
rect 22796 5216 22802 5228
rect 23569 5219 23627 5225
rect 23569 5216 23581 5219
rect 22796 5188 23581 5216
rect 22796 5176 22802 5188
rect 23569 5185 23581 5188
rect 23615 5185 23627 5219
rect 23569 5179 23627 5185
rect 23658 5222 23716 5228
rect 23658 5188 23670 5222
rect 23704 5188 23716 5222
rect 23658 5182 23716 5188
rect 18506 5108 18512 5160
rect 18564 5148 18570 5160
rect 18969 5151 19027 5157
rect 18969 5148 18981 5151
rect 18564 5120 18981 5148
rect 18564 5108 18570 5120
rect 18969 5117 18981 5120
rect 19015 5117 19027 5151
rect 18969 5111 19027 5117
rect 19978 5108 19984 5160
rect 20036 5148 20042 5160
rect 20438 5148 20444 5160
rect 20036 5120 20444 5148
rect 20036 5108 20042 5120
rect 20438 5108 20444 5120
rect 20496 5108 20502 5160
rect 20717 5151 20775 5157
rect 20717 5117 20729 5151
rect 20763 5117 20775 5151
rect 20717 5111 20775 5117
rect 14844 5052 17724 5080
rect 18138 5040 18144 5092
rect 18196 5080 18202 5092
rect 19426 5080 19432 5092
rect 18196 5052 19432 5080
rect 18196 5040 18202 5052
rect 19426 5040 19432 5052
rect 19484 5040 19490 5092
rect 20732 5080 20760 5111
rect 23382 5108 23388 5160
rect 23440 5148 23446 5160
rect 23673 5148 23701 5182
rect 23750 5174 23756 5226
rect 23808 5225 23814 5226
rect 23808 5216 23816 5225
rect 23937 5219 23995 5225
rect 23808 5188 23851 5216
rect 23808 5179 23816 5188
rect 23937 5185 23949 5219
rect 23983 5216 23995 5219
rect 24578 5216 24584 5228
rect 23983 5188 24584 5216
rect 23983 5185 23995 5188
rect 23937 5179 23995 5185
rect 23808 5174 23814 5179
rect 23440 5120 23701 5148
rect 23440 5108 23446 5120
rect 23198 5080 23204 5092
rect 20732 5052 23204 5080
rect 23198 5040 23204 5052
rect 23256 5080 23262 5092
rect 23952 5080 23980 5179
rect 24578 5176 24584 5188
rect 24636 5176 24642 5228
rect 24762 5216 24768 5228
rect 24723 5188 24768 5216
rect 24762 5176 24768 5188
rect 24820 5176 24826 5228
rect 24872 5225 24900 5256
rect 25038 5244 25044 5296
rect 25096 5284 25102 5296
rect 26053 5287 26111 5293
rect 26053 5284 26065 5287
rect 25096 5256 26065 5284
rect 25096 5244 25102 5256
rect 26053 5253 26065 5256
rect 26099 5284 26111 5287
rect 27341 5287 27399 5293
rect 27341 5284 27353 5287
rect 26099 5256 27353 5284
rect 26099 5253 26111 5256
rect 26053 5247 26111 5253
rect 27341 5253 27353 5256
rect 27387 5253 27399 5287
rect 27341 5247 27399 5253
rect 28994 5244 29000 5296
rect 29052 5284 29058 5296
rect 30834 5284 30840 5296
rect 29052 5256 30840 5284
rect 29052 5244 29058 5256
rect 30834 5244 30840 5256
rect 30892 5284 30898 5296
rect 31570 5284 31576 5296
rect 30892 5256 31576 5284
rect 30892 5244 30898 5256
rect 24857 5219 24915 5225
rect 24857 5185 24869 5219
rect 24903 5185 24915 5219
rect 24857 5179 24915 5185
rect 24872 5148 24900 5179
rect 24946 5176 24952 5228
rect 25004 5216 25010 5228
rect 26237 5219 26295 5225
rect 25004 5188 25049 5216
rect 25004 5176 25010 5188
rect 26237 5185 26249 5219
rect 26283 5216 26295 5219
rect 27246 5216 27252 5228
rect 26283 5188 27252 5216
rect 26283 5185 26295 5188
rect 26237 5179 26295 5185
rect 27246 5176 27252 5188
rect 27304 5176 27310 5228
rect 27525 5219 27583 5225
rect 27525 5185 27537 5219
rect 27571 5216 27583 5219
rect 27798 5216 27804 5228
rect 27571 5188 27804 5216
rect 27571 5185 27583 5188
rect 27525 5179 27583 5185
rect 27798 5176 27804 5188
rect 27856 5176 27862 5228
rect 30558 5176 30564 5228
rect 30616 5216 30622 5228
rect 31220 5225 31248 5256
rect 31570 5244 31576 5256
rect 31628 5244 31634 5296
rect 30938 5219 30996 5225
rect 30938 5216 30950 5219
rect 30616 5188 30950 5216
rect 30616 5176 30622 5188
rect 30938 5185 30950 5188
rect 30984 5185 30996 5219
rect 30938 5179 30996 5185
rect 31205 5219 31263 5225
rect 31205 5185 31217 5219
rect 31251 5185 31263 5219
rect 32876 5216 32904 5312
rect 37182 5284 37188 5296
rect 33244 5256 37188 5284
rect 33244 5225 33272 5256
rect 33137 5219 33195 5225
rect 33137 5216 33149 5219
rect 32876 5188 33149 5216
rect 31205 5179 31263 5185
rect 33137 5185 33149 5188
rect 33183 5185 33195 5219
rect 33137 5179 33195 5185
rect 33229 5219 33287 5225
rect 33229 5185 33241 5219
rect 33275 5185 33287 5219
rect 33229 5179 33287 5185
rect 33318 5176 33324 5228
rect 33376 5216 33382 5228
rect 33505 5219 33563 5225
rect 33376 5188 33421 5216
rect 33376 5176 33382 5188
rect 33505 5185 33517 5219
rect 33551 5185 33563 5219
rect 33505 5179 33563 5185
rect 26786 5148 26792 5160
rect 24872 5120 26792 5148
rect 26786 5108 26792 5120
rect 26844 5108 26850 5160
rect 33520 5148 33548 5179
rect 33870 5176 33876 5228
rect 33928 5216 33934 5228
rect 34348 5225 34376 5256
rect 34241 5219 34299 5225
rect 34241 5216 34253 5219
rect 33928 5188 34253 5216
rect 33928 5176 33934 5188
rect 34241 5185 34253 5188
rect 34287 5185 34299 5219
rect 34241 5179 34299 5185
rect 34333 5219 34391 5225
rect 34333 5185 34345 5219
rect 34379 5185 34391 5219
rect 34333 5179 34391 5185
rect 34422 5176 34428 5228
rect 34480 5216 34486 5228
rect 34609 5219 34667 5225
rect 34480 5188 34525 5216
rect 34480 5176 34486 5188
rect 34609 5185 34621 5219
rect 34655 5216 34667 5219
rect 35342 5216 35348 5228
rect 34655 5188 35348 5216
rect 34655 5185 34667 5188
rect 34609 5179 34667 5185
rect 34624 5148 34652 5179
rect 35342 5176 35348 5188
rect 35400 5176 35406 5228
rect 35986 5176 35992 5228
rect 36044 5216 36050 5228
rect 36188 5225 36216 5256
rect 37182 5244 37188 5256
rect 37240 5244 37246 5296
rect 37458 5284 37464 5296
rect 37419 5256 37464 5284
rect 37458 5244 37464 5256
rect 37516 5244 37522 5296
rect 38746 5244 38752 5296
rect 38804 5284 38810 5296
rect 39178 5287 39236 5293
rect 39178 5284 39190 5287
rect 38804 5256 39190 5284
rect 38804 5244 38810 5256
rect 39178 5253 39190 5256
rect 39224 5253 39236 5287
rect 39178 5247 39236 5253
rect 36081 5219 36139 5225
rect 36081 5216 36093 5219
rect 36044 5188 36093 5216
rect 36044 5176 36050 5188
rect 36081 5185 36093 5188
rect 36127 5185 36139 5219
rect 36081 5179 36139 5185
rect 36173 5219 36231 5225
rect 36173 5185 36185 5219
rect 36219 5185 36231 5219
rect 36173 5179 36231 5185
rect 36262 5176 36268 5228
rect 36320 5216 36326 5228
rect 36320 5188 36365 5216
rect 36320 5176 36326 5188
rect 36446 5176 36452 5228
rect 36504 5216 36510 5228
rect 37277 5219 37335 5225
rect 36504 5188 36549 5216
rect 36504 5176 36510 5188
rect 37277 5185 37289 5219
rect 37323 5216 37335 5219
rect 37366 5216 37372 5228
rect 37323 5188 37372 5216
rect 37323 5185 37335 5188
rect 37277 5179 37335 5185
rect 37366 5176 37372 5188
rect 37424 5176 37430 5228
rect 33520 5120 34652 5148
rect 38746 5108 38752 5160
rect 38804 5148 38810 5160
rect 38933 5151 38991 5157
rect 38933 5148 38945 5151
rect 38804 5120 38945 5148
rect 38804 5108 38810 5120
rect 38933 5117 38945 5120
rect 38979 5117 38991 5151
rect 38933 5111 38991 5117
rect 58802 5108 58808 5160
rect 58860 5148 58866 5160
rect 59449 5151 59507 5157
rect 59449 5148 59461 5151
rect 58860 5120 59461 5148
rect 58860 5108 58866 5120
rect 59449 5117 59461 5120
rect 59495 5117 59507 5151
rect 59449 5111 59507 5117
rect 23256 5052 23704 5080
rect 23256 5040 23262 5052
rect 12621 5015 12679 5021
rect 12621 5012 12633 5015
rect 12584 4984 12633 5012
rect 12584 4972 12590 4984
rect 12621 4981 12633 4984
rect 12667 4981 12679 5015
rect 12621 4975 12679 4981
rect 13081 5015 13139 5021
rect 13081 4981 13093 5015
rect 13127 4981 13139 5015
rect 13081 4975 13139 4981
rect 13998 4972 14004 5024
rect 14056 5012 14062 5024
rect 15013 5015 15071 5021
rect 15013 5012 15025 5015
rect 14056 4984 15025 5012
rect 14056 4972 14062 4984
rect 15013 4981 15025 4984
rect 15059 4981 15071 5015
rect 15013 4975 15071 4981
rect 16117 5015 16175 5021
rect 16117 4981 16129 5015
rect 16163 5012 16175 5015
rect 17862 5012 17868 5024
rect 16163 4984 17868 5012
rect 16163 4981 16175 4984
rect 16117 4975 16175 4981
rect 17862 4972 17868 4984
rect 17920 4972 17926 5024
rect 18509 5015 18567 5021
rect 18509 4981 18521 5015
rect 18555 5012 18567 5015
rect 19334 5012 19340 5024
rect 18555 4984 19340 5012
rect 18555 4981 18567 4984
rect 18509 4975 18567 4981
rect 19334 4972 19340 4984
rect 19392 4972 19398 5024
rect 19978 5012 19984 5024
rect 19939 4984 19984 5012
rect 19978 4972 19984 4984
rect 20036 4972 20042 5024
rect 20070 4972 20076 5024
rect 20128 5012 20134 5024
rect 21821 5015 21879 5021
rect 21821 5012 21833 5015
rect 20128 4984 21833 5012
rect 20128 4972 20134 4984
rect 21821 4981 21833 4984
rect 21867 4981 21879 5015
rect 22738 5012 22744 5024
rect 22699 4984 22744 5012
rect 21821 4975 21879 4981
rect 22738 4972 22744 4984
rect 22796 4972 22802 5024
rect 23676 5012 23704 5052
rect 23860 5052 23980 5080
rect 23860 5012 23888 5052
rect 59262 5040 59268 5092
rect 59320 5080 59326 5092
rect 60093 5083 60151 5089
rect 60093 5080 60105 5083
rect 59320 5052 60105 5080
rect 59320 5040 59326 5052
rect 60093 5049 60105 5052
rect 60139 5049 60151 5083
rect 60093 5043 60151 5049
rect 25222 5012 25228 5024
rect 23676 4984 23888 5012
rect 25183 4984 25228 5012
rect 25222 4972 25228 4984
rect 25280 4972 25286 5024
rect 26421 5015 26479 5021
rect 26421 4981 26433 5015
rect 26467 5012 26479 5015
rect 26694 5012 26700 5024
rect 26467 4984 26700 5012
rect 26467 4981 26479 4984
rect 26421 4975 26479 4981
rect 26694 4972 26700 4984
rect 26752 4972 26758 5024
rect 27614 4972 27620 5024
rect 27672 5012 27678 5024
rect 27709 5015 27767 5021
rect 27709 5012 27721 5015
rect 27672 4984 27721 5012
rect 27672 4972 27678 4984
rect 27709 4981 27721 4984
rect 27755 4981 27767 5015
rect 32858 5012 32864 5024
rect 32819 4984 32864 5012
rect 27709 4975 27767 4981
rect 32858 4972 32864 4984
rect 32916 4972 32922 5024
rect 33778 4972 33784 5024
rect 33836 5012 33842 5024
rect 33965 5015 34023 5021
rect 33965 5012 33977 5015
rect 33836 4984 33977 5012
rect 33836 4972 33842 4984
rect 33965 4981 33977 4984
rect 34011 4981 34023 5015
rect 33965 4975 34023 4981
rect 35618 4972 35624 5024
rect 35676 5012 35682 5024
rect 35805 5015 35863 5021
rect 35805 5012 35817 5015
rect 35676 4984 35817 5012
rect 35676 4972 35682 4984
rect 35805 4981 35817 4984
rect 35851 4981 35863 5015
rect 35805 4975 35863 4981
rect 58710 4972 58716 5024
rect 58768 5012 58774 5024
rect 58805 5015 58863 5021
rect 58805 5012 58817 5015
rect 58768 4984 58817 5012
rect 58768 4972 58774 4984
rect 58805 4981 58817 4984
rect 58851 4981 58863 5015
rect 67634 5012 67640 5024
rect 67595 4984 67640 5012
rect 58805 4975 58863 4981
rect 67634 4972 67640 4984
rect 67692 4972 67698 5024
rect 1104 4922 68816 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 65654 4922
rect 65706 4870 65718 4922
rect 65770 4870 65782 4922
rect 65834 4870 65846 4922
rect 65898 4870 65910 4922
rect 65962 4870 68816 4922
rect 1104 4848 68816 4870
rect 5813 4811 5871 4817
rect 5813 4777 5825 4811
rect 5859 4808 5871 4811
rect 6914 4808 6920 4820
rect 5859 4780 6920 4808
rect 5859 4777 5871 4780
rect 5813 4771 5871 4777
rect 6914 4768 6920 4780
rect 6972 4768 6978 4820
rect 9401 4811 9459 4817
rect 9401 4777 9413 4811
rect 9447 4808 9459 4811
rect 9766 4808 9772 4820
rect 9447 4780 9772 4808
rect 9447 4777 9459 4780
rect 9401 4771 9459 4777
rect 9766 4768 9772 4780
rect 9824 4808 9830 4820
rect 10594 4808 10600 4820
rect 9824 4780 10600 4808
rect 9824 4768 9830 4780
rect 10594 4768 10600 4780
rect 10652 4768 10658 4820
rect 11974 4808 11980 4820
rect 11935 4780 11980 4808
rect 11974 4768 11980 4780
rect 12032 4768 12038 4820
rect 13722 4768 13728 4820
rect 13780 4808 13786 4820
rect 14461 4811 14519 4817
rect 14461 4808 14473 4811
rect 13780 4780 14473 4808
rect 13780 4768 13786 4780
rect 14461 4777 14473 4780
rect 14507 4777 14519 4811
rect 14461 4771 14519 4777
rect 14921 4811 14979 4817
rect 14921 4777 14933 4811
rect 14967 4808 14979 4811
rect 17954 4808 17960 4820
rect 14967 4780 17960 4808
rect 14967 4777 14979 4780
rect 14921 4771 14979 4777
rect 17954 4768 17960 4780
rect 18012 4768 18018 4820
rect 18230 4808 18236 4820
rect 18143 4780 18236 4808
rect 18230 4768 18236 4780
rect 18288 4808 18294 4820
rect 20625 4811 20683 4817
rect 20625 4808 20637 4811
rect 18288 4780 20637 4808
rect 18288 4768 18294 4780
rect 20625 4777 20637 4780
rect 20671 4777 20683 4811
rect 20625 4771 20683 4777
rect 22094 4768 22100 4820
rect 22152 4808 22158 4820
rect 23477 4811 23535 4817
rect 22152 4780 22508 4808
rect 22152 4768 22158 4780
rect 1581 4743 1639 4749
rect 1581 4709 1593 4743
rect 1627 4740 1639 4743
rect 2774 4740 2780 4752
rect 1627 4712 2780 4740
rect 1627 4709 1639 4712
rect 1581 4703 1639 4709
rect 2774 4700 2780 4712
rect 2832 4700 2838 4752
rect 6457 4743 6515 4749
rect 6457 4709 6469 4743
rect 6503 4740 6515 4743
rect 6638 4740 6644 4752
rect 6503 4712 6644 4740
rect 6503 4709 6515 4712
rect 6457 4703 6515 4709
rect 6638 4700 6644 4712
rect 6696 4700 6702 4752
rect 10042 4740 10048 4752
rect 9324 4712 10048 4740
rect 2314 4632 2320 4684
rect 2372 4672 2378 4684
rect 2593 4675 2651 4681
rect 2593 4672 2605 4675
rect 2372 4644 2605 4672
rect 2372 4632 2378 4644
rect 2593 4641 2605 4644
rect 2639 4641 2651 4675
rect 7466 4672 7472 4684
rect 7427 4644 7472 4672
rect 2593 4635 2651 4641
rect 7466 4632 7472 4644
rect 7524 4632 7530 4684
rect 1394 4604 1400 4616
rect 1355 4576 1400 4604
rect 1394 4564 1400 4576
rect 1452 4564 1458 4616
rect 3789 4607 3847 4613
rect 3789 4573 3801 4607
rect 3835 4604 3847 4607
rect 3878 4604 3884 4616
rect 3835 4576 3884 4604
rect 3835 4573 3847 4576
rect 3789 4567 3847 4573
rect 3878 4564 3884 4576
rect 3936 4564 3942 4616
rect 4706 4613 4712 4616
rect 4433 4607 4491 4613
rect 4433 4573 4445 4607
rect 4479 4573 4491 4607
rect 4700 4604 4712 4613
rect 4667 4576 4712 4604
rect 4433 4567 4491 4573
rect 4700 4567 4712 4576
rect 2501 4539 2559 4545
rect 2501 4505 2513 4539
rect 2547 4536 2559 4539
rect 4246 4536 4252 4548
rect 2547 4508 4252 4536
rect 2547 4505 2559 4508
rect 2501 4499 2559 4505
rect 4246 4496 4252 4508
rect 4304 4496 4310 4548
rect 4448 4536 4476 4567
rect 4706 4564 4712 4567
rect 4764 4564 4770 4616
rect 8202 4604 8208 4616
rect 8163 4576 8208 4604
rect 8202 4564 8208 4576
rect 8260 4564 8266 4616
rect 8938 4604 8944 4616
rect 8899 4576 8944 4604
rect 8938 4564 8944 4576
rect 8996 4564 9002 4616
rect 9324 4613 9352 4712
rect 10042 4700 10048 4712
rect 10100 4700 10106 4752
rect 11698 4749 11704 4752
rect 11682 4743 11704 4749
rect 11682 4709 11694 4743
rect 11682 4703 11704 4709
rect 11698 4700 11704 4703
rect 11756 4700 11762 4752
rect 11790 4700 11796 4752
rect 11848 4740 11854 4752
rect 12066 4740 12072 4752
rect 11848 4712 11893 4740
rect 11992 4712 12072 4740
rect 11848 4700 11854 4712
rect 10321 4675 10379 4681
rect 10321 4672 10333 4675
rect 9508 4644 10333 4672
rect 9508 4616 9536 4644
rect 10321 4641 10333 4644
rect 10367 4641 10379 4675
rect 10321 4635 10379 4641
rect 11885 4675 11943 4681
rect 11885 4641 11897 4675
rect 11931 4672 11943 4675
rect 11992 4672 12020 4712
rect 12066 4700 12072 4712
rect 12124 4700 12130 4752
rect 12526 4700 12532 4752
rect 12584 4740 12590 4752
rect 13446 4740 13452 4752
rect 12584 4712 13452 4740
rect 12584 4700 12590 4712
rect 13446 4700 13452 4712
rect 13504 4740 13510 4752
rect 13814 4740 13820 4752
rect 13504 4712 13820 4740
rect 13504 4700 13510 4712
rect 13814 4700 13820 4712
rect 13872 4700 13878 4752
rect 14090 4740 14096 4752
rect 14051 4712 14096 4740
rect 14090 4700 14096 4712
rect 14148 4700 14154 4752
rect 14553 4743 14611 4749
rect 14553 4709 14565 4743
rect 14599 4709 14611 4743
rect 18138 4740 18144 4752
rect 14553 4703 14611 4709
rect 16040 4712 18144 4740
rect 11931 4644 12020 4672
rect 12084 4644 13032 4672
rect 11931 4641 11943 4644
rect 11885 4635 11943 4641
rect 9309 4607 9367 4613
rect 9309 4573 9321 4607
rect 9355 4573 9367 4607
rect 9490 4604 9496 4616
rect 9451 4576 9496 4604
rect 9309 4567 9367 4573
rect 9490 4564 9496 4576
rect 9548 4564 9554 4616
rect 10042 4564 10048 4616
rect 10100 4604 10106 4616
rect 10229 4607 10287 4613
rect 10229 4604 10241 4607
rect 10100 4576 10241 4604
rect 10100 4564 10106 4576
rect 10229 4573 10241 4576
rect 10275 4604 10287 4607
rect 12084 4604 12112 4644
rect 10275 4576 12112 4604
rect 10275 4573 10287 4576
rect 10229 4567 10287 4573
rect 12434 4564 12440 4616
rect 12492 4604 12498 4616
rect 13004 4613 13032 4644
rect 13630 4632 13636 4684
rect 13688 4672 13694 4684
rect 14568 4672 14596 4703
rect 16040 4684 16068 4712
rect 13688 4644 14596 4672
rect 14645 4675 14703 4681
rect 13688 4632 13694 4644
rect 14645 4641 14657 4675
rect 14691 4672 14703 4675
rect 14734 4672 14740 4684
rect 14691 4644 14740 4672
rect 14691 4641 14703 4644
rect 14645 4635 14703 4641
rect 12713 4607 12771 4613
rect 12713 4604 12725 4607
rect 12492 4576 12725 4604
rect 12492 4564 12498 4576
rect 12713 4573 12725 4576
rect 12759 4573 12771 4607
rect 12713 4567 12771 4573
rect 12989 4607 13047 4613
rect 12989 4573 13001 4607
rect 13035 4604 13047 4607
rect 13906 4604 13912 4616
rect 13035 4576 13912 4604
rect 13035 4573 13047 4576
rect 12989 4567 13047 4573
rect 4614 4536 4620 4548
rect 4448 4508 4620 4536
rect 4614 4496 4620 4508
rect 4672 4496 4678 4548
rect 6641 4539 6699 4545
rect 6641 4505 6653 4539
rect 6687 4536 6699 4539
rect 7285 4539 7343 4545
rect 7285 4536 7297 4539
rect 6687 4508 7297 4536
rect 6687 4505 6699 4508
rect 6641 4499 6699 4505
rect 7285 4505 7297 4508
rect 7331 4536 7343 4539
rect 7834 4536 7840 4548
rect 7331 4508 7840 4536
rect 7331 4505 7343 4508
rect 7285 4499 7343 4505
rect 7834 4496 7840 4508
rect 7892 4496 7898 4548
rect 9030 4496 9036 4548
rect 9088 4536 9094 4548
rect 10689 4539 10747 4545
rect 10689 4536 10701 4539
rect 9088 4508 10701 4536
rect 9088 4496 9094 4508
rect 10689 4505 10701 4508
rect 10735 4505 10747 4539
rect 10689 4499 10747 4505
rect 11146 4496 11152 4548
rect 11204 4536 11210 4548
rect 11517 4539 11575 4545
rect 11517 4536 11529 4539
rect 11204 4508 11529 4536
rect 11204 4496 11210 4508
rect 11517 4505 11529 4508
rect 11563 4505 11575 4539
rect 11517 4499 11575 4505
rect 11974 4496 11980 4548
rect 12032 4536 12038 4548
rect 12728 4536 12756 4567
rect 13906 4564 13912 4576
rect 13964 4564 13970 4616
rect 14458 4564 14464 4616
rect 14516 4604 14522 4616
rect 14660 4604 14688 4635
rect 14734 4632 14740 4644
rect 14792 4632 14798 4684
rect 15930 4672 15936 4684
rect 15891 4644 15936 4672
rect 15930 4632 15936 4644
rect 15988 4632 15994 4684
rect 16022 4632 16028 4684
rect 16080 4672 16086 4684
rect 16853 4675 16911 4681
rect 16080 4644 16125 4672
rect 16080 4632 16086 4644
rect 16853 4641 16865 4675
rect 16899 4672 16911 4675
rect 17954 4672 17960 4684
rect 16899 4644 17960 4672
rect 16899 4641 16911 4644
rect 16853 4635 16911 4641
rect 17954 4632 17960 4644
rect 18012 4632 18018 4684
rect 18064 4681 18092 4712
rect 18138 4700 18144 4712
rect 18196 4700 18202 4752
rect 18248 4681 18276 4768
rect 18690 4740 18696 4752
rect 18651 4712 18696 4740
rect 18690 4700 18696 4712
rect 18748 4700 18754 4752
rect 20254 4700 20260 4752
rect 20312 4740 20318 4752
rect 21085 4743 21143 4749
rect 21085 4740 21097 4743
rect 20312 4712 21097 4740
rect 20312 4700 20318 4712
rect 21085 4709 21097 4712
rect 21131 4709 21143 4743
rect 21085 4703 21143 4709
rect 22480 4681 22508 4780
rect 23477 4777 23489 4811
rect 23523 4808 23535 4811
rect 23750 4808 23756 4820
rect 23523 4780 23756 4808
rect 23523 4777 23535 4780
rect 23477 4771 23535 4777
rect 23750 4768 23756 4780
rect 23808 4768 23814 4820
rect 27154 4808 27160 4820
rect 27115 4780 27160 4808
rect 27154 4768 27160 4780
rect 27212 4768 27218 4820
rect 27338 4768 27344 4820
rect 27396 4808 27402 4820
rect 27617 4811 27675 4817
rect 27617 4808 27629 4811
rect 27396 4780 27629 4808
rect 27396 4768 27402 4780
rect 27617 4777 27629 4780
rect 27663 4777 27675 4811
rect 27617 4771 27675 4777
rect 32769 4811 32827 4817
rect 32769 4777 32781 4811
rect 32815 4808 32827 4811
rect 33318 4808 33324 4820
rect 32815 4780 33324 4808
rect 32815 4777 32827 4780
rect 32769 4771 32827 4777
rect 33318 4768 33324 4780
rect 33376 4768 33382 4820
rect 33870 4808 33876 4820
rect 33831 4780 33876 4808
rect 33870 4768 33876 4780
rect 33928 4768 33934 4820
rect 34422 4768 34428 4820
rect 34480 4808 34486 4820
rect 34701 4811 34759 4817
rect 34701 4808 34713 4811
rect 34480 4780 34713 4808
rect 34480 4768 34486 4780
rect 34701 4777 34713 4780
rect 34747 4777 34759 4811
rect 34701 4771 34759 4777
rect 36173 4811 36231 4817
rect 36173 4777 36185 4811
rect 36219 4808 36231 4811
rect 36262 4808 36268 4820
rect 36219 4780 36268 4808
rect 36219 4777 36231 4780
rect 36173 4771 36231 4777
rect 36262 4768 36268 4780
rect 36320 4768 36326 4820
rect 37369 4811 37427 4817
rect 37369 4777 37381 4811
rect 37415 4808 37427 4811
rect 37458 4808 37464 4820
rect 37415 4780 37464 4808
rect 37415 4777 37427 4780
rect 37369 4771 37427 4777
rect 37458 4768 37464 4780
rect 37516 4768 37522 4820
rect 22738 4700 22744 4752
rect 22796 4740 22802 4752
rect 25225 4743 25283 4749
rect 25225 4740 25237 4743
rect 22796 4712 25237 4740
rect 22796 4700 22802 4712
rect 25225 4709 25237 4712
rect 25271 4740 25283 4743
rect 25590 4740 25596 4752
rect 25271 4712 25596 4740
rect 25271 4709 25283 4712
rect 25225 4703 25283 4709
rect 25590 4700 25596 4712
rect 25648 4700 25654 4752
rect 57238 4700 57244 4752
rect 57296 4740 57302 4752
rect 57885 4743 57943 4749
rect 57885 4740 57897 4743
rect 57296 4712 57897 4740
rect 57296 4700 57302 4712
rect 57885 4709 57897 4712
rect 57931 4709 57943 4743
rect 57885 4703 57943 4709
rect 58250 4700 58256 4752
rect 58308 4740 58314 4752
rect 59173 4743 59231 4749
rect 59173 4740 59185 4743
rect 58308 4712 59185 4740
rect 58308 4700 58314 4712
rect 59173 4709 59185 4712
rect 59219 4709 59231 4743
rect 59173 4703 59231 4709
rect 18049 4675 18107 4681
rect 18049 4641 18061 4675
rect 18095 4641 18107 4675
rect 18049 4635 18107 4641
rect 18233 4675 18291 4681
rect 18233 4641 18245 4675
rect 18279 4641 18291 4675
rect 18233 4635 18291 4641
rect 22465 4675 22523 4681
rect 22465 4641 22477 4675
rect 22511 4672 22523 4675
rect 24302 4672 24308 4684
rect 22511 4644 24308 4672
rect 22511 4641 22523 4644
rect 22465 4635 22523 4641
rect 24302 4632 24308 4644
rect 24360 4672 24366 4684
rect 25777 4675 25835 4681
rect 25777 4672 25789 4675
rect 24360 4644 25789 4672
rect 24360 4632 24366 4644
rect 25777 4641 25789 4644
rect 25823 4641 25835 4675
rect 28994 4672 29000 4684
rect 28955 4644 29000 4672
rect 25777 4635 25835 4641
rect 28994 4632 29000 4644
rect 29052 4632 29058 4684
rect 38746 4672 38752 4684
rect 38707 4644 38752 4672
rect 38746 4632 38752 4644
rect 38804 4632 38810 4684
rect 58894 4632 58900 4684
rect 58952 4672 58958 4684
rect 60461 4675 60519 4681
rect 60461 4672 60473 4675
rect 58952 4644 60473 4672
rect 58952 4632 58958 4644
rect 60461 4641 60473 4644
rect 60507 4641 60519 4675
rect 60461 4635 60519 4641
rect 14516 4576 14688 4604
rect 17497 4607 17555 4613
rect 14516 4564 14522 4576
rect 17497 4573 17509 4607
rect 17543 4604 17555 4607
rect 19150 4604 19156 4616
rect 17543 4576 19156 4604
rect 17543 4573 17555 4576
rect 17497 4567 17555 4573
rect 19150 4564 19156 4576
rect 19208 4564 19214 4616
rect 19245 4607 19303 4613
rect 19245 4573 19257 4607
rect 19291 4573 19303 4607
rect 19245 4567 19303 4573
rect 13630 4536 13636 4548
rect 12032 4508 12664 4536
rect 12728 4508 13636 4536
rect 12032 4496 12038 4508
rect 1946 4428 1952 4480
rect 2004 4468 2010 4480
rect 2041 4471 2099 4477
rect 2041 4468 2053 4471
rect 2004 4440 2053 4468
rect 2004 4428 2010 4440
rect 2041 4437 2053 4440
rect 2087 4437 2099 4471
rect 2406 4468 2412 4480
rect 2367 4440 2412 4468
rect 2041 4431 2099 4437
rect 2406 4428 2412 4440
rect 2464 4468 2470 4480
rect 2682 4468 2688 4480
rect 2464 4440 2688 4468
rect 2464 4428 2470 4440
rect 2682 4428 2688 4440
rect 2740 4428 2746 4480
rect 3973 4471 4031 4477
rect 3973 4437 3985 4471
rect 4019 4468 4031 4471
rect 4706 4468 4712 4480
rect 4019 4440 4712 4468
rect 4019 4437 4031 4440
rect 3973 4431 4031 4437
rect 4706 4428 4712 4440
rect 4764 4428 4770 4480
rect 8386 4468 8392 4480
rect 8347 4440 8392 4468
rect 8386 4428 8392 4440
rect 8444 4428 8450 4480
rect 9125 4471 9183 4477
rect 9125 4437 9137 4471
rect 9171 4468 9183 4471
rect 9306 4468 9312 4480
rect 9171 4440 9312 4468
rect 9171 4437 9183 4440
rect 9125 4431 9183 4437
rect 9306 4428 9312 4440
rect 9364 4428 9370 4480
rect 10045 4471 10103 4477
rect 10045 4437 10057 4471
rect 10091 4468 10103 4471
rect 10134 4468 10140 4480
rect 10091 4440 10140 4468
rect 10091 4437 10103 4440
rect 10045 4431 10103 4437
rect 10134 4428 10140 4440
rect 10192 4428 10198 4480
rect 10318 4428 10324 4480
rect 10376 4468 10382 4480
rect 12526 4468 12532 4480
rect 10376 4440 12532 4468
rect 10376 4428 10382 4440
rect 12526 4428 12532 4440
rect 12584 4428 12590 4480
rect 12636 4468 12664 4508
rect 13630 4496 13636 4508
rect 13688 4496 13694 4548
rect 15396 4508 18000 4536
rect 15396 4468 15424 4508
rect 12636 4440 15424 4468
rect 15473 4471 15531 4477
rect 15473 4437 15485 4471
rect 15519 4468 15531 4471
rect 15562 4468 15568 4480
rect 15519 4440 15568 4468
rect 15519 4437 15531 4440
rect 15473 4431 15531 4437
rect 15562 4428 15568 4440
rect 15620 4428 15626 4480
rect 15838 4468 15844 4480
rect 15799 4440 15844 4468
rect 15838 4428 15844 4440
rect 15896 4428 15902 4480
rect 17972 4468 18000 4508
rect 18046 4496 18052 4548
rect 18104 4536 18110 4548
rect 19260 4536 19288 4567
rect 19978 4564 19984 4616
rect 20036 4604 20042 4616
rect 22198 4607 22256 4613
rect 22198 4604 22210 4607
rect 20036 4576 22210 4604
rect 20036 4564 20042 4576
rect 22198 4573 22210 4576
rect 22244 4573 22256 4607
rect 22198 4567 22256 4573
rect 23014 4564 23020 4616
rect 23072 4604 23078 4616
rect 23109 4607 23167 4613
rect 23109 4604 23121 4607
rect 23072 4576 23121 4604
rect 23072 4564 23078 4576
rect 23109 4573 23121 4576
rect 23155 4573 23167 4607
rect 23109 4567 23167 4573
rect 23293 4607 23351 4613
rect 23293 4573 23305 4607
rect 23339 4604 23351 4607
rect 23474 4604 23480 4616
rect 23339 4576 23480 4604
rect 23339 4573 23351 4576
rect 23293 4567 23351 4573
rect 23474 4564 23480 4576
rect 23532 4564 23538 4616
rect 25222 4564 25228 4616
rect 25280 4604 25286 4616
rect 26033 4607 26091 4613
rect 26033 4604 26045 4607
rect 25280 4576 26045 4604
rect 25280 4564 25286 4576
rect 26033 4573 26045 4576
rect 26079 4573 26091 4607
rect 26033 4567 26091 4573
rect 32398 4564 32404 4616
rect 32456 4604 32462 4616
rect 32953 4607 33011 4613
rect 32953 4604 32965 4607
rect 32456 4576 32965 4604
rect 32456 4564 32462 4576
rect 32953 4573 32965 4576
rect 32999 4573 33011 4607
rect 32953 4567 33011 4573
rect 34790 4564 34796 4616
rect 34848 4604 34854 4616
rect 34885 4607 34943 4613
rect 34885 4604 34897 4607
rect 34848 4576 34897 4604
rect 34848 4564 34854 4576
rect 34885 4573 34897 4576
rect 34931 4573 34943 4607
rect 34885 4567 34943 4573
rect 35989 4607 36047 4613
rect 35989 4573 36001 4607
rect 36035 4604 36047 4607
rect 36078 4604 36084 4616
rect 36035 4576 36084 4604
rect 36035 4573 36047 4576
rect 35989 4567 36047 4573
rect 36078 4564 36084 4576
rect 36136 4564 36142 4616
rect 37734 4564 37740 4616
rect 37792 4604 37798 4616
rect 38482 4607 38540 4613
rect 38482 4604 38494 4607
rect 37792 4576 38494 4604
rect 37792 4564 37798 4576
rect 38482 4573 38494 4576
rect 38528 4573 38540 4607
rect 38482 4567 38540 4573
rect 57146 4564 57152 4616
rect 57204 4604 57210 4616
rect 57241 4607 57299 4613
rect 57241 4604 57253 4607
rect 57204 4576 57253 4604
rect 57204 4564 57210 4576
rect 57241 4573 57253 4576
rect 57287 4573 57299 4607
rect 57241 4567 57299 4573
rect 57606 4564 57612 4616
rect 57664 4604 57670 4616
rect 58529 4607 58587 4613
rect 58529 4604 58541 4607
rect 57664 4576 58541 4604
rect 57664 4564 57670 4576
rect 58529 4573 58541 4576
rect 58575 4573 58587 4607
rect 58529 4567 58587 4573
rect 18104 4508 19288 4536
rect 19512 4539 19570 4545
rect 18104 4496 18110 4508
rect 19512 4505 19524 4539
rect 19558 4505 19570 4539
rect 19512 4499 19570 4505
rect 18230 4468 18236 4480
rect 17972 4440 18236 4468
rect 18230 4428 18236 4440
rect 18288 4428 18294 4480
rect 18325 4471 18383 4477
rect 18325 4437 18337 4471
rect 18371 4468 18383 4471
rect 18874 4468 18880 4480
rect 18371 4440 18880 4468
rect 18371 4437 18383 4440
rect 18325 4431 18383 4437
rect 18874 4428 18880 4440
rect 18932 4428 18938 4480
rect 19426 4428 19432 4480
rect 19484 4468 19490 4480
rect 19536 4468 19564 4499
rect 21266 4496 21272 4548
rect 21324 4536 21330 4548
rect 24397 4539 24455 4545
rect 24397 4536 24409 4539
rect 21324 4508 24409 4536
rect 21324 4496 21330 4508
rect 24397 4505 24409 4508
rect 24443 4536 24455 4539
rect 24946 4536 24952 4548
rect 24443 4508 24952 4536
rect 24443 4505 24455 4508
rect 24397 4499 24455 4505
rect 24946 4496 24952 4508
rect 25004 4496 25010 4548
rect 27706 4496 27712 4548
rect 27764 4536 27770 4548
rect 28730 4539 28788 4545
rect 28730 4536 28742 4539
rect 27764 4508 28742 4536
rect 27764 4496 27770 4508
rect 28730 4505 28742 4508
rect 28776 4505 28788 4539
rect 28730 4499 28788 4505
rect 33137 4539 33195 4545
rect 33137 4505 33149 4539
rect 33183 4536 33195 4539
rect 34698 4536 34704 4548
rect 33183 4508 34704 4536
rect 33183 4505 33195 4508
rect 33137 4499 33195 4505
rect 34698 4496 34704 4508
rect 34756 4536 34762 4548
rect 35069 4539 35127 4545
rect 35069 4536 35081 4539
rect 34756 4508 35081 4536
rect 34756 4496 34762 4508
rect 35069 4505 35081 4508
rect 35115 4536 35127 4539
rect 35805 4539 35863 4545
rect 35805 4536 35817 4539
rect 35115 4508 35817 4536
rect 35115 4505 35127 4508
rect 35069 4499 35127 4505
rect 35805 4505 35817 4508
rect 35851 4505 35863 4539
rect 35805 4499 35863 4505
rect 19484 4440 19564 4468
rect 19484 4428 19490 4440
rect 1104 4378 68816 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 68816 4378
rect 1104 4304 68816 4326
rect 2133 4267 2191 4273
rect 2133 4233 2145 4267
rect 2179 4264 2191 4267
rect 2222 4264 2228 4276
rect 2179 4236 2228 4264
rect 2179 4233 2191 4236
rect 2133 4227 2191 4233
rect 2222 4224 2228 4236
rect 2280 4224 2286 4276
rect 5169 4267 5227 4273
rect 5169 4233 5181 4267
rect 5215 4233 5227 4267
rect 5169 4227 5227 4233
rect 7561 4267 7619 4273
rect 7561 4233 7573 4267
rect 7607 4264 7619 4267
rect 8662 4264 8668 4276
rect 7607 4236 8668 4264
rect 7607 4233 7619 4236
rect 7561 4227 7619 4233
rect 2958 4156 2964 4208
rect 3016 4196 3022 4208
rect 3114 4199 3172 4205
rect 3114 4196 3126 4199
rect 3016 4168 3126 4196
rect 3016 4156 3022 4168
rect 3114 4165 3126 4168
rect 3160 4165 3172 4199
rect 5184 4196 5212 4227
rect 8662 4224 8668 4236
rect 8720 4264 8726 4276
rect 9398 4264 9404 4276
rect 8720 4236 9404 4264
rect 8720 4224 8726 4236
rect 9398 4224 9404 4236
rect 9456 4224 9462 4276
rect 9490 4224 9496 4276
rect 9548 4264 9554 4276
rect 9585 4267 9643 4273
rect 9585 4264 9597 4267
rect 9548 4236 9597 4264
rect 9548 4224 9554 4236
rect 9585 4233 9597 4236
rect 9631 4233 9643 4267
rect 10594 4264 10600 4276
rect 10555 4236 10600 4264
rect 9585 4227 9643 4233
rect 10594 4224 10600 4236
rect 10652 4224 10658 4276
rect 12066 4264 12072 4276
rect 10796 4236 12072 4264
rect 5184 4168 6684 4196
rect 3114 4159 3172 4165
rect 1946 4128 1952 4140
rect 1907 4100 1952 4128
rect 1946 4088 1952 4100
rect 2004 4088 2010 4140
rect 3694 4128 3700 4140
rect 2746 4100 3700 4128
rect 1762 4060 1768 4072
rect 1675 4032 1768 4060
rect 1762 4020 1768 4032
rect 1820 4020 1826 4072
rect 1780 3924 1808 4020
rect 1946 3924 1952 3936
rect 1780 3896 1952 3924
rect 1946 3884 1952 3896
rect 2004 3924 2010 3936
rect 2746 3924 2774 4100
rect 3694 4088 3700 4100
rect 3752 4088 3758 4140
rect 4985 4131 5043 4137
rect 4985 4097 4997 4131
rect 5031 4128 5043 4131
rect 5074 4128 5080 4140
rect 5031 4100 5080 4128
rect 5031 4097 5043 4100
rect 4985 4091 5043 4097
rect 5074 4088 5080 4100
rect 5132 4088 5138 4140
rect 5626 4128 5632 4140
rect 5587 4100 5632 4128
rect 5626 4088 5632 4100
rect 5684 4088 5690 4140
rect 6549 4131 6607 4137
rect 6549 4097 6561 4131
rect 6595 4097 6607 4131
rect 6656 4128 6684 4168
rect 8202 4156 8208 4208
rect 8260 4196 8266 4208
rect 10318 4196 10324 4208
rect 8260 4168 10324 4196
rect 8260 4156 8266 4168
rect 10318 4156 10324 4168
rect 10376 4156 10382 4208
rect 7653 4131 7711 4137
rect 6656 4100 7604 4128
rect 6549 4091 6607 4097
rect 2866 4020 2872 4072
rect 2924 4060 2930 4072
rect 2924 4032 2969 4060
rect 2924 4020 2930 4032
rect 6365 3995 6423 4001
rect 6365 3992 6377 3995
rect 3804 3964 6377 3992
rect 2004 3896 2774 3924
rect 2004 3884 2010 3896
rect 3050 3884 3056 3936
rect 3108 3924 3114 3936
rect 3804 3924 3832 3964
rect 6365 3961 6377 3964
rect 6411 3961 6423 3995
rect 6564 3992 6592 4091
rect 6730 4060 6736 4072
rect 6691 4032 6736 4060
rect 6730 4020 6736 4032
rect 6788 4020 6794 4072
rect 7193 3995 7251 4001
rect 7193 3992 7205 3995
rect 6564 3964 7205 3992
rect 6365 3955 6423 3961
rect 7193 3961 7205 3964
rect 7239 3961 7251 3995
rect 7576 3992 7604 4100
rect 7653 4097 7665 4131
rect 7699 4128 7711 4131
rect 8018 4128 8024 4140
rect 7699 4100 8024 4128
rect 7699 4097 7711 4100
rect 7653 4091 7711 4097
rect 8018 4088 8024 4100
rect 8076 4088 8082 4140
rect 8294 4088 8300 4140
rect 8352 4128 8358 4140
rect 8849 4131 8907 4137
rect 8849 4128 8861 4131
rect 8352 4100 8861 4128
rect 8352 4088 8358 4100
rect 8849 4097 8861 4100
rect 8895 4097 8907 4131
rect 9122 4128 9128 4140
rect 9083 4100 9128 4128
rect 8849 4091 8907 4097
rect 9122 4088 9128 4100
rect 9180 4088 9186 4140
rect 9766 4128 9772 4140
rect 9727 4100 9772 4128
rect 9766 4088 9772 4100
rect 9824 4088 9830 4140
rect 10686 4088 10692 4140
rect 10744 4128 10750 4140
rect 10796 4137 10824 4236
rect 12066 4224 12072 4236
rect 12124 4224 12130 4276
rect 13262 4224 13268 4276
rect 13320 4264 13326 4276
rect 14366 4264 14372 4276
rect 13320 4236 14372 4264
rect 13320 4224 13326 4236
rect 14366 4224 14372 4236
rect 14424 4224 14430 4276
rect 16206 4224 16212 4276
rect 16264 4264 16270 4276
rect 18138 4264 18144 4276
rect 16264 4236 18144 4264
rect 16264 4224 16270 4236
rect 18138 4224 18144 4236
rect 18196 4224 18202 4276
rect 18230 4224 18236 4276
rect 18288 4264 18294 4276
rect 18598 4264 18604 4276
rect 18288 4236 18604 4264
rect 18288 4224 18294 4236
rect 18598 4224 18604 4236
rect 18656 4224 18662 4276
rect 19426 4224 19432 4276
rect 19484 4264 19490 4276
rect 19521 4267 19579 4273
rect 19521 4264 19533 4267
rect 19484 4236 19533 4264
rect 19484 4224 19490 4236
rect 19521 4233 19533 4236
rect 19567 4233 19579 4267
rect 19521 4227 19579 4233
rect 20073 4267 20131 4273
rect 20073 4233 20085 4267
rect 20119 4264 20131 4267
rect 20438 4264 20444 4276
rect 20119 4236 20444 4264
rect 20119 4233 20131 4236
rect 20073 4227 20131 4233
rect 20438 4224 20444 4236
rect 20496 4224 20502 4276
rect 23382 4224 23388 4276
rect 23440 4264 23446 4276
rect 23440 4236 23507 4264
rect 23440 4224 23446 4236
rect 10965 4199 11023 4205
rect 10965 4165 10977 4199
rect 11011 4196 11023 4199
rect 11698 4196 11704 4208
rect 11011 4168 11704 4196
rect 11011 4165 11023 4168
rect 10965 4159 11023 4165
rect 11698 4156 11704 4168
rect 11756 4196 11762 4208
rect 11882 4196 11888 4208
rect 11756 4168 11888 4196
rect 11756 4156 11762 4168
rect 11882 4156 11888 4168
rect 11940 4156 11946 4208
rect 12342 4156 12348 4208
rect 12400 4156 12406 4208
rect 15102 4156 15108 4208
rect 15160 4156 15166 4208
rect 17954 4156 17960 4208
rect 18012 4196 18018 4208
rect 19058 4196 19064 4208
rect 18012 4168 19064 4196
rect 18012 4156 18018 4168
rect 19058 4156 19064 4168
rect 19116 4156 19122 4208
rect 10781 4131 10839 4137
rect 10781 4128 10793 4131
rect 10744 4100 10793 4128
rect 10744 4088 10750 4100
rect 10781 4097 10793 4100
rect 10827 4097 10839 4131
rect 12360 4128 12388 4156
rect 13722 4128 13728 4140
rect 10781 4091 10839 4097
rect 10980 4100 13728 4128
rect 7834 4060 7840 4072
rect 7795 4032 7840 4060
rect 7834 4020 7840 4032
rect 7892 4020 7898 4072
rect 9306 4020 9312 4072
rect 9364 4060 9370 4072
rect 9953 4063 10011 4069
rect 9953 4060 9965 4063
rect 9364 4032 9965 4060
rect 9364 4020 9370 4032
rect 9953 4029 9965 4032
rect 9999 4060 10011 4063
rect 10980 4060 11008 4100
rect 13722 4088 13728 4100
rect 13780 4088 13786 4140
rect 14369 4131 14427 4137
rect 14369 4097 14381 4131
rect 14415 4128 14427 4131
rect 15120 4128 15148 4156
rect 23479 4143 23507 4236
rect 34790 4224 34796 4276
rect 34848 4264 34854 4276
rect 34885 4267 34943 4273
rect 34885 4264 34897 4267
rect 34848 4236 34897 4264
rect 34848 4224 34854 4236
rect 34885 4233 34897 4236
rect 34931 4233 34943 4267
rect 34885 4227 34943 4233
rect 36078 4224 36084 4276
rect 36136 4264 36142 4276
rect 36725 4267 36783 4273
rect 36725 4264 36737 4267
rect 36136 4236 36737 4264
rect 36136 4224 36142 4236
rect 36725 4233 36737 4236
rect 36771 4233 36783 4267
rect 36725 4227 36783 4233
rect 26786 4156 26792 4208
rect 26844 4196 26850 4208
rect 35894 4196 35900 4208
rect 26844 4168 27660 4196
rect 26844 4156 26850 4168
rect 15378 4128 15384 4140
rect 14415 4100 15148 4128
rect 15339 4100 15384 4128
rect 14415 4097 14427 4100
rect 14369 4091 14427 4097
rect 15378 4088 15384 4100
rect 15436 4088 15442 4140
rect 15562 4128 15568 4140
rect 15523 4100 15568 4128
rect 15562 4088 15568 4100
rect 15620 4088 15626 4140
rect 17770 4088 17776 4140
rect 17828 4137 17834 4140
rect 17828 4128 17840 4137
rect 18046 4128 18052 4140
rect 17828 4100 17873 4128
rect 18007 4100 18052 4128
rect 17828 4091 17840 4100
rect 17828 4088 17834 4091
rect 18046 4088 18052 4100
rect 18104 4088 18110 4140
rect 18690 4128 18696 4140
rect 18651 4100 18696 4128
rect 18690 4088 18696 4100
rect 18748 4088 18754 4140
rect 18877 4131 18935 4137
rect 18877 4097 18889 4131
rect 18923 4128 18935 4131
rect 19337 4131 19395 4137
rect 19337 4128 19349 4131
rect 18923 4100 19349 4128
rect 18923 4097 18935 4100
rect 18877 4091 18935 4097
rect 19337 4097 19349 4100
rect 19383 4097 19395 4131
rect 23198 4128 23204 4140
rect 23159 4100 23204 4128
rect 19337 4091 19395 4097
rect 23198 4088 23204 4100
rect 23256 4088 23262 4140
rect 23364 4137 23422 4143
rect 23364 4134 23376 4137
rect 23308 4106 23376 4134
rect 9999 4032 11008 4060
rect 9999 4029 10011 4032
rect 9953 4023 10011 4029
rect 12066 4020 12072 4072
rect 12124 4060 12130 4072
rect 12342 4060 12348 4072
rect 12124 4032 12348 4060
rect 12124 4020 12130 4032
rect 12342 4020 12348 4032
rect 12400 4020 12406 4072
rect 12713 4063 12771 4069
rect 12713 4029 12725 4063
rect 12759 4060 12771 4063
rect 12802 4060 12808 4072
rect 12759 4032 12808 4060
rect 12759 4029 12771 4032
rect 12713 4023 12771 4029
rect 12802 4020 12808 4032
rect 12860 4020 12866 4072
rect 13446 4060 13452 4072
rect 13407 4032 13452 4060
rect 13446 4020 13452 4032
rect 13504 4020 13510 4072
rect 8202 3992 8208 4004
rect 7576 3964 8208 3992
rect 7193 3955 7251 3961
rect 8202 3952 8208 3964
rect 8260 3952 8266 4004
rect 10686 3992 10692 4004
rect 9048 3964 10692 3992
rect 4246 3924 4252 3936
rect 3108 3896 3832 3924
rect 4207 3896 4252 3924
rect 3108 3884 3114 3896
rect 4246 3884 4252 3896
rect 4304 3884 4310 3936
rect 5813 3927 5871 3933
rect 5813 3893 5825 3927
rect 5859 3924 5871 3927
rect 9048 3924 9076 3964
rect 10686 3952 10692 3964
rect 10744 3952 10750 4004
rect 11238 3992 11244 4004
rect 10888 3964 11244 3992
rect 5859 3896 9076 3924
rect 5859 3893 5871 3896
rect 5813 3887 5871 3893
rect 9122 3884 9128 3936
rect 9180 3924 9186 3936
rect 10888 3924 10916 3964
rect 11238 3952 11244 3964
rect 11296 3952 11302 4004
rect 11790 3992 11796 4004
rect 11751 3964 11796 3992
rect 11790 3952 11796 3964
rect 11848 3952 11854 4004
rect 11882 3952 11888 4004
rect 11940 3992 11946 4004
rect 12253 3995 12311 4001
rect 12253 3992 12265 3995
rect 11940 3964 12265 3992
rect 11940 3952 11946 3964
rect 12253 3961 12265 3964
rect 12299 3961 12311 3995
rect 12253 3955 12311 3961
rect 9180 3896 10916 3924
rect 9180 3884 9186 3896
rect 10962 3884 10968 3936
rect 11020 3924 11026 3936
rect 12066 3924 12072 3936
rect 11020 3896 12072 3924
rect 11020 3884 11026 3896
rect 12066 3884 12072 3896
rect 12124 3884 12130 3936
rect 12158 3884 12164 3936
rect 12216 3924 12222 3936
rect 13740 3924 13768 4088
rect 14001 4063 14059 4069
rect 14001 4029 14013 4063
rect 14047 4060 14059 4063
rect 14090 4060 14096 4072
rect 14047 4032 14096 4060
rect 14047 4029 14059 4032
rect 14001 4023 14059 4029
rect 14090 4020 14096 4032
rect 14148 4020 14154 4072
rect 15102 4020 15108 4072
rect 15160 4060 15166 4072
rect 15749 4063 15807 4069
rect 15749 4060 15761 4063
rect 15160 4032 15761 4060
rect 15160 4020 15166 4032
rect 15749 4029 15761 4032
rect 15795 4029 15807 4063
rect 18506 4060 18512 4072
rect 18419 4032 18512 4060
rect 15749 4023 15807 4029
rect 13906 3992 13912 4004
rect 13867 3964 13912 3992
rect 13906 3952 13912 3964
rect 13964 3952 13970 4004
rect 13814 3924 13820 3936
rect 12216 3896 12261 3924
rect 13727 3896 13820 3924
rect 12216 3884 12222 3896
rect 13814 3884 13820 3896
rect 13872 3884 13878 3936
rect 14921 3927 14979 3933
rect 14921 3893 14933 3927
rect 14967 3924 14979 3927
rect 15194 3924 15200 3936
rect 14967 3896 15200 3924
rect 14967 3893 14979 3896
rect 14921 3887 14979 3893
rect 15194 3884 15200 3896
rect 15252 3884 15258 3936
rect 15764 3924 15792 4023
rect 18506 4020 18512 4032
rect 18564 4020 18570 4072
rect 18598 4020 18604 4072
rect 18656 4060 18662 4072
rect 20162 4060 20168 4072
rect 18656 4032 20168 4060
rect 18656 4020 18662 4032
rect 20162 4020 20168 4032
rect 20220 4020 20226 4072
rect 23106 4020 23112 4072
rect 23164 4060 23170 4072
rect 23308 4060 23336 4106
rect 23364 4103 23376 4106
rect 23410 4103 23422 4137
rect 23364 4097 23422 4103
rect 23464 4137 23522 4143
rect 23658 4137 23664 4140
rect 23464 4103 23476 4137
rect 23510 4103 23522 4137
rect 23464 4097 23522 4103
rect 23615 4131 23664 4137
rect 23615 4097 23627 4131
rect 23661 4097 23664 4131
rect 23615 4091 23664 4097
rect 23658 4088 23664 4091
rect 23716 4128 23722 4140
rect 24302 4128 24308 4140
rect 23716 4100 23806 4128
rect 24263 4100 24308 4128
rect 23716 4088 23722 4100
rect 24302 4088 24308 4100
rect 24360 4088 24366 4140
rect 24561 4131 24619 4137
rect 24561 4128 24573 4131
rect 24412 4100 24573 4128
rect 23164 4032 23336 4060
rect 23164 4020 23170 4032
rect 15930 3952 15936 4004
rect 15988 3992 15994 4004
rect 16669 3995 16727 4001
rect 16669 3992 16681 3995
rect 15988 3964 16681 3992
rect 15988 3952 15994 3964
rect 16669 3961 16681 3964
rect 16715 3961 16727 3995
rect 16669 3955 16727 3961
rect 18524 3924 18552 4020
rect 18690 3952 18696 4004
rect 18748 3992 18754 4004
rect 18966 3992 18972 4004
rect 18748 3964 18972 3992
rect 18748 3952 18754 3964
rect 18966 3952 18972 3964
rect 19024 3952 19030 4004
rect 20254 3952 20260 4004
rect 20312 3992 20318 4004
rect 21821 3995 21879 4001
rect 21821 3992 21833 3995
rect 20312 3964 21833 3992
rect 20312 3952 20318 3964
rect 21821 3961 21833 3964
rect 21867 3961 21879 3995
rect 23673 3992 23701 4088
rect 23845 4063 23903 4069
rect 23845 4029 23857 4063
rect 23891 4060 23903 4063
rect 24412 4060 24440 4100
rect 24561 4097 24573 4100
rect 24607 4097 24619 4131
rect 27338 4128 27344 4140
rect 27299 4100 27344 4128
rect 24561 4091 24619 4097
rect 27338 4088 27344 4100
rect 27396 4088 27402 4140
rect 27522 4128 27528 4140
rect 27483 4100 27528 4128
rect 27522 4088 27528 4100
rect 27580 4088 27586 4140
rect 27632 4137 27660 4168
rect 33704 4168 34008 4196
rect 27617 4131 27675 4137
rect 27617 4097 27629 4131
rect 27663 4097 27675 4131
rect 27617 4091 27675 4097
rect 27709 4131 27767 4137
rect 27709 4097 27721 4131
rect 27755 4128 27767 4131
rect 27890 4128 27896 4140
rect 27755 4100 27896 4128
rect 27755 4097 27767 4100
rect 27709 4091 27767 4097
rect 27724 4060 27752 4091
rect 27890 4088 27896 4100
rect 27948 4088 27954 4140
rect 30662 4131 30720 4137
rect 30662 4128 30674 4131
rect 28000 4100 30674 4128
rect 28000 4069 28028 4100
rect 30662 4097 30674 4100
rect 30708 4097 30720 4131
rect 30662 4091 30720 4097
rect 30834 4088 30840 4140
rect 30892 4128 30898 4140
rect 30929 4131 30987 4137
rect 30929 4128 30941 4131
rect 30892 4100 30941 4128
rect 30892 4088 30898 4100
rect 30929 4097 30941 4100
rect 30975 4128 30987 4131
rect 33134 4128 33140 4140
rect 30975 4100 33140 4128
rect 30975 4097 30987 4100
rect 30929 4091 30987 4097
rect 33134 4088 33140 4100
rect 33192 4128 33198 4140
rect 33505 4131 33563 4137
rect 33505 4128 33517 4131
rect 33192 4100 33517 4128
rect 33192 4088 33198 4100
rect 33505 4097 33517 4100
rect 33551 4128 33563 4131
rect 33704 4128 33732 4168
rect 33778 4137 33784 4140
rect 33551 4100 33732 4128
rect 33551 4097 33563 4100
rect 33505 4091 33563 4097
rect 33772 4091 33784 4137
rect 33836 4128 33842 4140
rect 33980 4128 34008 4168
rect 35544 4168 35900 4196
rect 35345 4131 35403 4137
rect 35345 4128 35357 4131
rect 33836 4100 33872 4128
rect 33980 4100 35357 4128
rect 33778 4088 33784 4091
rect 33836 4088 33842 4100
rect 35345 4097 35357 4100
rect 35391 4128 35403 4131
rect 35544 4128 35572 4168
rect 35894 4156 35900 4168
rect 35952 4196 35958 4208
rect 38746 4196 38752 4208
rect 35952 4168 38752 4196
rect 35952 4156 35958 4168
rect 38746 4156 38752 4168
rect 38804 4156 38810 4208
rect 35618 4137 35624 4140
rect 35391 4100 35572 4128
rect 35391 4097 35403 4100
rect 35345 4091 35403 4097
rect 35612 4091 35624 4137
rect 35676 4128 35682 4140
rect 35676 4100 35712 4128
rect 35618 4088 35624 4091
rect 35676 4088 35682 4100
rect 57974 4088 57980 4140
rect 58032 4128 58038 4140
rect 59817 4131 59875 4137
rect 59817 4128 59829 4131
rect 58032 4100 59829 4128
rect 58032 4088 58038 4100
rect 59817 4097 59829 4100
rect 59863 4097 59875 4131
rect 59817 4091 59875 4097
rect 23891 4032 24440 4060
rect 26344 4032 27752 4060
rect 27985 4063 28043 4069
rect 23891 4029 23903 4032
rect 23845 4023 23903 4029
rect 21821 3955 21879 3961
rect 22296 3964 23701 3992
rect 25685 3995 25743 4001
rect 15764 3896 18552 3924
rect 20438 3884 20444 3936
rect 20496 3924 20502 3936
rect 20533 3927 20591 3933
rect 20533 3924 20545 3927
rect 20496 3896 20545 3924
rect 20496 3884 20502 3896
rect 20533 3893 20545 3896
rect 20579 3893 20591 3927
rect 21174 3924 21180 3936
rect 21135 3896 21180 3924
rect 20533 3887 20591 3893
rect 21174 3884 21180 3896
rect 21232 3924 21238 3936
rect 22296 3924 22324 3964
rect 25685 3961 25697 3995
rect 25731 3992 25743 3995
rect 25958 3992 25964 4004
rect 25731 3964 25964 3992
rect 25731 3961 25743 3964
rect 25685 3955 25743 3961
rect 25958 3952 25964 3964
rect 26016 3952 26022 4004
rect 26344 3936 26372 4032
rect 27985 4029 27997 4063
rect 28031 4029 28043 4063
rect 27985 4023 28043 4029
rect 59170 4020 59176 4072
rect 59228 4060 59234 4072
rect 61105 4063 61163 4069
rect 61105 4060 61117 4063
rect 59228 4032 61117 4060
rect 59228 4020 59234 4032
rect 61105 4029 61117 4032
rect 61151 4029 61163 4063
rect 61105 4023 61163 4029
rect 27798 3952 27804 4004
rect 27856 3992 27862 4004
rect 29549 3995 29607 4001
rect 29549 3992 29561 3995
rect 27856 3964 29561 3992
rect 27856 3952 27862 3964
rect 29549 3961 29561 3964
rect 29595 3961 29607 3995
rect 29549 3955 29607 3961
rect 57514 3952 57520 4004
rect 57572 3992 57578 4004
rect 58529 3995 58587 4001
rect 58529 3992 58541 3995
rect 57572 3964 58541 3992
rect 57572 3952 57578 3964
rect 58529 3961 58541 3964
rect 58575 3961 58587 3995
rect 58529 3955 58587 3961
rect 58618 3952 58624 4004
rect 58676 3992 58682 4004
rect 60461 3995 60519 4001
rect 60461 3992 60473 3995
rect 58676 3964 60473 3992
rect 58676 3952 58682 3964
rect 60461 3961 60473 3964
rect 60507 3961 60519 3995
rect 60461 3955 60519 3961
rect 21232 3896 22324 3924
rect 21232 3884 21238 3896
rect 22370 3884 22376 3936
rect 22428 3924 22434 3936
rect 22465 3927 22523 3933
rect 22465 3924 22477 3927
rect 22428 3896 22477 3924
rect 22428 3884 22434 3896
rect 22465 3893 22477 3896
rect 22511 3893 22523 3927
rect 26326 3924 26332 3936
rect 26287 3896 26332 3924
rect 22465 3887 22523 3893
rect 26326 3884 26332 3896
rect 26384 3884 26390 3936
rect 32582 3884 32588 3936
rect 32640 3924 32646 3936
rect 32677 3927 32735 3933
rect 32677 3924 32689 3927
rect 32640 3896 32689 3924
rect 32640 3884 32646 3896
rect 32677 3893 32689 3896
rect 32723 3893 32735 3927
rect 32677 3887 32735 3893
rect 56134 3884 56140 3936
rect 56192 3924 56198 3936
rect 56229 3927 56287 3933
rect 56229 3924 56241 3927
rect 56192 3896 56241 3924
rect 56192 3884 56198 3896
rect 56229 3893 56241 3896
rect 56275 3893 56287 3927
rect 56229 3887 56287 3893
rect 56318 3884 56324 3936
rect 56376 3924 56382 3936
rect 56873 3927 56931 3933
rect 56873 3924 56885 3927
rect 56376 3896 56885 3924
rect 56376 3884 56382 3896
rect 56873 3893 56885 3896
rect 56919 3893 56931 3927
rect 56873 3887 56931 3893
rect 56962 3884 56968 3936
rect 57020 3924 57026 3936
rect 57885 3927 57943 3933
rect 57885 3924 57897 3927
rect 57020 3896 57897 3924
rect 57020 3884 57026 3896
rect 57885 3893 57897 3896
rect 57931 3893 57943 3927
rect 57885 3887 57943 3893
rect 58066 3884 58072 3936
rect 58124 3924 58130 3936
rect 59173 3927 59231 3933
rect 59173 3924 59185 3927
rect 58124 3896 59185 3924
rect 58124 3884 58130 3896
rect 59173 3893 59185 3896
rect 59219 3893 59231 3927
rect 59173 3887 59231 3893
rect 1104 3834 68816 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 65654 3834
rect 65706 3782 65718 3834
rect 65770 3782 65782 3834
rect 65834 3782 65846 3834
rect 65898 3782 65910 3834
rect 65962 3782 68816 3834
rect 1104 3760 68816 3782
rect 3878 3680 3884 3732
rect 3936 3720 3942 3732
rect 4157 3723 4215 3729
rect 4157 3720 4169 3723
rect 3936 3692 4169 3720
rect 3936 3680 3942 3692
rect 4157 3689 4169 3692
rect 4203 3689 4215 3723
rect 7466 3720 7472 3732
rect 4157 3683 4215 3689
rect 5460 3692 7472 3720
rect 4893 3655 4951 3661
rect 4893 3621 4905 3655
rect 4939 3621 4951 3655
rect 4893 3615 4951 3621
rect 2314 3544 2320 3596
rect 2372 3584 2378 3596
rect 2409 3587 2467 3593
rect 2409 3584 2421 3587
rect 2372 3556 2421 3584
rect 2372 3544 2378 3556
rect 2409 3553 2421 3556
rect 2455 3553 2467 3587
rect 3786 3584 3792 3596
rect 3747 3556 3792 3584
rect 2409 3547 2467 3553
rect 3786 3544 3792 3556
rect 3844 3544 3850 3596
rect 3050 3516 3056 3528
rect 3011 3488 3056 3516
rect 3050 3476 3056 3488
rect 3108 3476 3114 3528
rect 3878 3516 3884 3528
rect 3160 3488 3884 3516
rect 2317 3451 2375 3457
rect 2317 3417 2329 3451
rect 2363 3448 2375 3451
rect 3160 3448 3188 3488
rect 3878 3476 3884 3488
rect 3936 3476 3942 3528
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3516 4031 3519
rect 4908 3516 4936 3615
rect 5460 3593 5488 3692
rect 7466 3680 7472 3692
rect 7524 3680 7530 3732
rect 7742 3720 7748 3732
rect 7703 3692 7748 3720
rect 7742 3680 7748 3692
rect 7800 3680 7806 3732
rect 8941 3723 8999 3729
rect 8941 3689 8953 3723
rect 8987 3720 8999 3723
rect 9030 3720 9036 3732
rect 8987 3692 9036 3720
rect 8987 3689 8999 3692
rect 8941 3683 8999 3689
rect 9030 3680 9036 3692
rect 9088 3680 9094 3732
rect 9306 3720 9312 3732
rect 9267 3692 9312 3720
rect 9306 3680 9312 3692
rect 9364 3680 9370 3732
rect 9858 3680 9864 3732
rect 9916 3720 9922 3732
rect 9953 3723 10011 3729
rect 9953 3720 9965 3723
rect 9916 3692 9965 3720
rect 9916 3680 9922 3692
rect 9953 3689 9965 3692
rect 9999 3689 10011 3723
rect 10778 3720 10784 3732
rect 10739 3692 10784 3720
rect 9953 3683 10011 3689
rect 10778 3680 10784 3692
rect 10836 3680 10842 3732
rect 10870 3680 10876 3732
rect 10928 3720 10934 3732
rect 10965 3723 11023 3729
rect 10965 3720 10977 3723
rect 10928 3692 10977 3720
rect 10928 3680 10934 3692
rect 10965 3689 10977 3692
rect 11011 3689 11023 3723
rect 11790 3720 11796 3732
rect 11751 3692 11796 3720
rect 10965 3683 11023 3689
rect 11790 3680 11796 3692
rect 11848 3680 11854 3732
rect 11882 3680 11888 3732
rect 11940 3720 11946 3732
rect 12253 3723 12311 3729
rect 11940 3692 11985 3720
rect 11940 3680 11946 3692
rect 12253 3689 12265 3723
rect 12299 3720 12311 3723
rect 12894 3720 12900 3732
rect 12299 3692 12900 3720
rect 12299 3689 12311 3692
rect 12253 3683 12311 3689
rect 12894 3680 12900 3692
rect 12952 3680 12958 3732
rect 14090 3680 14096 3732
rect 14148 3720 14154 3732
rect 14277 3723 14335 3729
rect 14277 3720 14289 3723
rect 14148 3692 14289 3720
rect 14148 3680 14154 3692
rect 14277 3689 14289 3692
rect 14323 3689 14335 3723
rect 14277 3683 14335 3689
rect 14366 3680 14372 3732
rect 14424 3720 14430 3732
rect 15013 3723 15071 3729
rect 15013 3720 15025 3723
rect 14424 3692 15025 3720
rect 14424 3680 14430 3692
rect 15013 3689 15025 3692
rect 15059 3689 15071 3723
rect 15013 3683 15071 3689
rect 15749 3723 15807 3729
rect 15749 3689 15761 3723
rect 15795 3720 15807 3723
rect 15838 3720 15844 3732
rect 15795 3692 15844 3720
rect 15795 3689 15807 3692
rect 15749 3683 15807 3689
rect 15838 3680 15844 3692
rect 15896 3720 15902 3732
rect 21174 3720 21180 3732
rect 15896 3692 21180 3720
rect 15896 3680 15902 3692
rect 21174 3680 21180 3692
rect 21232 3680 21238 3732
rect 23106 3680 23112 3732
rect 23164 3720 23170 3732
rect 23477 3723 23535 3729
rect 23477 3720 23489 3723
rect 23164 3692 23489 3720
rect 23164 3680 23170 3692
rect 23477 3689 23489 3692
rect 23523 3689 23535 3723
rect 23477 3683 23535 3689
rect 27157 3723 27215 3729
rect 27157 3689 27169 3723
rect 27203 3720 27215 3723
rect 27706 3720 27712 3732
rect 27203 3692 27712 3720
rect 27203 3689 27215 3692
rect 27157 3683 27215 3689
rect 27706 3680 27712 3692
rect 27764 3680 27770 3732
rect 31757 3723 31815 3729
rect 31757 3689 31769 3723
rect 31803 3720 31815 3723
rect 32398 3720 32404 3732
rect 31803 3692 32404 3720
rect 31803 3689 31815 3692
rect 31757 3683 31815 3689
rect 32398 3680 32404 3692
rect 32456 3680 32462 3732
rect 57790 3680 57796 3732
rect 57848 3720 57854 3732
rect 58066 3720 58072 3732
rect 57848 3692 58072 3720
rect 57848 3680 57854 3692
rect 58066 3680 58072 3692
rect 58124 3680 58130 3732
rect 7285 3655 7343 3661
rect 7285 3621 7297 3655
rect 7331 3652 7343 3655
rect 7926 3652 7932 3664
rect 7331 3624 7932 3652
rect 7331 3621 7343 3624
rect 7285 3615 7343 3621
rect 7926 3612 7932 3624
rect 7984 3612 7990 3664
rect 8386 3612 8392 3664
rect 8444 3652 8450 3664
rect 13357 3655 13415 3661
rect 8444 3624 11744 3652
rect 8444 3612 8450 3624
rect 5445 3587 5503 3593
rect 5445 3553 5457 3587
rect 5491 3553 5503 3587
rect 5445 3547 5503 3553
rect 8202 3544 8208 3596
rect 8260 3584 8266 3596
rect 8260 3556 9812 3584
rect 8260 3544 8266 3556
rect 4019 3488 4936 3516
rect 4019 3485 4031 3488
rect 3973 3479 4031 3485
rect 6362 3476 6368 3528
rect 6420 3516 6426 3528
rect 6457 3519 6515 3525
rect 6457 3516 6469 3519
rect 6420 3488 6469 3516
rect 6420 3476 6426 3488
rect 6457 3485 6469 3488
rect 6503 3516 6515 3519
rect 6546 3516 6552 3528
rect 6503 3488 6552 3516
rect 6503 3485 6515 3488
rect 6457 3479 6515 3485
rect 6546 3476 6552 3488
rect 6604 3476 6610 3528
rect 7101 3519 7159 3525
rect 7101 3485 7113 3519
rect 7147 3516 7159 3519
rect 7282 3516 7288 3528
rect 7147 3488 7288 3516
rect 7147 3485 7159 3488
rect 7101 3479 7159 3485
rect 7282 3476 7288 3488
rect 7340 3476 7346 3528
rect 7926 3516 7932 3528
rect 7887 3488 7932 3516
rect 7926 3476 7932 3488
rect 7984 3476 7990 3528
rect 8113 3519 8171 3525
rect 8113 3485 8125 3519
rect 8159 3485 8171 3519
rect 9122 3516 9128 3528
rect 9035 3488 9128 3516
rect 8113 3479 8171 3485
rect 2363 3420 3188 3448
rect 3252 3420 6500 3448
rect 2363 3417 2375 3420
rect 2317 3411 2375 3417
rect 1762 3340 1768 3392
rect 1820 3380 1826 3392
rect 1857 3383 1915 3389
rect 1857 3380 1869 3383
rect 1820 3352 1869 3380
rect 1820 3340 1826 3352
rect 1857 3349 1869 3352
rect 1903 3349 1915 3383
rect 2222 3380 2228 3392
rect 2183 3352 2228 3380
rect 1857 3343 1915 3349
rect 2222 3340 2228 3352
rect 2280 3340 2286 3392
rect 3252 3389 3280 3420
rect 6472 3392 6500 3420
rect 7558 3408 7564 3460
rect 7616 3448 7622 3460
rect 8128 3448 8156 3479
rect 7616 3420 8156 3448
rect 7616 3408 7622 3420
rect 3237 3383 3295 3389
rect 3237 3349 3249 3383
rect 3283 3349 3295 3383
rect 5258 3380 5264 3392
rect 5219 3352 5264 3380
rect 3237 3343 3295 3349
rect 5258 3340 5264 3352
rect 5316 3340 5322 3392
rect 5350 3340 5356 3392
rect 5408 3380 5414 3392
rect 5408 3352 5453 3380
rect 5408 3340 5414 3352
rect 6454 3340 6460 3392
rect 6512 3340 6518 3392
rect 6641 3383 6699 3389
rect 6641 3349 6653 3383
rect 6687 3380 6699 3383
rect 7098 3380 7104 3392
rect 6687 3352 7104 3380
rect 6687 3349 6699 3352
rect 6641 3343 6699 3349
rect 7098 3340 7104 3352
rect 7156 3340 7162 3392
rect 7190 3340 7196 3392
rect 7248 3380 7254 3392
rect 9048 3380 9076 3488
rect 9122 3476 9128 3488
rect 9180 3476 9186 3528
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3485 9367 3519
rect 9309 3479 9367 3485
rect 7248 3352 9076 3380
rect 9324 3380 9352 3479
rect 9784 3457 9812 3556
rect 11238 3544 11244 3596
rect 11296 3584 11302 3596
rect 11425 3587 11483 3593
rect 11425 3584 11437 3587
rect 11296 3556 11437 3584
rect 11296 3544 11302 3556
rect 11425 3553 11437 3556
rect 11471 3553 11483 3587
rect 11425 3547 11483 3553
rect 9769 3451 9827 3457
rect 9769 3417 9781 3451
rect 9815 3417 9827 3451
rect 9769 3411 9827 3417
rect 9985 3451 10043 3457
rect 9985 3417 9997 3451
rect 10031 3448 10043 3451
rect 10410 3448 10416 3460
rect 10031 3420 10416 3448
rect 10031 3417 10043 3420
rect 9985 3411 10043 3417
rect 10410 3408 10416 3420
rect 10468 3408 10474 3460
rect 10594 3448 10600 3460
rect 10555 3420 10600 3448
rect 10594 3408 10600 3420
rect 10652 3408 10658 3460
rect 9674 3380 9680 3392
rect 9324 3352 9680 3380
rect 7248 3340 7254 3352
rect 9674 3340 9680 3352
rect 9732 3340 9738 3392
rect 10134 3380 10140 3392
rect 10047 3352 10140 3380
rect 10134 3340 10140 3352
rect 10192 3380 10198 3392
rect 10797 3383 10855 3389
rect 10797 3380 10809 3383
rect 10192 3352 10809 3380
rect 10192 3340 10198 3352
rect 10797 3349 10809 3352
rect 10843 3349 10855 3383
rect 11716 3380 11744 3624
rect 13357 3621 13369 3655
rect 13403 3652 13415 3655
rect 14734 3652 14740 3664
rect 13403 3624 14740 3652
rect 13403 3621 13415 3624
rect 13357 3615 13415 3621
rect 14734 3612 14740 3624
rect 14792 3612 14798 3664
rect 15194 3612 15200 3664
rect 15252 3652 15258 3664
rect 17954 3652 17960 3664
rect 15252 3624 17960 3652
rect 15252 3612 15258 3624
rect 17954 3612 17960 3624
rect 18012 3652 18018 3664
rect 18966 3652 18972 3664
rect 18012 3624 18972 3652
rect 18012 3612 18018 3624
rect 18966 3612 18972 3624
rect 19024 3612 19030 3664
rect 19334 3652 19340 3664
rect 19295 3624 19340 3652
rect 19334 3612 19340 3624
rect 19392 3612 19398 3664
rect 22005 3655 22063 3661
rect 22005 3621 22017 3655
rect 22051 3652 22063 3655
rect 22646 3652 22652 3664
rect 22051 3624 22652 3652
rect 22051 3621 22063 3624
rect 22005 3615 22063 3621
rect 22646 3612 22652 3624
rect 22704 3612 22710 3664
rect 41138 3612 41144 3664
rect 41196 3652 41202 3664
rect 41785 3655 41843 3661
rect 41785 3652 41797 3655
rect 41196 3624 41797 3652
rect 41196 3612 41202 3624
rect 41785 3621 41797 3624
rect 41831 3621 41843 3655
rect 41785 3615 41843 3621
rect 56502 3612 56508 3664
rect 56560 3652 56566 3664
rect 57885 3655 57943 3661
rect 57885 3652 57897 3655
rect 56560 3624 57897 3652
rect 56560 3612 56566 3624
rect 57885 3621 57897 3624
rect 57931 3621 57943 3655
rect 57885 3615 57943 3621
rect 58342 3612 58348 3664
rect 58400 3652 58406 3664
rect 61105 3655 61163 3661
rect 61105 3652 61117 3655
rect 58400 3624 61117 3652
rect 58400 3612 58406 3624
rect 61105 3621 61117 3624
rect 61151 3621 61163 3655
rect 61105 3615 61163 3621
rect 11977 3587 12035 3593
rect 11977 3553 11989 3587
rect 12023 3584 12035 3587
rect 12342 3584 12348 3596
rect 12023 3556 12348 3584
rect 12023 3553 12035 3556
rect 11977 3547 12035 3553
rect 12342 3544 12348 3556
rect 12400 3544 12406 3596
rect 14369 3587 14427 3593
rect 14369 3584 14381 3587
rect 12452 3556 14381 3584
rect 12452 3516 12480 3556
rect 14369 3553 14381 3556
rect 14415 3553 14427 3587
rect 14369 3547 14427 3553
rect 17313 3587 17371 3593
rect 17313 3553 17325 3587
rect 17359 3584 17371 3587
rect 18874 3584 18880 3596
rect 17359 3556 18880 3584
rect 17359 3553 17371 3556
rect 17313 3547 17371 3553
rect 18874 3544 18880 3556
rect 18932 3544 18938 3596
rect 19797 3587 19855 3593
rect 19797 3553 19809 3587
rect 19843 3584 19855 3587
rect 20070 3584 20076 3596
rect 19843 3556 20076 3584
rect 19843 3553 19855 3556
rect 19797 3547 19855 3553
rect 20070 3544 20076 3556
rect 20128 3544 20134 3596
rect 24578 3544 24584 3596
rect 24636 3584 24642 3596
rect 27338 3584 27344 3596
rect 24636 3556 27344 3584
rect 24636 3544 24642 3556
rect 12084 3488 12480 3516
rect 11790 3408 11796 3460
rect 11848 3448 11854 3460
rect 12084 3448 12112 3488
rect 12894 3476 12900 3528
rect 12952 3516 12958 3528
rect 13541 3519 13599 3525
rect 12952 3488 13492 3516
rect 12952 3476 12958 3488
rect 11848 3420 12112 3448
rect 13464 3448 13492 3488
rect 13541 3485 13553 3519
rect 13587 3516 13599 3519
rect 13587 3488 14412 3516
rect 13587 3485 13599 3488
rect 13541 3479 13599 3485
rect 14274 3448 14280 3460
rect 13464 3420 14280 3448
rect 11848 3408 11854 3420
rect 14274 3408 14280 3420
rect 14332 3408 14338 3460
rect 14384 3448 14412 3488
rect 14458 3476 14464 3528
rect 14516 3516 14522 3528
rect 15197 3519 15255 3525
rect 15197 3516 15209 3519
rect 14516 3488 14561 3516
rect 14936 3488 15209 3516
rect 14516 3476 14522 3488
rect 14826 3448 14832 3460
rect 14384 3420 14832 3448
rect 14826 3408 14832 3420
rect 14884 3408 14890 3460
rect 12434 3380 12440 3392
rect 11716 3352 12440 3380
rect 10797 3343 10855 3349
rect 12434 3340 12440 3352
rect 12492 3340 12498 3392
rect 13354 3340 13360 3392
rect 13412 3380 13418 3392
rect 14093 3383 14151 3389
rect 14093 3380 14105 3383
rect 13412 3352 14105 3380
rect 13412 3340 13418 3352
rect 14093 3349 14105 3352
rect 14139 3349 14151 3383
rect 14093 3343 14151 3349
rect 14366 3340 14372 3392
rect 14424 3380 14430 3392
rect 14936 3380 14964 3488
rect 15197 3485 15209 3488
rect 15243 3516 15255 3519
rect 15654 3516 15660 3528
rect 15243 3488 15660 3516
rect 15243 3485 15255 3488
rect 15197 3479 15255 3485
rect 15654 3476 15660 3488
rect 15712 3476 15718 3528
rect 16669 3519 16727 3525
rect 16669 3485 16681 3519
rect 16715 3516 16727 3519
rect 17402 3516 17408 3528
rect 16715 3488 17408 3516
rect 16715 3485 16727 3488
rect 16669 3479 16727 3485
rect 17402 3476 17408 3488
rect 17460 3476 17466 3528
rect 17862 3516 17868 3528
rect 17823 3488 17868 3516
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 18693 3519 18751 3525
rect 18693 3485 18705 3519
rect 18739 3516 18751 3519
rect 19978 3516 19984 3528
rect 18739 3488 19984 3516
rect 18739 3485 18751 3488
rect 18693 3479 18751 3485
rect 19978 3476 19984 3488
rect 20036 3476 20042 3528
rect 20990 3476 20996 3528
rect 21048 3516 21054 3528
rect 21085 3519 21143 3525
rect 21085 3516 21097 3519
rect 21048 3488 21097 3516
rect 21048 3476 21054 3488
rect 21085 3485 21097 3488
rect 21131 3485 21143 3519
rect 21085 3479 21143 3485
rect 22649 3519 22707 3525
rect 22649 3485 22661 3519
rect 22695 3516 22707 3519
rect 23198 3516 23204 3528
rect 22695 3488 23204 3516
rect 22695 3485 22707 3488
rect 22649 3479 22707 3485
rect 23198 3476 23204 3488
rect 23256 3476 23262 3528
rect 24765 3519 24823 3525
rect 24765 3485 24777 3519
rect 24811 3516 24823 3519
rect 24854 3516 24860 3528
rect 24811 3488 24860 3516
rect 24811 3485 24823 3488
rect 24765 3479 24823 3485
rect 24854 3476 24860 3488
rect 24912 3476 24918 3528
rect 25409 3519 25467 3525
rect 25409 3485 25421 3519
rect 25455 3516 25467 3519
rect 25682 3516 25688 3528
rect 25455 3488 25688 3516
rect 25455 3485 25467 3488
rect 25409 3479 25467 3485
rect 25682 3476 25688 3488
rect 25740 3476 25746 3528
rect 26053 3519 26111 3525
rect 26053 3485 26065 3519
rect 26099 3516 26111 3519
rect 26234 3516 26240 3528
rect 26099 3488 26240 3516
rect 26099 3485 26111 3488
rect 26053 3479 26111 3485
rect 26234 3476 26240 3488
rect 26292 3476 26298 3528
rect 26528 3525 26556 3556
rect 27338 3544 27344 3556
rect 27396 3544 27402 3596
rect 33134 3584 33140 3596
rect 33095 3556 33140 3584
rect 33134 3544 33140 3556
rect 33192 3544 33198 3596
rect 55766 3544 55772 3596
rect 55824 3584 55830 3596
rect 56597 3587 56655 3593
rect 56597 3584 56609 3587
rect 55824 3556 56609 3584
rect 55824 3544 55830 3556
rect 56597 3553 56609 3556
rect 56643 3553 56655 3587
rect 56597 3547 56655 3553
rect 56778 3544 56784 3596
rect 56836 3584 56842 3596
rect 58529 3587 58587 3593
rect 58529 3584 58541 3587
rect 56836 3556 58541 3584
rect 56836 3544 56842 3556
rect 58529 3553 58541 3556
rect 58575 3553 58587 3587
rect 58529 3547 58587 3553
rect 58986 3544 58992 3596
rect 59044 3584 59050 3596
rect 61749 3587 61807 3593
rect 61749 3584 61761 3587
rect 59044 3556 61761 3584
rect 59044 3544 59050 3556
rect 61749 3553 61761 3556
rect 61795 3553 61807 3587
rect 61749 3547 61807 3553
rect 26513 3519 26571 3525
rect 26513 3485 26525 3519
rect 26559 3485 26571 3519
rect 26694 3516 26700 3528
rect 26655 3488 26700 3516
rect 26513 3479 26571 3485
rect 26694 3476 26700 3488
rect 26752 3476 26758 3528
rect 26786 3476 26792 3528
rect 26844 3516 26850 3528
rect 26970 3525 26976 3528
rect 26927 3519 26976 3525
rect 26844 3488 26889 3516
rect 26844 3476 26850 3488
rect 26927 3485 26939 3519
rect 26973 3485 26976 3519
rect 26927 3479 26976 3485
rect 26970 3476 26976 3479
rect 27028 3476 27034 3528
rect 27890 3476 27896 3528
rect 27948 3516 27954 3528
rect 27985 3519 28043 3525
rect 27985 3516 27997 3519
rect 27948 3488 27997 3516
rect 27948 3476 27954 3488
rect 27985 3485 27997 3488
rect 28031 3485 28043 3519
rect 27985 3479 28043 3485
rect 28718 3476 28724 3528
rect 28776 3516 28782 3528
rect 28813 3519 28871 3525
rect 28813 3516 28825 3519
rect 28776 3488 28825 3516
rect 28776 3476 28782 3488
rect 28813 3485 28825 3488
rect 28859 3485 28871 3519
rect 28813 3479 28871 3485
rect 29546 3476 29552 3528
rect 29604 3516 29610 3528
rect 29641 3519 29699 3525
rect 29641 3516 29653 3519
rect 29604 3488 29653 3516
rect 29604 3476 29610 3488
rect 29641 3485 29653 3488
rect 29687 3485 29699 3519
rect 30650 3516 30656 3528
rect 30611 3488 30656 3516
rect 29641 3479 29699 3485
rect 30650 3476 30656 3488
rect 30708 3476 30714 3528
rect 31113 3519 31171 3525
rect 31113 3485 31125 3519
rect 31159 3516 31171 3519
rect 31202 3516 31208 3528
rect 31159 3488 31208 3516
rect 31159 3485 31171 3488
rect 31113 3479 31171 3485
rect 31202 3476 31208 3488
rect 31260 3476 31266 3528
rect 32858 3476 32864 3528
rect 32916 3525 32922 3528
rect 32916 3516 32928 3525
rect 32916 3488 32961 3516
rect 32916 3479 32928 3488
rect 32916 3476 32922 3479
rect 39206 3476 39212 3528
rect 39264 3516 39270 3528
rect 39853 3519 39911 3525
rect 39853 3516 39865 3519
rect 39264 3488 39865 3516
rect 39264 3476 39270 3488
rect 39853 3485 39865 3488
rect 39899 3485 39911 3519
rect 39853 3479 39911 3485
rect 40034 3476 40040 3528
rect 40092 3516 40098 3528
rect 40497 3519 40555 3525
rect 40497 3516 40509 3519
rect 40092 3488 40509 3516
rect 40092 3476 40098 3488
rect 40497 3485 40509 3488
rect 40543 3485 40555 3519
rect 40497 3479 40555 3485
rect 40862 3476 40868 3528
rect 40920 3516 40926 3528
rect 41141 3519 41199 3525
rect 41141 3516 41153 3519
rect 40920 3488 41153 3516
rect 40920 3476 40926 3488
rect 41141 3485 41153 3488
rect 41187 3485 41199 3519
rect 41141 3479 41199 3485
rect 42518 3476 42524 3528
rect 42576 3516 42582 3528
rect 42613 3519 42671 3525
rect 42613 3516 42625 3519
rect 42576 3488 42625 3516
rect 42576 3476 42582 3488
rect 42613 3485 42625 3488
rect 42659 3485 42671 3519
rect 42613 3479 42671 3485
rect 43070 3476 43076 3528
rect 43128 3516 43134 3528
rect 43257 3519 43315 3525
rect 43257 3516 43269 3519
rect 43128 3488 43269 3516
rect 43128 3476 43134 3488
rect 43257 3485 43269 3488
rect 43303 3485 43315 3519
rect 43257 3479 43315 3485
rect 45002 3476 45008 3528
rect 45060 3516 45066 3528
rect 45097 3519 45155 3525
rect 45097 3516 45109 3519
rect 45060 3488 45109 3516
rect 45060 3476 45066 3488
rect 45097 3485 45109 3488
rect 45143 3485 45155 3519
rect 45097 3479 45155 3485
rect 45278 3476 45284 3528
rect 45336 3516 45342 3528
rect 45741 3519 45799 3525
rect 45741 3516 45753 3519
rect 45336 3488 45753 3516
rect 45336 3476 45342 3488
rect 45741 3485 45753 3488
rect 45787 3485 45799 3519
rect 45741 3479 45799 3485
rect 46106 3476 46112 3528
rect 46164 3516 46170 3528
rect 46385 3519 46443 3525
rect 46385 3516 46397 3519
rect 46164 3488 46397 3516
rect 46164 3476 46170 3488
rect 46385 3485 46397 3488
rect 46431 3485 46443 3519
rect 46385 3479 46443 3485
rect 46934 3476 46940 3528
rect 46992 3516 46998 3528
rect 47029 3519 47087 3525
rect 47029 3516 47041 3519
rect 46992 3488 47041 3516
rect 46992 3476 46998 3488
rect 47029 3485 47041 3488
rect 47075 3485 47087 3519
rect 47029 3479 47087 3485
rect 47762 3476 47768 3528
rect 47820 3516 47826 3528
rect 47857 3519 47915 3525
rect 47857 3516 47869 3519
rect 47820 3488 47869 3516
rect 47820 3476 47826 3488
rect 47857 3485 47869 3488
rect 47903 3485 47915 3519
rect 47857 3479 47915 3485
rect 48866 3476 48872 3528
rect 48924 3516 48930 3528
rect 48961 3519 49019 3525
rect 48961 3516 48973 3519
rect 48924 3488 48973 3516
rect 48924 3476 48930 3488
rect 48961 3485 48973 3488
rect 49007 3485 49019 3519
rect 48961 3479 49019 3485
rect 50154 3476 50160 3528
rect 50212 3516 50218 3528
rect 50341 3519 50399 3525
rect 50341 3516 50353 3519
rect 50212 3488 50353 3516
rect 50212 3476 50218 3488
rect 50341 3485 50353 3488
rect 50387 3485 50399 3519
rect 50341 3479 50399 3485
rect 50798 3476 50804 3528
rect 50856 3516 50862 3528
rect 50985 3519 51043 3525
rect 50985 3516 50997 3519
rect 50856 3488 50997 3516
rect 50856 3476 50862 3488
rect 50985 3485 50997 3488
rect 51031 3485 51043 3519
rect 50985 3479 51043 3485
rect 51350 3476 51356 3528
rect 51408 3516 51414 3528
rect 51629 3519 51687 3525
rect 51629 3516 51641 3519
rect 51408 3488 51641 3516
rect 51408 3476 51414 3488
rect 51629 3485 51641 3488
rect 51675 3485 51687 3519
rect 51629 3479 51687 3485
rect 52730 3476 52736 3528
rect 52788 3516 52794 3528
rect 52825 3519 52883 3525
rect 52825 3516 52837 3519
rect 52788 3488 52837 3516
rect 52788 3476 52794 3488
rect 52825 3485 52837 3488
rect 52871 3485 52883 3519
rect 52825 3479 52883 3485
rect 53006 3476 53012 3528
rect 53064 3516 53070 3528
rect 53469 3519 53527 3525
rect 53469 3516 53481 3519
rect 53064 3488 53481 3516
rect 53064 3476 53070 3488
rect 53469 3485 53481 3488
rect 53515 3485 53527 3519
rect 53469 3479 53527 3485
rect 54662 3476 54668 3528
rect 54720 3516 54726 3528
rect 55309 3519 55367 3525
rect 55309 3516 55321 3519
rect 54720 3488 55321 3516
rect 54720 3476 54726 3488
rect 55309 3485 55321 3488
rect 55355 3485 55367 3519
rect 55309 3479 55367 3485
rect 55490 3476 55496 3528
rect 55548 3516 55554 3528
rect 55953 3519 56011 3525
rect 55953 3516 55965 3519
rect 55548 3488 55965 3516
rect 55548 3476 55554 3488
rect 55953 3485 55965 3488
rect 55999 3485 56011 3519
rect 55953 3479 56011 3485
rect 56226 3476 56232 3528
rect 56284 3516 56290 3528
rect 57241 3519 57299 3525
rect 57241 3516 57253 3519
rect 56284 3488 57253 3516
rect 56284 3476 56290 3488
rect 57241 3485 57253 3488
rect 57287 3485 57299 3519
rect 57241 3479 57299 3485
rect 57330 3476 57336 3528
rect 57388 3516 57394 3528
rect 59173 3519 59231 3525
rect 59173 3516 59185 3519
rect 57388 3488 59185 3516
rect 57388 3476 57394 3488
rect 59173 3485 59185 3488
rect 59219 3485 59231 3519
rect 60458 3516 60464 3528
rect 60419 3488 60464 3516
rect 59173 3479 59231 3485
rect 60458 3476 60464 3488
rect 60516 3476 60522 3528
rect 68094 3516 68100 3528
rect 68055 3488 68100 3516
rect 68094 3476 68100 3488
rect 68152 3476 68158 3528
rect 15102 3408 15108 3460
rect 15160 3448 15166 3460
rect 15841 3451 15899 3457
rect 15841 3448 15853 3451
rect 15160 3420 15853 3448
rect 15160 3408 15166 3420
rect 15841 3417 15853 3420
rect 15887 3448 15899 3451
rect 18414 3448 18420 3460
rect 15887 3420 18420 3448
rect 15887 3417 15899 3420
rect 15841 3411 15899 3417
rect 18414 3408 18420 3420
rect 18472 3408 18478 3460
rect 19337 3451 19395 3457
rect 19337 3417 19349 3451
rect 19383 3417 19395 3451
rect 19337 3411 19395 3417
rect 16482 3380 16488 3392
rect 14424 3352 14964 3380
rect 16443 3352 16488 3380
rect 14424 3340 14430 3352
rect 16482 3340 16488 3352
rect 16540 3340 16546 3392
rect 18049 3383 18107 3389
rect 18049 3349 18061 3383
rect 18095 3380 18107 3383
rect 19352 3380 19380 3411
rect 19426 3408 19432 3460
rect 19484 3448 19490 3460
rect 19889 3451 19947 3457
rect 19889 3448 19901 3451
rect 19484 3420 19901 3448
rect 19484 3408 19490 3420
rect 19889 3417 19901 3420
rect 19935 3417 19947 3451
rect 20070 3448 20076 3460
rect 20031 3420 20076 3448
rect 19889 3411 19947 3417
rect 20070 3408 20076 3420
rect 20128 3408 20134 3460
rect 23014 3408 23020 3460
rect 23072 3448 23078 3460
rect 23109 3451 23167 3457
rect 23109 3448 23121 3451
rect 23072 3420 23121 3448
rect 23072 3408 23078 3420
rect 23109 3417 23121 3420
rect 23155 3417 23167 3451
rect 23109 3411 23167 3417
rect 23293 3451 23351 3457
rect 23293 3417 23305 3451
rect 23339 3448 23351 3451
rect 25958 3448 25964 3460
rect 23339 3420 25964 3448
rect 23339 3417 23351 3420
rect 23293 3411 23351 3417
rect 25958 3408 25964 3420
rect 26016 3408 26022 3460
rect 18095 3352 19380 3380
rect 18095 3349 18107 3352
rect 18049 3343 18107 3349
rect 20162 3340 20168 3392
rect 20220 3380 20226 3392
rect 20533 3383 20591 3389
rect 20533 3380 20545 3383
rect 20220 3352 20545 3380
rect 20220 3340 20226 3352
rect 20533 3349 20545 3352
rect 20579 3349 20591 3383
rect 20533 3343 20591 3349
rect 1104 3290 68816 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 68816 3290
rect 1104 3216 68816 3238
rect 1394 3136 1400 3188
rect 1452 3176 1458 3188
rect 1581 3179 1639 3185
rect 1581 3176 1593 3179
rect 1452 3148 1593 3176
rect 1452 3136 1458 3148
rect 1581 3145 1593 3148
rect 1627 3145 1639 3179
rect 3970 3176 3976 3188
rect 3931 3148 3976 3176
rect 1581 3139 1639 3145
rect 3970 3136 3976 3148
rect 4028 3136 4034 3188
rect 4614 3176 4620 3188
rect 4448 3148 4620 3176
rect 2958 3108 2964 3120
rect 2608 3080 2964 3108
rect 1762 3040 1768 3052
rect 1723 3012 1768 3040
rect 1762 3000 1768 3012
rect 1820 3000 1826 3052
rect 1946 3040 1952 3052
rect 1907 3012 1952 3040
rect 1946 3000 1952 3012
rect 2004 3000 2010 3052
rect 2608 3049 2636 3080
rect 2958 3068 2964 3080
rect 3016 3108 3022 3120
rect 3016 3080 3832 3108
rect 3016 3068 3022 3080
rect 2866 3049 2872 3052
rect 2593 3043 2651 3049
rect 2593 3009 2605 3043
rect 2639 3009 2651 3043
rect 2593 3003 2651 3009
rect 2860 3003 2872 3049
rect 2924 3040 2930 3052
rect 3804 3040 3832 3080
rect 4448 3049 4476 3148
rect 4614 3136 4620 3148
rect 4672 3136 4678 3188
rect 5350 3136 5356 3188
rect 5408 3176 5414 3188
rect 5813 3179 5871 3185
rect 5813 3176 5825 3179
rect 5408 3148 5825 3176
rect 5408 3136 5414 3148
rect 5813 3145 5825 3148
rect 5859 3176 5871 3179
rect 7006 3176 7012 3188
rect 5859 3148 7012 3176
rect 5859 3145 5871 3148
rect 5813 3139 5871 3145
rect 7006 3136 7012 3148
rect 7064 3136 7070 3188
rect 7745 3179 7803 3185
rect 7745 3145 7757 3179
rect 7791 3176 7803 3179
rect 8018 3176 8024 3188
rect 7791 3148 8024 3176
rect 7791 3145 7803 3148
rect 7745 3139 7803 3145
rect 8018 3136 8024 3148
rect 8076 3136 8082 3188
rect 8110 3136 8116 3188
rect 8168 3176 8174 3188
rect 8938 3176 8944 3188
rect 8168 3148 8944 3176
rect 8168 3136 8174 3148
rect 8938 3136 8944 3148
rect 8996 3176 9002 3188
rect 10134 3176 10140 3188
rect 8996 3148 10140 3176
rect 8996 3136 9002 3148
rect 10134 3136 10140 3148
rect 10192 3136 10198 3188
rect 11606 3136 11612 3188
rect 11664 3176 11670 3188
rect 11882 3176 11888 3188
rect 11664 3148 11888 3176
rect 11664 3136 11670 3148
rect 11882 3136 11888 3148
rect 11940 3136 11946 3188
rect 11974 3136 11980 3188
rect 12032 3176 12038 3188
rect 12250 3176 12256 3188
rect 12032 3148 12256 3176
rect 12032 3136 12038 3148
rect 12250 3136 12256 3148
rect 12308 3136 12314 3188
rect 12529 3179 12587 3185
rect 12529 3145 12541 3179
rect 12575 3176 12587 3179
rect 12986 3176 12992 3188
rect 12575 3148 12992 3176
rect 12575 3145 12587 3148
rect 12529 3139 12587 3145
rect 12986 3136 12992 3148
rect 13044 3136 13050 3188
rect 13354 3136 13360 3188
rect 13412 3176 13418 3188
rect 16482 3176 16488 3188
rect 13412 3148 16488 3176
rect 13412 3136 13418 3148
rect 16482 3136 16488 3148
rect 16540 3136 16546 3188
rect 18693 3179 18751 3185
rect 18693 3145 18705 3179
rect 18739 3176 18751 3179
rect 19334 3176 19340 3188
rect 18739 3148 19340 3176
rect 18739 3145 18751 3148
rect 18693 3139 18751 3145
rect 19334 3136 19340 3148
rect 19392 3136 19398 3188
rect 19426 3136 19432 3188
rect 19484 3176 19490 3188
rect 20254 3176 20260 3188
rect 19484 3148 20260 3176
rect 19484 3136 19490 3148
rect 20254 3136 20260 3148
rect 20312 3136 20318 3188
rect 21913 3179 21971 3185
rect 21913 3145 21925 3179
rect 21959 3176 21971 3179
rect 22002 3176 22008 3188
rect 21959 3148 22008 3176
rect 21959 3145 21971 3148
rect 21913 3139 21971 3145
rect 22002 3136 22008 3148
rect 22060 3136 22066 3188
rect 26418 3136 26424 3188
rect 26476 3176 26482 3188
rect 26970 3176 26976 3188
rect 26476 3148 26976 3176
rect 26476 3136 26482 3148
rect 26970 3136 26976 3148
rect 27028 3136 27034 3188
rect 55950 3136 55956 3188
rect 56008 3176 56014 3188
rect 58066 3176 58072 3188
rect 56008 3148 58072 3176
rect 56008 3136 56014 3148
rect 58066 3136 58072 3148
rect 58124 3136 58130 3188
rect 4706 3117 4712 3120
rect 4700 3108 4712 3117
rect 4667 3080 4712 3108
rect 4700 3071 4712 3080
rect 4706 3068 4712 3071
rect 4764 3068 4770 3120
rect 9950 3108 9956 3120
rect 6380 3080 9956 3108
rect 6380 3049 6408 3080
rect 4433 3043 4491 3049
rect 4433 3040 4445 3043
rect 2924 3012 2960 3040
rect 3804 3012 4445 3040
rect 2866 3000 2872 3003
rect 2924 3000 2930 3012
rect 4433 3009 4445 3012
rect 4479 3009 4491 3043
rect 4433 3003 4491 3009
rect 6365 3043 6423 3049
rect 6365 3009 6377 3043
rect 6411 3009 6423 3043
rect 6365 3003 6423 3009
rect 6454 3000 6460 3052
rect 6512 3040 6518 3052
rect 6621 3043 6679 3049
rect 6621 3040 6633 3043
rect 6512 3012 6633 3040
rect 6512 3000 6518 3012
rect 6621 3009 6633 3012
rect 6667 3009 6679 3043
rect 6621 3003 6679 3009
rect 7098 3000 7104 3052
rect 7156 3040 7162 3052
rect 7156 3012 8892 3040
rect 7156 3000 7162 3012
rect 8481 2907 8539 2913
rect 8481 2904 8493 2907
rect 7300 2876 8493 2904
rect 6362 2796 6368 2848
rect 6420 2836 6426 2848
rect 7300 2836 7328 2876
rect 8481 2873 8493 2876
rect 8527 2873 8539 2907
rect 8481 2867 8539 2873
rect 6420 2808 7328 2836
rect 8864 2836 8892 3012
rect 9214 3000 9220 3052
rect 9272 3040 9278 3052
rect 9876 3049 9904 3080
rect 9950 3068 9956 3080
rect 10008 3068 10014 3120
rect 10042 3068 10048 3120
rect 10100 3108 10106 3120
rect 10505 3111 10563 3117
rect 10505 3108 10517 3111
rect 10100 3080 10517 3108
rect 10100 3068 10106 3080
rect 10505 3077 10517 3080
rect 10551 3108 10563 3111
rect 12894 3108 12900 3120
rect 10551 3080 12900 3108
rect 10551 3077 10563 3080
rect 10505 3071 10563 3077
rect 12894 3068 12900 3080
rect 12952 3068 12958 3120
rect 13078 3108 13084 3120
rect 13039 3080 13084 3108
rect 13078 3068 13084 3080
rect 13136 3068 13142 3120
rect 13814 3068 13820 3120
rect 13872 3108 13878 3120
rect 15102 3108 15108 3120
rect 13872 3080 15108 3108
rect 13872 3068 13878 3080
rect 15102 3068 15108 3080
rect 15160 3068 15166 3120
rect 17862 3068 17868 3120
rect 17920 3108 17926 3120
rect 20622 3108 20628 3120
rect 17920 3080 20628 3108
rect 17920 3068 17926 3080
rect 20622 3068 20628 3080
rect 20680 3068 20686 3120
rect 57698 3068 57704 3120
rect 57756 3108 57762 3120
rect 60458 3108 60464 3120
rect 57756 3080 60464 3108
rect 57756 3068 57762 3080
rect 60458 3068 60464 3080
rect 60516 3068 60522 3120
rect 9594 3043 9652 3049
rect 9594 3040 9606 3043
rect 9272 3012 9606 3040
rect 9272 3000 9278 3012
rect 9594 3009 9606 3012
rect 9640 3009 9652 3043
rect 9594 3003 9652 3009
rect 9861 3043 9919 3049
rect 9861 3009 9873 3043
rect 9907 3009 9919 3043
rect 9861 3003 9919 3009
rect 10873 3043 10931 3049
rect 10873 3009 10885 3043
rect 10919 3040 10931 3043
rect 11606 3040 11612 3052
rect 10919 3012 11612 3040
rect 10919 3009 10931 3012
rect 10873 3003 10931 3009
rect 11606 3000 11612 3012
rect 11664 3000 11670 3052
rect 11790 3000 11796 3052
rect 11848 3040 11854 3052
rect 11885 3043 11943 3049
rect 11885 3040 11897 3043
rect 11848 3012 11897 3040
rect 11848 3000 11854 3012
rect 11885 3009 11897 3012
rect 11931 3009 11943 3043
rect 11885 3003 11943 3009
rect 11977 3043 12035 3049
rect 11977 3009 11989 3043
rect 12023 3040 12035 3043
rect 12158 3040 12164 3052
rect 12023 3012 12164 3040
rect 12023 3009 12035 3012
rect 11977 3003 12035 3009
rect 11238 2932 11244 2984
rect 11296 2972 11302 2984
rect 11992 2972 12020 3003
rect 12158 3000 12164 3012
rect 12216 3000 12222 3052
rect 12342 3040 12348 3052
rect 12303 3012 12348 3040
rect 12342 3000 12348 3012
rect 12400 3000 12406 3052
rect 13096 3040 13124 3068
rect 13096 3012 13492 3040
rect 11296 2944 12020 2972
rect 11296 2932 11302 2944
rect 12434 2932 12440 2984
rect 12492 2972 12498 2984
rect 13357 2975 13415 2981
rect 13357 2972 13369 2975
rect 12492 2944 13369 2972
rect 12492 2932 12498 2944
rect 13357 2941 13369 2944
rect 13403 2941 13415 2975
rect 13464 2972 13492 3012
rect 13538 3000 13544 3052
rect 13596 3040 13602 3052
rect 13596 3012 13641 3040
rect 13596 3000 13602 3012
rect 13906 3000 13912 3052
rect 13964 3040 13970 3052
rect 14461 3043 14519 3049
rect 14461 3040 14473 3043
rect 13964 3012 14473 3040
rect 13964 3000 13970 3012
rect 14461 3009 14473 3012
rect 14507 3009 14519 3043
rect 14461 3003 14519 3009
rect 14550 3000 14556 3052
rect 14608 3040 14614 3052
rect 15473 3043 15531 3049
rect 15473 3040 15485 3043
rect 14608 3012 15485 3040
rect 14608 3000 14614 3012
rect 15473 3009 15485 3012
rect 15519 3009 15531 3043
rect 15473 3003 15531 3009
rect 16850 3000 16856 3052
rect 16908 3040 16914 3052
rect 16945 3043 17003 3049
rect 16945 3040 16957 3043
rect 16908 3012 16957 3040
rect 16908 3000 16914 3012
rect 16945 3009 16957 3012
rect 16991 3009 17003 3043
rect 17586 3040 17592 3052
rect 17547 3012 17592 3040
rect 16945 3003 17003 3009
rect 17586 3000 17592 3012
rect 17644 3000 17650 3052
rect 18509 3043 18567 3049
rect 18509 3009 18521 3043
rect 18555 3040 18567 3043
rect 20070 3040 20076 3052
rect 18555 3012 20076 3040
rect 18555 3009 18567 3012
rect 18509 3003 18567 3009
rect 20070 3000 20076 3012
rect 20128 3000 20134 3052
rect 58158 3000 58164 3052
rect 58216 3040 58222 3052
rect 61105 3043 61163 3049
rect 61105 3040 61117 3043
rect 58216 3012 61117 3040
rect 58216 3000 58222 3012
rect 61105 3009 61117 3012
rect 61151 3009 61163 3043
rect 61105 3003 61163 3009
rect 14185 2975 14243 2981
rect 14185 2972 14197 2975
rect 13464 2944 14197 2972
rect 13357 2935 13415 2941
rect 14185 2941 14197 2944
rect 14231 2941 14243 2975
rect 14185 2935 14243 2941
rect 14274 2932 14280 2984
rect 14332 2972 14338 2984
rect 18690 2972 18696 2984
rect 14332 2944 18696 2972
rect 14332 2932 14338 2944
rect 18690 2932 18696 2944
rect 18748 2932 18754 2984
rect 19981 2975 20039 2981
rect 19981 2941 19993 2975
rect 20027 2972 20039 2975
rect 20714 2972 20720 2984
rect 20027 2944 20720 2972
rect 20027 2941 20039 2944
rect 19981 2935 20039 2941
rect 20714 2932 20720 2944
rect 20772 2932 20778 2984
rect 21269 2975 21327 2981
rect 21269 2941 21281 2975
rect 21315 2972 21327 2975
rect 21818 2972 21824 2984
rect 21315 2944 21824 2972
rect 21315 2941 21327 2944
rect 21269 2935 21327 2941
rect 21818 2932 21824 2944
rect 21876 2932 21882 2984
rect 24489 2975 24547 2981
rect 24489 2941 24501 2975
rect 24535 2972 24547 2975
rect 25130 2972 25136 2984
rect 24535 2944 25136 2972
rect 24535 2941 24547 2944
rect 24489 2935 24547 2941
rect 25130 2932 25136 2944
rect 25188 2932 25194 2984
rect 28353 2975 28411 2981
rect 28353 2941 28365 2975
rect 28399 2972 28411 2975
rect 28994 2972 29000 2984
rect 28399 2944 29000 2972
rect 28399 2941 28411 2944
rect 28353 2935 28411 2941
rect 28994 2932 29000 2944
rect 29052 2932 29058 2984
rect 30285 2975 30343 2981
rect 30285 2941 30297 2975
rect 30331 2972 30343 2975
rect 30926 2972 30932 2984
rect 30331 2944 30932 2972
rect 30331 2941 30343 2944
rect 30285 2935 30343 2941
rect 30926 2932 30932 2944
rect 30984 2932 30990 2984
rect 37274 2932 37280 2984
rect 37332 2972 37338 2984
rect 37921 2975 37979 2981
rect 37921 2972 37933 2975
rect 37332 2944 37933 2972
rect 37332 2932 37338 2944
rect 37921 2941 37933 2944
rect 37967 2941 37979 2975
rect 37921 2935 37979 2941
rect 44726 2932 44732 2984
rect 44784 2972 44790 2984
rect 45649 2975 45707 2981
rect 45649 2972 45661 2975
rect 44784 2944 45661 2972
rect 44784 2932 44790 2944
rect 45649 2941 45661 2944
rect 45695 2941 45707 2975
rect 45649 2935 45707 2941
rect 48590 2932 48596 2984
rect 48648 2972 48654 2984
rect 49513 2975 49571 2981
rect 49513 2972 49525 2975
rect 48648 2944 49525 2972
rect 48648 2932 48654 2944
rect 49513 2941 49525 2944
rect 49559 2941 49571 2975
rect 49513 2935 49571 2941
rect 52454 2932 52460 2984
rect 52512 2972 52518 2984
rect 53377 2975 53435 2981
rect 53377 2972 53389 2975
rect 52512 2944 53389 2972
rect 52512 2932 52518 2944
rect 53377 2941 53389 2944
rect 53423 2941 53435 2975
rect 53377 2935 53435 2941
rect 53558 2932 53564 2984
rect 53616 2972 53622 2984
rect 55214 2972 55220 2984
rect 53616 2944 55220 2972
rect 53616 2932 53622 2944
rect 55214 2932 55220 2944
rect 55272 2932 55278 2984
rect 56686 2932 56692 2984
rect 56744 2972 56750 2984
rect 56744 2944 58204 2972
rect 56744 2932 56750 2944
rect 11790 2904 11796 2916
rect 11624 2876 11796 2904
rect 11624 2836 11652 2876
rect 11790 2864 11796 2876
rect 11848 2864 11854 2916
rect 11882 2864 11888 2916
rect 11940 2904 11946 2916
rect 11940 2876 13216 2904
rect 11940 2864 11946 2876
rect 8864 2808 11652 2836
rect 6420 2796 6426 2808
rect 11698 2796 11704 2848
rect 11756 2836 11762 2848
rect 13188 2845 13216 2876
rect 13262 2864 13268 2916
rect 13320 2864 13326 2916
rect 13630 2864 13636 2916
rect 13688 2904 13694 2916
rect 16761 2907 16819 2913
rect 16761 2904 16773 2907
rect 13688 2876 16773 2904
rect 13688 2864 13694 2876
rect 16761 2873 16773 2876
rect 16807 2873 16819 2907
rect 16761 2867 16819 2873
rect 19337 2907 19395 2913
rect 19337 2873 19349 2907
rect 19383 2904 19395 2907
rect 20254 2904 20260 2916
rect 19383 2876 20260 2904
rect 19383 2873 19395 2876
rect 19337 2867 19395 2873
rect 20254 2864 20260 2876
rect 20312 2864 20318 2916
rect 22002 2904 22008 2916
rect 20364 2876 22008 2904
rect 12345 2839 12403 2845
rect 12345 2836 12357 2839
rect 11756 2808 12357 2836
rect 11756 2796 11762 2808
rect 12345 2805 12357 2808
rect 12391 2805 12403 2839
rect 12345 2799 12403 2805
rect 13173 2839 13231 2845
rect 13173 2805 13185 2839
rect 13219 2805 13231 2839
rect 13280 2836 13308 2864
rect 13725 2839 13783 2845
rect 13725 2836 13737 2839
rect 13280 2808 13737 2836
rect 13173 2799 13231 2805
rect 13725 2805 13737 2808
rect 13771 2805 13783 2839
rect 13725 2799 13783 2805
rect 14182 2796 14188 2848
rect 14240 2836 14246 2848
rect 15657 2839 15715 2845
rect 15657 2836 15669 2839
rect 14240 2808 15669 2836
rect 14240 2796 14246 2808
rect 15657 2805 15669 2808
rect 15703 2805 15715 2839
rect 15657 2799 15715 2805
rect 17497 2839 17555 2845
rect 17497 2805 17509 2839
rect 17543 2836 17555 2839
rect 17770 2836 17776 2848
rect 17543 2808 17776 2836
rect 17543 2805 17555 2808
rect 17497 2799 17555 2805
rect 17770 2796 17776 2808
rect 17828 2796 17834 2848
rect 20162 2796 20168 2848
rect 20220 2836 20226 2848
rect 20364 2836 20392 2876
rect 22002 2864 22008 2876
rect 22060 2864 22066 2916
rect 22557 2907 22615 2913
rect 22557 2873 22569 2907
rect 22603 2904 22615 2907
rect 23474 2904 23480 2916
rect 22603 2876 23480 2904
rect 22603 2873 22615 2876
rect 22557 2867 22615 2873
rect 23474 2864 23480 2876
rect 23532 2864 23538 2916
rect 25958 2904 25964 2916
rect 25148 2876 25964 2904
rect 20220 2808 20392 2836
rect 20625 2839 20683 2845
rect 20220 2796 20226 2808
rect 20625 2805 20637 2839
rect 20671 2836 20683 2839
rect 21266 2836 21272 2848
rect 20671 2808 21272 2836
rect 20671 2805 20683 2808
rect 20625 2799 20683 2805
rect 21266 2796 21272 2808
rect 21324 2796 21330 2848
rect 23201 2839 23259 2845
rect 23201 2805 23213 2839
rect 23247 2836 23259 2839
rect 23750 2836 23756 2848
rect 23247 2808 23756 2836
rect 23247 2805 23259 2808
rect 23201 2799 23259 2805
rect 23750 2796 23756 2808
rect 23808 2796 23814 2848
rect 23845 2839 23903 2845
rect 23845 2805 23857 2839
rect 23891 2836 23903 2839
rect 24302 2836 24308 2848
rect 23891 2808 24308 2836
rect 23891 2805 23903 2808
rect 23845 2799 23903 2805
rect 24302 2796 24308 2808
rect 24360 2796 24366 2848
rect 25148 2845 25176 2876
rect 25958 2864 25964 2876
rect 26016 2864 26022 2916
rect 26421 2907 26479 2913
rect 26421 2873 26433 2907
rect 26467 2904 26479 2907
rect 27062 2904 27068 2916
rect 26467 2876 27068 2904
rect 26467 2873 26479 2876
rect 26421 2867 26479 2873
rect 27062 2864 27068 2876
rect 27120 2864 27126 2916
rect 38378 2864 38384 2916
rect 38436 2904 38442 2916
rect 39209 2907 39267 2913
rect 39209 2904 39221 2907
rect 38436 2876 39221 2904
rect 38436 2864 38442 2876
rect 39209 2873 39221 2876
rect 39255 2873 39267 2907
rect 39209 2867 39267 2873
rect 39758 2864 39764 2916
rect 39816 2904 39822 2916
rect 40497 2907 40555 2913
rect 40497 2904 40509 2907
rect 39816 2876 40509 2904
rect 39816 2864 39822 2876
rect 40497 2873 40509 2876
rect 40543 2873 40555 2907
rect 40497 2867 40555 2873
rect 42242 2864 42248 2916
rect 42300 2904 42306 2916
rect 43073 2907 43131 2913
rect 43073 2904 43085 2907
rect 42300 2876 43085 2904
rect 42300 2864 42306 2876
rect 43073 2873 43085 2876
rect 43119 2873 43131 2907
rect 43073 2867 43131 2873
rect 43622 2864 43628 2916
rect 43680 2904 43686 2916
rect 44361 2907 44419 2913
rect 44361 2904 44373 2907
rect 43680 2876 44373 2904
rect 43680 2864 43686 2876
rect 44361 2873 44373 2876
rect 44407 2873 44419 2907
rect 44361 2867 44419 2873
rect 47486 2864 47492 2916
rect 47544 2904 47550 2916
rect 48225 2907 48283 2913
rect 48225 2904 48237 2907
rect 47544 2876 48237 2904
rect 47544 2864 47550 2876
rect 48225 2873 48237 2876
rect 48271 2873 48283 2907
rect 48225 2867 48283 2873
rect 49418 2864 49424 2916
rect 49476 2904 49482 2916
rect 50157 2907 50215 2913
rect 50157 2904 50169 2907
rect 49476 2876 50169 2904
rect 49476 2864 49482 2876
rect 50157 2873 50169 2876
rect 50203 2873 50215 2907
rect 50157 2867 50215 2873
rect 50614 2864 50620 2916
rect 50672 2904 50678 2916
rect 51445 2907 51503 2913
rect 51445 2904 51457 2907
rect 50672 2876 51457 2904
rect 50672 2864 50678 2876
rect 51445 2873 51457 2876
rect 51491 2873 51503 2907
rect 51445 2867 51503 2873
rect 53282 2864 53288 2916
rect 53340 2904 53346 2916
rect 54021 2907 54079 2913
rect 54021 2904 54033 2907
rect 53340 2876 54033 2904
rect 53340 2864 53346 2876
rect 54021 2873 54033 2876
rect 54067 2873 54079 2907
rect 54021 2867 54079 2873
rect 54386 2864 54392 2916
rect 54444 2904 54450 2916
rect 55309 2907 55367 2913
rect 55309 2904 55321 2907
rect 54444 2876 55321 2904
rect 54444 2864 54450 2876
rect 55309 2873 55321 2876
rect 55355 2873 55367 2907
rect 55309 2867 55367 2873
rect 55674 2864 55680 2916
rect 55732 2904 55738 2916
rect 56597 2907 56655 2913
rect 56597 2904 56609 2907
rect 55732 2876 56609 2904
rect 55732 2864 55738 2876
rect 56597 2873 56609 2876
rect 56643 2873 56655 2907
rect 56597 2867 56655 2873
rect 57054 2864 57060 2916
rect 57112 2904 57118 2916
rect 58176 2904 58204 2944
rect 58434 2932 58440 2984
rect 58492 2972 58498 2984
rect 61749 2975 61807 2981
rect 61749 2972 61761 2975
rect 58492 2944 61761 2972
rect 58492 2932 58498 2944
rect 61749 2941 61761 2944
rect 61795 2941 61807 2975
rect 61749 2935 61807 2941
rect 58529 2907 58587 2913
rect 58529 2904 58541 2907
rect 57112 2876 58020 2904
rect 58176 2876 58541 2904
rect 57112 2864 57118 2876
rect 25133 2839 25191 2845
rect 25133 2805 25145 2839
rect 25179 2805 25191 2839
rect 25133 2799 25191 2805
rect 25777 2839 25835 2845
rect 25777 2805 25789 2839
rect 25823 2836 25835 2839
rect 26786 2836 26792 2848
rect 25823 2808 26792 2836
rect 25823 2805 25835 2808
rect 25777 2799 25835 2805
rect 26786 2796 26792 2808
rect 26844 2796 26850 2848
rect 27709 2839 27767 2845
rect 27709 2805 27721 2839
rect 27755 2836 27767 2839
rect 28166 2836 28172 2848
rect 27755 2808 28172 2836
rect 27755 2805 27767 2808
rect 27709 2799 27767 2805
rect 28166 2796 28172 2808
rect 28224 2796 28230 2848
rect 28997 2839 29055 2845
rect 28997 2805 29009 2839
rect 29043 2836 29055 2839
rect 29270 2836 29276 2848
rect 29043 2808 29276 2836
rect 29043 2805 29055 2808
rect 28997 2799 29055 2805
rect 29270 2796 29276 2808
rect 29328 2796 29334 2848
rect 29641 2839 29699 2845
rect 29641 2805 29653 2839
rect 29687 2836 29699 2839
rect 30098 2836 30104 2848
rect 29687 2808 30104 2836
rect 29687 2805 29699 2808
rect 29641 2799 29699 2805
rect 30098 2796 30104 2808
rect 30156 2796 30162 2848
rect 30929 2839 30987 2845
rect 30929 2805 30941 2839
rect 30975 2836 30987 2839
rect 31478 2836 31484 2848
rect 30975 2808 31484 2836
rect 30975 2805 30987 2808
rect 30929 2799 30987 2805
rect 31478 2796 31484 2808
rect 31536 2796 31542 2848
rect 31573 2839 31631 2845
rect 31573 2805 31585 2839
rect 31619 2836 31631 2839
rect 32030 2836 32036 2848
rect 31619 2808 32036 2836
rect 31619 2805 31631 2808
rect 31573 2799 31631 2805
rect 32030 2796 32036 2808
rect 32088 2796 32094 2848
rect 32861 2839 32919 2845
rect 32861 2805 32873 2839
rect 32907 2836 32919 2839
rect 33134 2836 33140 2848
rect 32907 2808 33140 2836
rect 32907 2805 32919 2808
rect 32861 2799 32919 2805
rect 33134 2796 33140 2808
rect 33192 2796 33198 2848
rect 33505 2839 33563 2845
rect 33505 2805 33517 2839
rect 33551 2836 33563 2839
rect 33686 2836 33692 2848
rect 33551 2808 33692 2836
rect 33551 2805 33563 2808
rect 33505 2799 33563 2805
rect 33686 2796 33692 2808
rect 33744 2796 33750 2848
rect 34149 2839 34207 2845
rect 34149 2805 34161 2839
rect 34195 2836 34207 2839
rect 34238 2836 34244 2848
rect 34195 2808 34244 2836
rect 34195 2805 34207 2808
rect 34149 2799 34207 2805
rect 34238 2796 34244 2808
rect 34296 2796 34302 2848
rect 34514 2796 34520 2848
rect 34572 2836 34578 2848
rect 34609 2839 34667 2845
rect 34609 2836 34621 2839
rect 34572 2808 34621 2836
rect 34572 2796 34578 2808
rect 34609 2805 34621 2808
rect 34655 2805 34667 2839
rect 34609 2799 34667 2805
rect 35342 2796 35348 2848
rect 35400 2836 35406 2848
rect 35437 2839 35495 2845
rect 35437 2836 35449 2839
rect 35400 2808 35449 2836
rect 35400 2796 35406 2808
rect 35437 2805 35449 2808
rect 35483 2805 35495 2839
rect 35437 2799 35495 2805
rect 36170 2796 36176 2848
rect 36228 2836 36234 2848
rect 36265 2839 36323 2845
rect 36265 2836 36277 2839
rect 36228 2808 36277 2836
rect 36228 2796 36234 2808
rect 36265 2805 36277 2808
rect 36311 2805 36323 2839
rect 36265 2799 36323 2805
rect 36722 2796 36728 2848
rect 36780 2836 36786 2848
rect 37277 2839 37335 2845
rect 37277 2836 37289 2839
rect 36780 2808 37289 2836
rect 36780 2796 36786 2808
rect 37277 2805 37289 2808
rect 37323 2805 37335 2839
rect 37277 2799 37335 2805
rect 37826 2796 37832 2848
rect 37884 2836 37890 2848
rect 38565 2839 38623 2845
rect 38565 2836 38577 2839
rect 37884 2808 38577 2836
rect 37884 2796 37890 2808
rect 38565 2805 38577 2808
rect 38611 2805 38623 2839
rect 38565 2799 38623 2805
rect 38930 2796 38936 2848
rect 38988 2836 38994 2848
rect 39853 2839 39911 2845
rect 39853 2836 39865 2839
rect 38988 2808 39865 2836
rect 38988 2796 38994 2808
rect 39853 2805 39865 2808
rect 39899 2805 39911 2839
rect 39853 2799 39911 2805
rect 40310 2796 40316 2848
rect 40368 2836 40374 2848
rect 41141 2839 41199 2845
rect 41141 2836 41153 2839
rect 40368 2808 41153 2836
rect 40368 2796 40374 2808
rect 41141 2805 41153 2808
rect 41187 2805 41199 2839
rect 41141 2799 41199 2805
rect 41690 2796 41696 2848
rect 41748 2836 41754 2848
rect 42429 2839 42487 2845
rect 42429 2836 42441 2839
rect 41748 2808 42441 2836
rect 41748 2796 41754 2808
rect 42429 2805 42441 2808
rect 42475 2805 42487 2839
rect 42429 2799 42487 2805
rect 42794 2796 42800 2848
rect 42852 2836 42858 2848
rect 43717 2839 43775 2845
rect 43717 2836 43729 2839
rect 42852 2808 43729 2836
rect 42852 2796 42858 2808
rect 43717 2805 43729 2808
rect 43763 2805 43775 2839
rect 43717 2799 43775 2805
rect 44174 2796 44180 2848
rect 44232 2836 44238 2848
rect 45005 2839 45063 2845
rect 45005 2836 45017 2839
rect 44232 2808 45017 2836
rect 44232 2796 44238 2808
rect 45005 2805 45017 2808
rect 45051 2805 45063 2839
rect 45005 2799 45063 2805
rect 45554 2796 45560 2848
rect 45612 2836 45618 2848
rect 46293 2839 46351 2845
rect 46293 2836 46305 2839
rect 45612 2808 46305 2836
rect 45612 2796 45618 2808
rect 46293 2805 46305 2808
rect 46339 2805 46351 2839
rect 46293 2799 46351 2805
rect 46658 2796 46664 2848
rect 46716 2836 46722 2848
rect 47581 2839 47639 2845
rect 47581 2836 47593 2839
rect 46716 2808 47593 2836
rect 46716 2796 46722 2808
rect 47581 2805 47593 2808
rect 47627 2805 47639 2839
rect 47581 2799 47639 2805
rect 48038 2796 48044 2848
rect 48096 2836 48102 2848
rect 48869 2839 48927 2845
rect 48869 2836 48881 2839
rect 48096 2808 48881 2836
rect 48096 2796 48102 2808
rect 48869 2805 48881 2808
rect 48915 2805 48927 2839
rect 48869 2799 48927 2805
rect 49970 2796 49976 2848
rect 50028 2836 50034 2848
rect 50801 2839 50859 2845
rect 50801 2836 50813 2839
rect 50028 2808 50813 2836
rect 50028 2796 50034 2808
rect 50801 2805 50813 2808
rect 50847 2805 50859 2839
rect 50801 2799 50859 2805
rect 51902 2796 51908 2848
rect 51960 2836 51966 2848
rect 52733 2839 52791 2845
rect 52733 2836 52745 2839
rect 51960 2808 52745 2836
rect 51960 2796 51966 2808
rect 52733 2805 52745 2808
rect 52779 2805 52791 2839
rect 52733 2799 52791 2805
rect 53834 2796 53840 2848
rect 53892 2836 53898 2848
rect 54665 2839 54723 2845
rect 54665 2836 54677 2839
rect 53892 2808 54677 2836
rect 53892 2796 53898 2808
rect 54665 2805 54677 2808
rect 54711 2805 54723 2839
rect 54665 2799 54723 2805
rect 55398 2796 55404 2848
rect 55456 2836 55462 2848
rect 55953 2839 56011 2845
rect 55953 2836 55965 2839
rect 55456 2808 55965 2836
rect 55456 2796 55462 2808
rect 55953 2805 55965 2808
rect 55999 2805 56011 2839
rect 55953 2799 56011 2805
rect 56042 2796 56048 2848
rect 56100 2836 56106 2848
rect 57885 2839 57943 2845
rect 57885 2836 57897 2839
rect 56100 2808 57897 2836
rect 56100 2796 56106 2808
rect 57885 2805 57897 2808
rect 57931 2805 57943 2839
rect 57992 2836 58020 2876
rect 58529 2873 58541 2876
rect 58575 2873 58587 2907
rect 58529 2867 58587 2873
rect 59354 2864 59360 2916
rect 59412 2904 59418 2916
rect 63037 2907 63095 2913
rect 63037 2904 63049 2907
rect 59412 2876 63049 2904
rect 59412 2864 59418 2876
rect 63037 2873 63049 2876
rect 63083 2873 63095 2907
rect 63037 2867 63095 2873
rect 59173 2839 59231 2845
rect 59173 2836 59185 2839
rect 57992 2808 59185 2836
rect 57885 2799 57943 2805
rect 59173 2805 59185 2808
rect 59219 2805 59231 2839
rect 59173 2799 59231 2805
rect 59446 2796 59452 2848
rect 59504 2836 59510 2848
rect 59817 2839 59875 2845
rect 59817 2836 59829 2839
rect 59504 2808 59829 2836
rect 59504 2796 59510 2808
rect 59817 2805 59829 2808
rect 59863 2805 59875 2839
rect 60458 2836 60464 2848
rect 60419 2808 60464 2836
rect 59817 2799 59875 2805
rect 60458 2796 60464 2808
rect 60516 2796 60522 2848
rect 1104 2746 68816 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 65654 2746
rect 65706 2694 65718 2746
rect 65770 2694 65782 2746
rect 65834 2694 65846 2746
rect 65898 2694 65910 2746
rect 65962 2694 68816 2746
rect 1104 2672 68816 2694
rect 1949 2635 2007 2641
rect 1949 2601 1961 2635
rect 1995 2632 2007 2635
rect 8294 2632 8300 2644
rect 1995 2604 8300 2632
rect 1995 2601 2007 2604
rect 1949 2595 2007 2601
rect 8294 2592 8300 2604
rect 8352 2592 8358 2644
rect 9861 2635 9919 2641
rect 9861 2601 9873 2635
rect 9907 2632 9919 2635
rect 10410 2632 10416 2644
rect 9907 2604 10416 2632
rect 9907 2601 9919 2604
rect 9861 2595 9919 2601
rect 10410 2592 10416 2604
rect 10468 2592 10474 2644
rect 10502 2592 10508 2644
rect 10560 2632 10566 2644
rect 12802 2632 12808 2644
rect 10560 2604 12808 2632
rect 10560 2592 10566 2604
rect 12802 2592 12808 2604
rect 12860 2592 12866 2644
rect 14826 2632 14832 2644
rect 14787 2604 14832 2632
rect 14826 2592 14832 2604
rect 14884 2592 14890 2644
rect 17497 2635 17555 2641
rect 17497 2601 17509 2635
rect 17543 2632 17555 2635
rect 17954 2632 17960 2644
rect 17543 2604 17960 2632
rect 17543 2601 17555 2604
rect 17497 2595 17555 2601
rect 17954 2592 17960 2604
rect 18012 2592 18018 2644
rect 24397 2635 24455 2641
rect 24397 2632 24409 2635
rect 18064 2604 24409 2632
rect 5629 2567 5687 2573
rect 5629 2533 5641 2567
rect 5675 2564 5687 2567
rect 10778 2564 10784 2576
rect 5675 2536 10784 2564
rect 5675 2533 5687 2536
rect 5629 2527 5687 2533
rect 10778 2524 10784 2536
rect 10836 2524 10842 2576
rect 11054 2524 11060 2576
rect 11112 2564 11118 2576
rect 12434 2564 12440 2576
rect 11112 2536 12440 2564
rect 11112 2524 11118 2536
rect 12434 2524 12440 2536
rect 12492 2524 12498 2576
rect 14458 2524 14464 2576
rect 14516 2564 14522 2576
rect 15933 2567 15991 2573
rect 15933 2564 15945 2567
rect 14516 2536 15945 2564
rect 14516 2524 14522 2536
rect 15933 2533 15945 2536
rect 15979 2533 15991 2567
rect 15933 2527 15991 2533
rect 17586 2524 17592 2576
rect 17644 2564 17650 2576
rect 18064 2564 18092 2604
rect 24397 2601 24409 2604
rect 24443 2601 24455 2635
rect 24397 2595 24455 2601
rect 55214 2592 55220 2644
rect 55272 2632 55278 2644
rect 55309 2635 55367 2641
rect 55309 2632 55321 2635
rect 55272 2604 55321 2632
rect 55272 2592 55278 2604
rect 55309 2601 55321 2604
rect 55355 2601 55367 2635
rect 55309 2595 55367 2601
rect 57422 2592 57428 2644
rect 57480 2632 57486 2644
rect 61105 2635 61163 2641
rect 61105 2632 61117 2635
rect 57480 2604 61117 2632
rect 57480 2592 57486 2604
rect 61105 2601 61117 2604
rect 61151 2601 61163 2635
rect 61105 2595 61163 2601
rect 17644 2536 18092 2564
rect 18325 2567 18383 2573
rect 17644 2524 17650 2536
rect 18325 2533 18337 2567
rect 18371 2533 18383 2567
rect 18325 2527 18383 2533
rect 19981 2567 20039 2573
rect 19981 2533 19993 2567
rect 20027 2564 20039 2567
rect 21542 2564 21548 2576
rect 20027 2536 21548 2564
rect 20027 2533 20039 2536
rect 19981 2527 20039 2533
rect 5166 2496 5172 2508
rect 4264 2468 5172 2496
rect 1762 2428 1768 2440
rect 1723 2400 1768 2428
rect 1762 2388 1768 2400
rect 1820 2388 1826 2440
rect 2409 2431 2467 2437
rect 2409 2397 2421 2431
rect 2455 2428 2467 2431
rect 2498 2428 2504 2440
rect 2455 2400 2504 2428
rect 2455 2397 2467 2400
rect 2409 2391 2467 2397
rect 2498 2388 2504 2400
rect 2556 2388 2562 2440
rect 2958 2388 2964 2440
rect 3016 2428 3022 2440
rect 4264 2437 4292 2468
rect 5166 2456 5172 2468
rect 5224 2456 5230 2508
rect 8478 2496 8484 2508
rect 6932 2468 8484 2496
rect 3053 2431 3111 2437
rect 3053 2428 3065 2431
rect 3016 2400 3065 2428
rect 3016 2388 3022 2400
rect 3053 2397 3065 2400
rect 3099 2397 3111 2431
rect 3053 2391 3111 2397
rect 4249 2431 4307 2437
rect 4249 2397 4261 2431
rect 4295 2397 4307 2431
rect 4890 2428 4896 2440
rect 4851 2400 4896 2428
rect 4249 2391 4307 2397
rect 4890 2388 4896 2400
rect 4948 2388 4954 2440
rect 5813 2431 5871 2437
rect 5813 2397 5825 2431
rect 5859 2428 5871 2431
rect 6362 2428 6368 2440
rect 5859 2400 6368 2428
rect 5859 2397 5871 2400
rect 5813 2391 5871 2397
rect 6362 2388 6368 2400
rect 6420 2388 6426 2440
rect 6932 2437 6960 2468
rect 8478 2456 8484 2468
rect 8536 2456 8542 2508
rect 10042 2456 10048 2508
rect 10100 2496 10106 2508
rect 10597 2499 10655 2505
rect 10597 2496 10609 2499
rect 10100 2468 10609 2496
rect 10100 2456 10106 2468
rect 10597 2465 10609 2468
rect 10643 2465 10655 2499
rect 10597 2459 10655 2465
rect 11072 2468 11652 2496
rect 6917 2431 6975 2437
rect 6917 2397 6929 2431
rect 6963 2397 6975 2431
rect 7650 2428 7656 2440
rect 7611 2400 7656 2428
rect 6917 2391 6975 2397
rect 7650 2388 7656 2400
rect 7708 2388 7714 2440
rect 8389 2431 8447 2437
rect 8128 2400 8340 2428
rect 4338 2360 4344 2372
rect 2608 2332 4344 2360
rect 2608 2301 2636 2332
rect 4338 2320 4344 2332
rect 4396 2320 4402 2372
rect 7190 2360 7196 2372
rect 4448 2332 7196 2360
rect 2593 2295 2651 2301
rect 2593 2261 2605 2295
rect 2639 2261 2651 2295
rect 3234 2292 3240 2304
rect 3195 2264 3240 2292
rect 2593 2255 2651 2261
rect 3234 2252 3240 2264
rect 3292 2252 3298 2304
rect 4448 2301 4476 2332
rect 7190 2320 7196 2332
rect 7248 2320 7254 2372
rect 8128 2360 8156 2400
rect 7484 2332 8156 2360
rect 8312 2360 8340 2400
rect 8389 2397 8401 2431
rect 8435 2428 8447 2431
rect 8754 2428 8760 2440
rect 8435 2400 8760 2428
rect 8435 2397 8447 2400
rect 8389 2391 8447 2397
rect 8754 2388 8760 2400
rect 8812 2388 8818 2440
rect 9122 2428 9128 2440
rect 9083 2400 9128 2428
rect 9122 2388 9128 2400
rect 9180 2388 9186 2440
rect 10502 2428 10508 2440
rect 9232 2400 10508 2428
rect 8312 2332 8432 2360
rect 4433 2295 4491 2301
rect 4433 2261 4445 2295
rect 4479 2261 4491 2295
rect 5074 2292 5080 2304
rect 5035 2264 5080 2292
rect 4433 2255 4491 2261
rect 5074 2252 5080 2264
rect 5132 2252 5138 2304
rect 6730 2292 6736 2304
rect 6691 2264 6736 2292
rect 6730 2252 6736 2264
rect 6788 2252 6794 2304
rect 7484 2301 7512 2332
rect 7469 2295 7527 2301
rect 7469 2261 7481 2295
rect 7515 2261 7527 2295
rect 7469 2255 7527 2261
rect 8202 2252 8208 2304
rect 8260 2292 8266 2304
rect 8404 2292 8432 2332
rect 8478 2320 8484 2372
rect 8536 2360 8542 2372
rect 9232 2360 9260 2400
rect 10502 2388 10508 2400
rect 10560 2388 10566 2440
rect 10612 2428 10640 2459
rect 11072 2428 11100 2468
rect 10612 2400 11100 2428
rect 11146 2388 11152 2440
rect 11204 2428 11210 2440
rect 11517 2431 11575 2437
rect 11517 2428 11529 2431
rect 11204 2400 11529 2428
rect 11204 2388 11210 2400
rect 11517 2397 11529 2400
rect 11563 2397 11575 2431
rect 11624 2428 11652 2468
rect 11698 2456 11704 2508
rect 11756 2496 11762 2508
rect 11793 2499 11851 2505
rect 11793 2496 11805 2499
rect 11756 2468 11805 2496
rect 11756 2456 11762 2468
rect 11793 2465 11805 2468
rect 11839 2465 11851 2499
rect 11793 2459 11851 2465
rect 12158 2456 12164 2508
rect 12216 2496 12222 2508
rect 13538 2496 13544 2508
rect 12216 2468 13544 2496
rect 12216 2456 12222 2468
rect 13538 2456 13544 2468
rect 13596 2456 13602 2508
rect 18340 2496 18368 2527
rect 21542 2524 21548 2536
rect 21600 2524 21606 2576
rect 22557 2567 22615 2573
rect 22557 2533 22569 2567
rect 22603 2564 22615 2567
rect 24026 2564 24032 2576
rect 22603 2536 24032 2564
rect 22603 2533 22615 2536
rect 22557 2527 22615 2533
rect 24026 2524 24032 2536
rect 24084 2524 24090 2576
rect 25777 2567 25835 2573
rect 25777 2533 25789 2567
rect 25823 2564 25835 2567
rect 27338 2564 27344 2576
rect 25823 2536 27344 2564
rect 25823 2533 25835 2536
rect 25777 2527 25835 2533
rect 27338 2524 27344 2536
rect 27396 2524 27402 2576
rect 31573 2567 31631 2573
rect 31573 2533 31585 2567
rect 31619 2564 31631 2567
rect 32858 2564 32864 2576
rect 31619 2536 32864 2564
rect 31619 2533 31631 2536
rect 31573 2527 31631 2533
rect 32858 2524 32864 2536
rect 32916 2524 32922 2576
rect 40586 2524 40592 2576
rect 40644 2564 40650 2576
rect 42429 2567 42487 2573
rect 42429 2564 42441 2567
rect 40644 2536 42441 2564
rect 40644 2524 40650 2536
rect 42429 2533 42441 2536
rect 42475 2533 42487 2567
rect 42429 2527 42487 2533
rect 44450 2524 44456 2576
rect 44508 2564 44514 2576
rect 46293 2567 46351 2573
rect 46293 2564 46305 2567
rect 44508 2536 46305 2564
rect 44508 2524 44514 2536
rect 46293 2533 46305 2536
rect 46339 2533 46351 2567
rect 46293 2527 46351 2533
rect 48314 2524 48320 2576
rect 48372 2564 48378 2576
rect 50157 2567 50215 2573
rect 50157 2564 50169 2567
rect 48372 2536 50169 2564
rect 48372 2524 48378 2536
rect 50157 2533 50169 2536
rect 50203 2533 50215 2567
rect 50157 2527 50215 2533
rect 52178 2524 52184 2576
rect 52236 2564 52242 2576
rect 54021 2567 54079 2573
rect 54021 2564 54033 2567
rect 52236 2536 54033 2564
rect 52236 2524 52242 2536
rect 54021 2533 54033 2536
rect 54067 2533 54079 2567
rect 54021 2527 54079 2533
rect 55858 2524 55864 2576
rect 55916 2564 55922 2576
rect 57885 2567 57943 2573
rect 57885 2564 57897 2567
rect 55916 2536 57897 2564
rect 55916 2524 55922 2536
rect 57885 2533 57897 2536
rect 57931 2533 57943 2567
rect 57885 2527 57943 2533
rect 58066 2524 58072 2576
rect 58124 2564 58130 2576
rect 58529 2567 58587 2573
rect 58529 2564 58541 2567
rect 58124 2536 58541 2564
rect 58124 2524 58130 2536
rect 58529 2533 58541 2536
rect 58575 2533 58587 2567
rect 58529 2527 58587 2533
rect 60461 2567 60519 2573
rect 60461 2533 60473 2567
rect 60507 2533 60519 2567
rect 60461 2527 60519 2533
rect 20625 2499 20683 2505
rect 13740 2468 18368 2496
rect 18524 2468 20576 2496
rect 13170 2428 13176 2440
rect 11624 2400 13176 2428
rect 11517 2391 11575 2397
rect 13170 2388 13176 2400
rect 13228 2388 13234 2440
rect 13740 2428 13768 2468
rect 13556 2400 13768 2428
rect 13556 2372 13584 2400
rect 14918 2388 14924 2440
rect 14976 2428 14982 2440
rect 15749 2431 15807 2437
rect 15749 2428 15761 2431
rect 14976 2400 15761 2428
rect 14976 2388 14982 2400
rect 15749 2397 15761 2400
rect 15795 2397 15807 2431
rect 16945 2431 17003 2437
rect 16945 2428 16957 2431
rect 15749 2391 15807 2397
rect 16684 2400 16957 2428
rect 8536 2332 9260 2360
rect 8536 2320 8542 2332
rect 9950 2320 9956 2372
rect 10008 2360 10014 2372
rect 10873 2363 10931 2369
rect 10008 2332 10053 2360
rect 10008 2320 10014 2332
rect 10873 2329 10885 2363
rect 10919 2360 10931 2363
rect 11882 2360 11888 2372
rect 10919 2332 11888 2360
rect 10919 2329 10931 2332
rect 10873 2323 10931 2329
rect 11882 2320 11888 2332
rect 11940 2320 11946 2372
rect 12710 2320 12716 2372
rect 12768 2360 12774 2372
rect 12897 2363 12955 2369
rect 12897 2360 12909 2363
rect 12768 2332 12909 2360
rect 12768 2320 12774 2332
rect 12897 2329 12909 2332
rect 12943 2329 12955 2363
rect 12897 2323 12955 2329
rect 13538 2320 13544 2372
rect 13596 2320 13602 2372
rect 13722 2320 13728 2372
rect 13780 2360 13786 2372
rect 14553 2363 14611 2369
rect 14553 2360 14565 2363
rect 13780 2332 14565 2360
rect 13780 2320 13786 2332
rect 14553 2329 14565 2332
rect 14599 2329 14611 2363
rect 14553 2323 14611 2329
rect 11054 2292 11060 2304
rect 8260 2264 8305 2292
rect 8404 2264 11060 2292
rect 8260 2252 8266 2264
rect 11054 2252 11060 2264
rect 11112 2252 11118 2304
rect 12986 2292 12992 2304
rect 12947 2264 12992 2292
rect 12986 2252 12992 2264
rect 13044 2252 13050 2304
rect 14090 2252 14096 2304
rect 14148 2292 14154 2304
rect 16684 2292 16712 2400
rect 16945 2397 16957 2400
rect 16991 2397 17003 2431
rect 18138 2428 18144 2440
rect 18099 2400 18144 2428
rect 16945 2391 17003 2397
rect 14148 2264 16712 2292
rect 14148 2252 14154 2264
rect 16758 2252 16764 2304
rect 16816 2292 16822 2304
rect 16960 2292 16988 2391
rect 18138 2388 18144 2400
rect 18196 2388 18202 2440
rect 17586 2360 17592 2372
rect 17547 2332 17592 2360
rect 17586 2320 17592 2332
rect 17644 2360 17650 2372
rect 18524 2360 18552 2468
rect 20548 2428 20576 2468
rect 20625 2465 20637 2499
rect 20671 2496 20683 2499
rect 22094 2496 22100 2508
rect 20671 2468 22100 2496
rect 20671 2465 20683 2468
rect 20625 2459 20683 2465
rect 22094 2456 22100 2468
rect 22152 2456 22158 2508
rect 23201 2499 23259 2505
rect 23201 2465 23213 2499
rect 23247 2496 23259 2499
rect 24578 2496 24584 2508
rect 23247 2468 24584 2496
rect 23247 2465 23259 2468
rect 23201 2459 23259 2465
rect 24578 2456 24584 2468
rect 24636 2456 24642 2508
rect 25133 2499 25191 2505
rect 25133 2465 25145 2499
rect 25179 2496 25191 2499
rect 26510 2496 26516 2508
rect 25179 2468 26516 2496
rect 25179 2465 25191 2468
rect 25133 2459 25191 2465
rect 26510 2456 26516 2468
rect 26568 2456 26574 2508
rect 27709 2499 27767 2505
rect 27709 2465 27721 2499
rect 27755 2496 27767 2499
rect 28442 2496 28448 2508
rect 27755 2468 28448 2496
rect 27755 2465 27767 2468
rect 27709 2459 27767 2465
rect 28442 2456 28448 2468
rect 28500 2456 28506 2508
rect 28997 2499 29055 2505
rect 28997 2465 29009 2499
rect 29043 2496 29055 2499
rect 30374 2496 30380 2508
rect 29043 2468 30380 2496
rect 29043 2465 29055 2468
rect 28997 2459 29055 2465
rect 30374 2456 30380 2468
rect 30432 2456 30438 2508
rect 36998 2456 37004 2508
rect 37056 2496 37062 2508
rect 37921 2499 37979 2505
rect 37921 2496 37933 2499
rect 37056 2468 37933 2496
rect 37056 2456 37062 2468
rect 37921 2465 37933 2468
rect 37967 2465 37979 2499
rect 37921 2459 37979 2465
rect 38102 2456 38108 2508
rect 38160 2496 38166 2508
rect 39853 2499 39911 2505
rect 39853 2496 39865 2499
rect 38160 2468 39865 2496
rect 38160 2456 38166 2468
rect 39853 2465 39865 2468
rect 39899 2465 39911 2499
rect 39853 2459 39911 2465
rect 41414 2456 41420 2508
rect 41472 2496 41478 2508
rect 43073 2499 43131 2505
rect 43073 2496 43085 2499
rect 41472 2468 43085 2496
rect 41472 2456 41478 2468
rect 43073 2465 43085 2468
rect 43119 2465 43131 2499
rect 43073 2459 43131 2465
rect 43346 2456 43352 2508
rect 43404 2496 43410 2508
rect 45005 2499 45063 2505
rect 45005 2496 45017 2499
rect 43404 2468 45017 2496
rect 43404 2456 43410 2468
rect 45005 2465 45017 2468
rect 45051 2465 45063 2499
rect 45005 2459 45063 2465
rect 46382 2456 46388 2508
rect 46440 2496 46446 2508
rect 48225 2499 48283 2505
rect 48225 2496 48237 2499
rect 46440 2468 48237 2496
rect 46440 2456 46446 2468
rect 48225 2465 48237 2468
rect 48271 2465 48283 2499
rect 48225 2459 48283 2465
rect 49142 2456 49148 2508
rect 49200 2496 49206 2508
rect 50801 2499 50859 2505
rect 50801 2496 50813 2499
rect 49200 2468 50813 2496
rect 49200 2456 49206 2468
rect 50801 2465 50813 2468
rect 50847 2465 50859 2499
rect 50801 2459 50859 2465
rect 51074 2456 51080 2508
rect 51132 2496 51138 2508
rect 52733 2499 52791 2505
rect 52733 2496 52745 2499
rect 51132 2468 52745 2496
rect 51132 2456 51138 2468
rect 52733 2465 52745 2468
rect 52779 2465 52791 2499
rect 52733 2459 52791 2465
rect 54938 2456 54944 2508
rect 54996 2496 55002 2508
rect 56597 2499 56655 2505
rect 56597 2496 56609 2499
rect 54996 2468 56609 2496
rect 54996 2456 55002 2468
rect 56597 2465 56609 2468
rect 56643 2465 56655 2499
rect 60476 2496 60504 2527
rect 63678 2496 63684 2508
rect 60476 2468 60596 2496
rect 63639 2468 63684 2496
rect 56597 2459 56655 2465
rect 21269 2431 21327 2437
rect 20548 2400 20668 2428
rect 20530 2360 20536 2372
rect 17644 2332 18552 2360
rect 18708 2332 20536 2360
rect 17644 2320 17650 2332
rect 18708 2292 18736 2332
rect 20530 2320 20536 2332
rect 20588 2320 20594 2372
rect 20640 2360 20668 2400
rect 21269 2397 21281 2431
rect 21315 2428 21327 2431
rect 22922 2428 22928 2440
rect 21315 2400 22928 2428
rect 21315 2397 21327 2400
rect 21269 2391 21327 2397
rect 22922 2388 22928 2400
rect 22980 2388 22986 2440
rect 23845 2431 23903 2437
rect 23845 2397 23857 2431
rect 23891 2428 23903 2431
rect 25406 2428 25412 2440
rect 23891 2400 25412 2428
rect 23891 2397 23903 2400
rect 23845 2391 23903 2397
rect 25406 2388 25412 2400
rect 25464 2388 25470 2440
rect 26421 2431 26479 2437
rect 26421 2397 26433 2431
rect 26467 2428 26479 2431
rect 27614 2428 27620 2440
rect 26467 2400 27620 2428
rect 26467 2397 26479 2400
rect 26421 2391 26479 2397
rect 27614 2388 27620 2400
rect 27672 2388 27678 2440
rect 28353 2431 28411 2437
rect 28353 2397 28365 2431
rect 28399 2428 28411 2431
rect 29822 2428 29828 2440
rect 28399 2400 29828 2428
rect 28399 2397 28411 2400
rect 28353 2391 28411 2397
rect 29822 2388 29828 2400
rect 29880 2388 29886 2440
rect 30285 2431 30343 2437
rect 30285 2397 30297 2431
rect 30331 2397 30343 2431
rect 30285 2391 30343 2397
rect 30929 2431 30987 2437
rect 30929 2397 30941 2431
rect 30975 2428 30987 2431
rect 32306 2428 32312 2440
rect 30975 2400 32312 2428
rect 30975 2397 30987 2400
rect 30929 2391 30987 2397
rect 26973 2363 27031 2369
rect 26973 2360 26985 2363
rect 20640 2332 26985 2360
rect 26973 2329 26985 2332
rect 27019 2329 27031 2363
rect 30300 2360 30328 2391
rect 32306 2388 32312 2400
rect 32364 2388 32370 2440
rect 32861 2431 32919 2437
rect 32861 2397 32873 2431
rect 32907 2428 32919 2431
rect 33410 2428 33416 2440
rect 32907 2400 33416 2428
rect 32907 2397 32919 2400
rect 32861 2391 32919 2397
rect 33410 2388 33416 2400
rect 33468 2388 33474 2440
rect 33505 2431 33563 2437
rect 33505 2397 33517 2431
rect 33551 2428 33563 2431
rect 33962 2428 33968 2440
rect 33551 2400 33968 2428
rect 33551 2397 33563 2400
rect 33505 2391 33563 2397
rect 33962 2388 33968 2400
rect 34020 2388 34026 2440
rect 34149 2431 34207 2437
rect 34149 2397 34161 2431
rect 34195 2428 34207 2431
rect 34790 2428 34796 2440
rect 34195 2400 34796 2428
rect 34195 2397 34207 2400
rect 34149 2391 34207 2397
rect 34790 2388 34796 2400
rect 34848 2388 34854 2440
rect 34885 2431 34943 2437
rect 34885 2397 34897 2431
rect 34931 2428 34943 2431
rect 35066 2428 35072 2440
rect 34931 2400 35072 2428
rect 34931 2397 34943 2400
rect 34885 2391 34943 2397
rect 35066 2388 35072 2400
rect 35124 2388 35130 2440
rect 35529 2431 35587 2437
rect 35529 2397 35541 2431
rect 35575 2428 35587 2431
rect 35618 2428 35624 2440
rect 35575 2400 35624 2428
rect 35575 2397 35587 2400
rect 35529 2391 35587 2397
rect 35618 2388 35624 2400
rect 35676 2388 35682 2440
rect 35894 2388 35900 2440
rect 35952 2428 35958 2440
rect 35989 2431 36047 2437
rect 35989 2428 36001 2431
rect 35952 2400 36001 2428
rect 35952 2388 35958 2400
rect 35989 2397 36001 2400
rect 36035 2397 36047 2431
rect 35989 2391 36047 2397
rect 36446 2388 36452 2440
rect 36504 2428 36510 2440
rect 37277 2431 37335 2437
rect 37277 2428 37289 2431
rect 36504 2400 37289 2428
rect 36504 2388 36510 2400
rect 37277 2397 37289 2400
rect 37323 2397 37335 2431
rect 37277 2391 37335 2397
rect 37550 2388 37556 2440
rect 37608 2428 37614 2440
rect 38565 2431 38623 2437
rect 38565 2428 38577 2431
rect 37608 2400 38577 2428
rect 37608 2388 37614 2400
rect 38565 2397 38577 2400
rect 38611 2397 38623 2431
rect 38565 2391 38623 2397
rect 38654 2388 38660 2440
rect 38712 2428 38718 2440
rect 40497 2431 40555 2437
rect 40497 2428 40509 2431
rect 38712 2400 40509 2428
rect 38712 2388 38718 2400
rect 40497 2397 40509 2400
rect 40543 2397 40555 2431
rect 40497 2391 40555 2397
rect 41141 2431 41199 2437
rect 41141 2397 41153 2431
rect 41187 2397 41199 2431
rect 41141 2391 41199 2397
rect 31754 2360 31760 2372
rect 30300 2332 31760 2360
rect 26973 2323 27031 2329
rect 31754 2320 31760 2332
rect 31812 2320 31818 2372
rect 39482 2320 39488 2372
rect 39540 2360 39546 2372
rect 41156 2360 41184 2391
rect 41966 2388 41972 2440
rect 42024 2428 42030 2440
rect 43717 2431 43775 2437
rect 43717 2428 43729 2431
rect 42024 2400 43729 2428
rect 42024 2388 42030 2400
rect 43717 2397 43729 2400
rect 43763 2397 43775 2431
rect 45649 2431 45707 2437
rect 45649 2428 45661 2431
rect 43717 2391 43775 2397
rect 45526 2400 45661 2428
rect 39540 2332 41184 2360
rect 39540 2320 39546 2332
rect 43898 2320 43904 2372
rect 43956 2360 43962 2372
rect 45526 2360 45554 2400
rect 45649 2397 45661 2400
rect 45695 2397 45707 2431
rect 45649 2391 45707 2397
rect 45830 2388 45836 2440
rect 45888 2428 45894 2440
rect 47581 2431 47639 2437
rect 47581 2428 47593 2431
rect 45888 2400 47593 2428
rect 45888 2388 45894 2400
rect 47581 2397 47593 2400
rect 47627 2397 47639 2431
rect 47581 2391 47639 2397
rect 48869 2431 48927 2437
rect 48869 2397 48881 2431
rect 48915 2397 48927 2431
rect 48869 2391 48927 2397
rect 43956 2332 45554 2360
rect 43956 2320 43962 2332
rect 47210 2320 47216 2372
rect 47268 2360 47274 2372
rect 48884 2360 48912 2391
rect 49694 2388 49700 2440
rect 49752 2428 49758 2440
rect 51445 2431 51503 2437
rect 51445 2428 51457 2431
rect 49752 2400 51457 2428
rect 49752 2388 49758 2400
rect 51445 2397 51457 2400
rect 51491 2397 51503 2431
rect 51445 2391 51503 2397
rect 51626 2388 51632 2440
rect 51684 2428 51690 2440
rect 53377 2431 53435 2437
rect 53377 2428 53389 2431
rect 51684 2400 53389 2428
rect 51684 2388 51690 2400
rect 53377 2397 53389 2400
rect 53423 2397 53435 2431
rect 53377 2391 53435 2397
rect 55953 2431 56011 2437
rect 55953 2397 55965 2431
rect 55999 2397 56011 2431
rect 55953 2391 56011 2397
rect 47268 2332 48912 2360
rect 47268 2320 47274 2332
rect 54110 2320 54116 2372
rect 54168 2360 54174 2372
rect 55968 2360 55996 2391
rect 56410 2388 56416 2440
rect 56468 2428 56474 2440
rect 59173 2431 59231 2437
rect 59173 2428 59185 2431
rect 56468 2400 59185 2428
rect 56468 2388 56474 2400
rect 59173 2397 59185 2400
rect 59219 2397 59231 2431
rect 59173 2391 59231 2397
rect 54168 2332 55996 2360
rect 54168 2320 54174 2332
rect 16816 2264 16861 2292
rect 16960 2264 18736 2292
rect 16816 2252 16822 2264
rect 18782 2252 18788 2304
rect 18840 2292 18846 2304
rect 19242 2292 19248 2304
rect 18840 2264 19248 2292
rect 18840 2252 18846 2264
rect 19242 2252 19248 2264
rect 19300 2292 19306 2304
rect 19337 2295 19395 2301
rect 19337 2292 19349 2295
rect 19300 2264 19349 2292
rect 19300 2252 19306 2264
rect 19337 2261 19349 2264
rect 19383 2261 19395 2295
rect 19337 2255 19395 2261
rect 20622 2252 20628 2304
rect 20680 2292 20686 2304
rect 21821 2295 21879 2301
rect 21821 2292 21833 2295
rect 20680 2264 21833 2292
rect 20680 2252 20686 2264
rect 21821 2261 21833 2264
rect 21867 2261 21879 2295
rect 21821 2255 21879 2261
rect 56870 2252 56876 2304
rect 56928 2292 56934 2304
rect 60568 2292 60596 2468
rect 63678 2456 63684 2468
rect 63736 2456 63742 2508
rect 61746 2428 61752 2440
rect 61707 2400 61752 2428
rect 61746 2388 61752 2400
rect 61804 2388 61810 2440
rect 63034 2428 63040 2440
rect 62995 2400 63040 2428
rect 63034 2388 63040 2400
rect 63092 2388 63098 2440
rect 66990 2428 66996 2440
rect 66951 2400 66996 2428
rect 66990 2388 66996 2400
rect 67048 2388 67054 2440
rect 67542 2388 67548 2440
rect 67600 2428 67606 2440
rect 67637 2431 67695 2437
rect 67637 2428 67649 2431
rect 67600 2400 67649 2428
rect 67600 2388 67606 2400
rect 67637 2397 67649 2400
rect 67683 2397 67695 2431
rect 67637 2391 67695 2397
rect 56928 2264 60596 2292
rect 56928 2252 56934 2264
rect 1104 2202 68816 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 68816 2202
rect 1104 2128 68816 2150
rect 6730 2048 6736 2100
rect 6788 2088 6794 2100
rect 11698 2088 11704 2100
rect 6788 2060 11704 2088
rect 6788 2048 6794 2060
rect 11698 2048 11704 2060
rect 11756 2048 11762 2100
rect 13170 2048 13176 2100
rect 13228 2088 13234 2100
rect 20346 2088 20352 2100
rect 13228 2060 20352 2088
rect 13228 2048 13234 2060
rect 20346 2048 20352 2060
rect 20404 2048 20410 2100
rect 58066 2048 58072 2100
rect 58124 2088 58130 2100
rect 61746 2088 61752 2100
rect 58124 2060 61752 2088
rect 58124 2048 58130 2060
rect 61746 2048 61752 2060
rect 61804 2048 61810 2100
rect 5074 1980 5080 2032
rect 5132 2020 5138 2032
rect 12158 2020 12164 2032
rect 5132 1992 12164 2020
rect 5132 1980 5138 1992
rect 12158 1980 12164 1992
rect 12216 1980 12222 2032
rect 12342 1980 12348 2032
rect 12400 2020 12406 2032
rect 13722 2020 13728 2032
rect 12400 1992 13728 2020
rect 12400 1980 12406 1992
rect 13722 1980 13728 1992
rect 13780 1980 13786 2032
rect 16758 1980 16764 2032
rect 16816 2020 16822 2032
rect 22738 2020 22744 2032
rect 16816 1992 22744 2020
rect 16816 1980 16822 1992
rect 22738 1980 22744 1992
rect 22796 1980 22802 2032
rect 59078 1980 59084 2032
rect 59136 2020 59142 2032
rect 63678 2020 63684 2032
rect 59136 1992 63684 2020
rect 59136 1980 59142 1992
rect 63678 1980 63684 1992
rect 63736 1980 63742 2032
rect 8846 1912 8852 1964
rect 8904 1952 8910 1964
rect 9950 1952 9956 1964
rect 8904 1924 9956 1952
rect 8904 1912 8910 1924
rect 9950 1912 9956 1924
rect 10008 1952 10014 1964
rect 11238 1952 11244 1964
rect 10008 1924 11244 1952
rect 10008 1912 10014 1924
rect 11238 1912 11244 1924
rect 11296 1912 11302 1964
rect 58526 1912 58532 1964
rect 58584 1952 58590 1964
rect 63034 1952 63040 1964
rect 58584 1924 63040 1952
rect 58584 1912 58590 1924
rect 63034 1912 63040 1924
rect 63092 1912 63098 1964
rect 9122 1844 9128 1896
rect 9180 1884 9186 1896
rect 16666 1884 16672 1896
rect 9180 1856 16672 1884
rect 9180 1844 9186 1856
rect 16666 1844 16672 1856
rect 16724 1844 16730 1896
rect 4338 1776 4344 1828
rect 4396 1816 4402 1828
rect 9858 1816 9864 1828
rect 4396 1788 9864 1816
rect 4396 1776 4402 1788
rect 9858 1776 9864 1788
rect 9916 1776 9922 1828
rect 3234 1708 3240 1760
rect 3292 1748 3298 1760
rect 10594 1748 10600 1760
rect 3292 1720 10600 1748
rect 3292 1708 3298 1720
rect 10594 1708 10600 1720
rect 10652 1708 10658 1760
rect 19794 1708 19800 1760
rect 19852 1748 19858 1760
rect 20622 1748 20628 1760
rect 19852 1720 20628 1748
rect 19852 1708 19858 1720
rect 20622 1708 20628 1720
rect 20680 1708 20686 1760
rect 2958 1640 2964 1692
rect 3016 1680 3022 1692
rect 11054 1680 11060 1692
rect 3016 1652 11060 1680
rect 3016 1640 3022 1652
rect 11054 1640 11060 1652
rect 11112 1640 11118 1692
rect 12618 1368 12624 1420
rect 12676 1408 12682 1420
rect 13170 1408 13176 1420
rect 12676 1380 13176 1408
rect 12676 1368 12682 1380
rect 13170 1368 13176 1380
rect 13228 1368 13234 1420
rect 13538 1408 13544 1420
rect 13280 1380 13544 1408
rect 1762 1300 1768 1352
rect 1820 1340 1826 1352
rect 10318 1340 10324 1352
rect 1820 1312 10324 1340
rect 1820 1300 1826 1312
rect 10318 1300 10324 1312
rect 10376 1340 10382 1352
rect 10686 1340 10692 1352
rect 10376 1312 10692 1340
rect 10376 1300 10382 1312
rect 10686 1300 10692 1312
rect 10744 1300 10750 1352
rect 13078 1300 13084 1352
rect 13136 1340 13142 1352
rect 13280 1340 13308 1380
rect 13538 1368 13544 1380
rect 13596 1368 13602 1420
rect 17586 1408 17592 1420
rect 13648 1380 17592 1408
rect 13648 1340 13676 1380
rect 17586 1368 17592 1380
rect 17644 1368 17650 1420
rect 13136 1312 13308 1340
rect 13556 1312 13676 1340
rect 13136 1300 13142 1312
rect 13556 1284 13584 1312
rect 19518 1300 19524 1352
rect 19576 1340 19582 1352
rect 20162 1340 20168 1352
rect 19576 1312 20168 1340
rect 19576 1300 19582 1312
rect 20162 1300 20168 1312
rect 20220 1300 20226 1352
rect 5166 1232 5172 1284
rect 5224 1272 5230 1284
rect 11882 1272 11888 1284
rect 5224 1244 11888 1272
rect 5224 1232 5230 1244
rect 11882 1232 11888 1244
rect 11940 1232 11946 1284
rect 13538 1232 13544 1284
rect 13596 1232 13602 1284
rect 56778 1164 56784 1216
rect 56836 1204 56842 1216
rect 57054 1204 57060 1216
rect 56836 1176 57060 1204
rect 56836 1164 56842 1176
rect 57054 1164 57060 1176
rect 57112 1164 57118 1216
rect 57054 1028 57060 1080
rect 57112 1068 57118 1080
rect 59446 1068 59452 1080
rect 57112 1040 59452 1068
rect 57112 1028 57118 1040
rect 59446 1028 59452 1040
rect 59504 1028 59510 1080
rect 4890 960 4896 1012
rect 4948 1000 4954 1012
rect 4948 972 12434 1000
rect 4948 960 4954 972
rect 9674 892 9680 944
rect 9732 932 9738 944
rect 10870 932 10876 944
rect 9732 904 10876 932
rect 9732 892 9738 904
rect 10870 892 10876 904
rect 10928 892 10934 944
rect 12406 932 12434 972
rect 12894 932 12900 944
rect 12406 904 12900 932
rect 12894 892 12900 904
rect 12952 892 12958 944
rect 2498 144 2504 196
rect 2556 184 2562 196
rect 9674 184 9680 196
rect 2556 156 9680 184
rect 2556 144 2562 156
rect 9674 144 9680 156
rect 9732 144 9738 196
<< via1 >>
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 5172 57400 5224 57452
rect 15200 57443 15252 57452
rect 15200 57409 15209 57443
rect 15209 57409 15243 57443
rect 15243 57409 15252 57443
rect 15200 57400 15252 57409
rect 25044 57400 25096 57452
rect 34980 57400 35032 57452
rect 44916 57400 44968 57452
rect 54852 57400 54904 57452
rect 64788 57400 64840 57452
rect 66996 57443 67048 57452
rect 66996 57409 67005 57443
rect 67005 57409 67039 57443
rect 67039 57409 67048 57443
rect 66996 57400 67048 57409
rect 67548 57400 67600 57452
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 65654 57094 65706 57146
rect 65718 57094 65770 57146
rect 65782 57094 65834 57146
rect 65846 57094 65898 57146
rect 65910 57094 65962 57146
rect 68100 56831 68152 56840
rect 68100 56797 68109 56831
rect 68109 56797 68143 56831
rect 68143 56797 68152 56831
rect 68100 56788 68152 56797
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 65654 56006 65706 56058
rect 65718 56006 65770 56058
rect 65782 56006 65834 56058
rect 65846 56006 65898 56058
rect 65910 56006 65962 56058
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 67640 55131 67692 55140
rect 67640 55097 67649 55131
rect 67649 55097 67683 55131
rect 67683 55097 67692 55131
rect 67640 55088 67692 55097
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 65654 54918 65706 54970
rect 65718 54918 65770 54970
rect 65782 54918 65834 54970
rect 65846 54918 65898 54970
rect 65910 54918 65962 54970
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 67548 53932 67600 53984
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 65654 53830 65706 53882
rect 65718 53830 65770 53882
rect 65782 53830 65834 53882
rect 65846 53830 65898 53882
rect 65910 53830 65962 53882
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 65654 52742 65706 52794
rect 65718 52742 65770 52794
rect 65782 52742 65834 52794
rect 65846 52742 65898 52794
rect 65910 52742 65962 52794
rect 68100 52479 68152 52488
rect 68100 52445 68109 52479
rect 68109 52445 68143 52479
rect 68143 52445 68152 52479
rect 68100 52436 68152 52445
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 65654 51654 65706 51706
rect 65718 51654 65770 51706
rect 65782 51654 65834 51706
rect 65846 51654 65898 51706
rect 65910 51654 65962 51706
rect 68100 51391 68152 51400
rect 68100 51357 68109 51391
rect 68109 51357 68143 51391
rect 68143 51357 68152 51391
rect 68100 51348 68152 51357
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 65654 50566 65706 50618
rect 65718 50566 65770 50618
rect 65782 50566 65834 50618
rect 65846 50566 65898 50618
rect 65910 50566 65962 50618
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 67640 49759 67692 49768
rect 67640 49725 67649 49759
rect 67649 49725 67683 49759
rect 67683 49725 67692 49759
rect 67640 49716 67692 49725
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 65654 49478 65706 49530
rect 65718 49478 65770 49530
rect 65782 49478 65834 49530
rect 65846 49478 65898 49530
rect 65910 49478 65962 49530
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 67640 48535 67692 48544
rect 67640 48501 67649 48535
rect 67649 48501 67683 48535
rect 67683 48501 67692 48535
rect 67640 48492 67692 48501
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 65654 48390 65706 48442
rect 65718 48390 65770 48442
rect 65782 48390 65834 48442
rect 65846 48390 65898 48442
rect 65910 48390 65962 48442
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 65654 47302 65706 47354
rect 65718 47302 65770 47354
rect 65782 47302 65834 47354
rect 65846 47302 65898 47354
rect 65910 47302 65962 47354
rect 68100 47039 68152 47048
rect 68100 47005 68109 47039
rect 68109 47005 68143 47039
rect 68143 47005 68152 47039
rect 68100 46996 68152 47005
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 65654 46214 65706 46266
rect 65718 46214 65770 46266
rect 65782 46214 65834 46266
rect 65846 46214 65898 46266
rect 65910 46214 65962 46266
rect 68100 45951 68152 45960
rect 68100 45917 68109 45951
rect 68109 45917 68143 45951
rect 68143 45917 68152 45951
rect 68100 45908 68152 45917
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 65654 45126 65706 45178
rect 65718 45126 65770 45178
rect 65782 45126 65834 45178
rect 65846 45126 65898 45178
rect 65910 45126 65962 45178
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 67640 44251 67692 44260
rect 67640 44217 67649 44251
rect 67649 44217 67683 44251
rect 67683 44217 67692 44251
rect 67640 44208 67692 44217
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 65654 44038 65706 44090
rect 65718 44038 65770 44090
rect 65782 44038 65834 44090
rect 65846 44038 65898 44090
rect 65910 44038 65962 44090
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 67640 43095 67692 43104
rect 67640 43061 67649 43095
rect 67649 43061 67683 43095
rect 67683 43061 67692 43095
rect 67640 43052 67692 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 65654 42950 65706 43002
rect 65718 42950 65770 43002
rect 65782 42950 65834 43002
rect 65846 42950 65898 43002
rect 65910 42950 65962 43002
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 65654 41862 65706 41914
rect 65718 41862 65770 41914
rect 65782 41862 65834 41914
rect 65846 41862 65898 41914
rect 65910 41862 65962 41914
rect 68100 41599 68152 41608
rect 68100 41565 68109 41599
rect 68109 41565 68143 41599
rect 68143 41565 68152 41599
rect 68100 41556 68152 41565
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 65654 40774 65706 40826
rect 65718 40774 65770 40826
rect 65782 40774 65834 40826
rect 65846 40774 65898 40826
rect 65910 40774 65962 40826
rect 68100 40511 68152 40520
rect 68100 40477 68109 40511
rect 68109 40477 68143 40511
rect 68143 40477 68152 40511
rect 68100 40468 68152 40477
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 65654 39686 65706 39738
rect 65718 39686 65770 39738
rect 65782 39686 65834 39738
rect 65846 39686 65898 39738
rect 65910 39686 65962 39738
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 67640 38811 67692 38820
rect 67640 38777 67649 38811
rect 67649 38777 67683 38811
rect 67683 38777 67692 38811
rect 67640 38768 67692 38777
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 65654 38598 65706 38650
rect 65718 38598 65770 38650
rect 65782 38598 65834 38650
rect 65846 38598 65898 38650
rect 65910 38598 65962 38650
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 67640 37655 67692 37664
rect 67640 37621 67649 37655
rect 67649 37621 67683 37655
rect 67683 37621 67692 37655
rect 67640 37612 67692 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 65654 37510 65706 37562
rect 65718 37510 65770 37562
rect 65782 37510 65834 37562
rect 65846 37510 65898 37562
rect 65910 37510 65962 37562
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 65654 36422 65706 36474
rect 65718 36422 65770 36474
rect 65782 36422 65834 36474
rect 65846 36422 65898 36474
rect 65910 36422 65962 36474
rect 68100 36159 68152 36168
rect 68100 36125 68109 36159
rect 68109 36125 68143 36159
rect 68143 36125 68152 36159
rect 68100 36116 68152 36125
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 65654 35334 65706 35386
rect 65718 35334 65770 35386
rect 65782 35334 65834 35386
rect 65846 35334 65898 35386
rect 65910 35334 65962 35386
rect 68100 35071 68152 35080
rect 68100 35037 68109 35071
rect 68109 35037 68143 35071
rect 68143 35037 68152 35071
rect 68100 35028 68152 35037
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 65654 34246 65706 34298
rect 65718 34246 65770 34298
rect 65782 34246 65834 34298
rect 65846 34246 65898 34298
rect 65910 34246 65962 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 67640 33371 67692 33380
rect 67640 33337 67649 33371
rect 67649 33337 67683 33371
rect 67683 33337 67692 33371
rect 67640 33328 67692 33337
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 65654 33158 65706 33210
rect 65718 33158 65770 33210
rect 65782 33158 65834 33210
rect 65846 33158 65898 33210
rect 65910 33158 65962 33210
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 21364 32172 21416 32224
rect 22468 32172 22520 32224
rect 67640 32215 67692 32224
rect 67640 32181 67649 32215
rect 67649 32181 67683 32215
rect 67683 32181 67692 32215
rect 67640 32172 67692 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 65654 32070 65706 32122
rect 65718 32070 65770 32122
rect 65782 32070 65834 32122
rect 65846 32070 65898 32122
rect 65910 32070 65962 32122
rect 21824 31968 21876 32020
rect 21364 31875 21416 31884
rect 21364 31841 21373 31875
rect 21373 31841 21407 31875
rect 21407 31841 21416 31875
rect 21364 31832 21416 31841
rect 15108 31739 15160 31748
rect 15108 31705 15117 31739
rect 15117 31705 15151 31739
rect 15151 31705 15160 31739
rect 15108 31696 15160 31705
rect 15292 31739 15344 31748
rect 15292 31705 15301 31739
rect 15301 31705 15335 31739
rect 15335 31705 15344 31739
rect 15292 31696 15344 31705
rect 21364 31696 21416 31748
rect 15568 31628 15620 31680
rect 18512 31628 18564 31680
rect 22376 31764 22428 31816
rect 23296 31807 23348 31816
rect 23296 31773 23305 31807
rect 23305 31773 23339 31807
rect 23339 31773 23348 31807
rect 23296 31764 23348 31773
rect 22192 31696 22244 31748
rect 23572 31696 23624 31748
rect 23388 31628 23440 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 12624 31356 12676 31408
rect 3424 31288 3476 31340
rect 12440 31288 12492 31340
rect 15108 31288 15160 31340
rect 15936 31356 15988 31408
rect 4804 31220 4856 31272
rect 15568 31331 15620 31340
rect 15568 31297 15577 31331
rect 15577 31297 15611 31331
rect 15611 31297 15620 31331
rect 15568 31288 15620 31297
rect 15752 31331 15804 31340
rect 15752 31297 15761 31331
rect 15761 31297 15795 31331
rect 15795 31297 15804 31331
rect 17408 31331 17460 31340
rect 15752 31288 15804 31297
rect 17408 31297 17417 31331
rect 17417 31297 17451 31331
rect 17451 31297 17460 31331
rect 17408 31288 17460 31297
rect 17592 31331 17644 31340
rect 17592 31297 17601 31331
rect 17601 31297 17635 31331
rect 17635 31297 17644 31331
rect 17592 31288 17644 31297
rect 18512 31331 18564 31340
rect 18512 31297 18521 31331
rect 18521 31297 18555 31331
rect 18555 31297 18564 31331
rect 18512 31288 18564 31297
rect 19524 31331 19576 31340
rect 2872 31127 2924 31136
rect 2872 31093 2881 31127
rect 2881 31093 2915 31127
rect 2915 31093 2924 31127
rect 15660 31152 15712 31204
rect 19524 31297 19533 31331
rect 19533 31297 19567 31331
rect 19567 31297 19576 31331
rect 19524 31288 19576 31297
rect 22284 31288 22336 31340
rect 22376 31288 22428 31340
rect 23480 31331 23532 31340
rect 23480 31297 23489 31331
rect 23489 31297 23523 31331
rect 23523 31297 23532 31331
rect 23480 31288 23532 31297
rect 20076 31220 20128 31272
rect 23388 31220 23440 31272
rect 2872 31084 2924 31093
rect 13636 31084 13688 31136
rect 15108 31127 15160 31136
rect 15108 31093 15117 31127
rect 15117 31093 15151 31127
rect 15151 31093 15160 31127
rect 15108 31084 15160 31093
rect 15200 31084 15252 31136
rect 17408 31084 17460 31136
rect 18236 31127 18288 31136
rect 18236 31093 18245 31127
rect 18245 31093 18279 31127
rect 18279 31093 18288 31127
rect 18236 31084 18288 31093
rect 19984 31127 20036 31136
rect 19984 31093 19993 31127
rect 19993 31093 20027 31127
rect 20027 31093 20036 31127
rect 19984 31084 20036 31093
rect 22192 31152 22244 31204
rect 25596 31152 25648 31204
rect 24860 31084 24912 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 65654 30982 65706 31034
rect 65718 30982 65770 31034
rect 65782 30982 65834 31034
rect 65846 30982 65898 31034
rect 65910 30982 65962 31034
rect 15292 30880 15344 30932
rect 19524 30880 19576 30932
rect 17408 30744 17460 30796
rect 6736 30719 6788 30728
rect 6736 30685 6745 30719
rect 6745 30685 6779 30719
rect 6779 30685 6788 30719
rect 6736 30676 6788 30685
rect 11060 30676 11112 30728
rect 13820 30676 13872 30728
rect 18236 30676 18288 30728
rect 22468 30719 22520 30728
rect 22468 30685 22486 30719
rect 22486 30685 22520 30719
rect 22468 30676 22520 30685
rect 24032 30676 24084 30728
rect 68100 30719 68152 30728
rect 68100 30685 68109 30719
rect 68109 30685 68143 30719
rect 68143 30685 68152 30719
rect 68100 30676 68152 30685
rect 7104 30608 7156 30660
rect 9220 30608 9272 30660
rect 10968 30608 11020 30660
rect 13176 30608 13228 30660
rect 15108 30608 15160 30660
rect 19432 30651 19484 30660
rect 19432 30617 19441 30651
rect 19441 30617 19475 30651
rect 19475 30617 19484 30651
rect 19432 30608 19484 30617
rect 8116 30583 8168 30592
rect 8116 30549 8125 30583
rect 8125 30549 8159 30583
rect 8159 30549 8168 30583
rect 8116 30540 8168 30549
rect 9772 30540 9824 30592
rect 12624 30540 12676 30592
rect 14096 30540 14148 30592
rect 15752 30540 15804 30592
rect 17408 30540 17460 30592
rect 17592 30540 17644 30592
rect 21364 30583 21416 30592
rect 21364 30549 21373 30583
rect 21373 30549 21407 30583
rect 21407 30549 21416 30583
rect 21364 30540 21416 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 12900 30336 12952 30388
rect 1676 30268 1728 30320
rect 2688 30200 2740 30252
rect 2872 30132 2924 30184
rect 2136 29996 2188 30048
rect 2504 29996 2556 30048
rect 4804 30268 4856 30320
rect 6736 30268 6788 30320
rect 13176 30311 13228 30320
rect 13176 30277 13185 30311
rect 13185 30277 13219 30311
rect 13219 30277 13228 30311
rect 13176 30268 13228 30277
rect 15936 30336 15988 30388
rect 18236 30336 18288 30388
rect 23296 30336 23348 30388
rect 17132 30268 17184 30320
rect 19984 30268 20036 30320
rect 21824 30311 21876 30320
rect 21824 30277 21833 30311
rect 21833 30277 21867 30311
rect 21867 30277 21876 30311
rect 21824 30268 21876 30277
rect 4712 30243 4764 30252
rect 4712 30209 4746 30243
rect 4746 30209 4764 30243
rect 9312 30243 9364 30252
rect 4712 30200 4764 30209
rect 9312 30209 9321 30243
rect 9321 30209 9355 30243
rect 9355 30209 9364 30243
rect 9312 30200 9364 30209
rect 13452 30243 13504 30252
rect 13452 30209 13461 30243
rect 13461 30209 13495 30243
rect 13495 30209 13504 30243
rect 13452 30200 13504 30209
rect 13636 30243 13688 30252
rect 13636 30209 13650 30243
rect 13650 30209 13684 30243
rect 13684 30209 13688 30243
rect 13636 30200 13688 30209
rect 14096 30200 14148 30252
rect 15292 30200 15344 30252
rect 15660 30243 15712 30252
rect 15660 30209 15669 30243
rect 15669 30209 15703 30243
rect 15703 30209 15712 30243
rect 15660 30200 15712 30209
rect 16580 30132 16632 30184
rect 21456 30132 21508 30184
rect 22560 30200 22612 30252
rect 24032 30243 24084 30252
rect 24032 30209 24041 30243
rect 24041 30209 24075 30243
rect 24075 30209 24084 30243
rect 24032 30200 24084 30209
rect 25596 30243 25648 30252
rect 25596 30209 25614 30243
rect 25614 30209 25648 30243
rect 25596 30200 25648 30209
rect 5816 30107 5868 30116
rect 5816 30073 5825 30107
rect 5825 30073 5859 30107
rect 5859 30073 5868 30107
rect 5816 30064 5868 30073
rect 6736 30064 6788 30116
rect 7748 30064 7800 30116
rect 11060 30064 11112 30116
rect 13452 30064 13504 30116
rect 18052 29996 18104 30048
rect 19524 30039 19576 30048
rect 19524 30005 19533 30039
rect 19533 30005 19567 30039
rect 19567 30005 19576 30039
rect 19524 29996 19576 30005
rect 22008 30064 22060 30116
rect 20996 29996 21048 30048
rect 22100 29996 22152 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 65654 29894 65706 29946
rect 65718 29894 65770 29946
rect 65782 29894 65834 29946
rect 65846 29894 65898 29946
rect 65910 29894 65962 29946
rect 3424 29792 3476 29844
rect 10968 29835 11020 29844
rect 10968 29801 10977 29835
rect 10977 29801 11011 29835
rect 11011 29801 11020 29835
rect 10968 29792 11020 29801
rect 1952 29631 2004 29640
rect 1952 29597 1961 29631
rect 1961 29597 1995 29631
rect 1995 29597 2004 29631
rect 1952 29588 2004 29597
rect 2136 29631 2188 29640
rect 2136 29597 2145 29631
rect 2145 29597 2179 29631
rect 2179 29597 2188 29631
rect 2136 29588 2188 29597
rect 2780 29724 2832 29776
rect 9404 29724 9456 29776
rect 13268 29724 13320 29776
rect 12900 29656 12952 29708
rect 7288 29631 7340 29640
rect 7288 29597 7297 29631
rect 7297 29597 7331 29631
rect 7331 29597 7340 29631
rect 7288 29588 7340 29597
rect 2412 29520 2464 29572
rect 2688 29520 2740 29572
rect 5448 29520 5500 29572
rect 7196 29520 7248 29572
rect 11060 29588 11112 29640
rect 12992 29588 13044 29640
rect 13084 29588 13136 29640
rect 13452 29656 13504 29708
rect 17040 29656 17092 29708
rect 13360 29631 13412 29640
rect 13360 29597 13369 29631
rect 13369 29597 13403 29631
rect 13403 29597 13412 29631
rect 13360 29588 13412 29597
rect 14096 29588 14148 29640
rect 14740 29588 14792 29640
rect 4160 29495 4212 29504
rect 4160 29461 4169 29495
rect 4169 29461 4203 29495
rect 4203 29461 4212 29495
rect 4160 29452 4212 29461
rect 6644 29452 6696 29504
rect 7656 29452 7708 29504
rect 9220 29520 9272 29572
rect 10232 29520 10284 29572
rect 12440 29563 12492 29572
rect 12440 29529 12449 29563
rect 12449 29529 12483 29563
rect 12483 29529 12492 29563
rect 12440 29520 12492 29529
rect 17316 29631 17368 29640
rect 17316 29597 17325 29631
rect 17325 29597 17359 29631
rect 17359 29597 17368 29631
rect 17316 29588 17368 29597
rect 17132 29520 17184 29572
rect 19524 29792 19576 29844
rect 22560 29835 22612 29844
rect 22560 29801 22569 29835
rect 22569 29801 22603 29835
rect 22603 29801 22612 29835
rect 22560 29792 22612 29801
rect 18052 29631 18104 29640
rect 18052 29597 18061 29631
rect 18061 29597 18095 29631
rect 18095 29597 18104 29631
rect 18052 29588 18104 29597
rect 18236 29631 18288 29640
rect 18236 29597 18243 29631
rect 18243 29597 18288 29631
rect 18236 29588 18288 29597
rect 18512 29631 18564 29640
rect 18512 29597 18526 29631
rect 18526 29597 18560 29631
rect 18560 29597 18564 29631
rect 18512 29588 18564 29597
rect 19248 29631 19300 29640
rect 19248 29597 19257 29631
rect 19257 29597 19291 29631
rect 19291 29597 19300 29631
rect 19248 29588 19300 29597
rect 21364 29656 21416 29708
rect 19064 29520 19116 29572
rect 19616 29563 19668 29572
rect 19616 29529 19625 29563
rect 19625 29529 19659 29563
rect 19659 29529 19668 29563
rect 22100 29724 22152 29776
rect 22192 29724 22244 29776
rect 19616 29520 19668 29529
rect 9128 29452 9180 29504
rect 12808 29452 12860 29504
rect 16580 29495 16632 29504
rect 16580 29461 16589 29495
rect 16589 29461 16623 29495
rect 16623 29461 16632 29495
rect 16580 29452 16632 29461
rect 18604 29452 18656 29504
rect 19156 29452 19208 29504
rect 19432 29452 19484 29504
rect 20260 29452 20312 29504
rect 22376 29588 22428 29640
rect 26976 29631 27028 29640
rect 26976 29597 26985 29631
rect 26985 29597 27019 29631
rect 27019 29597 27028 29631
rect 26976 29588 27028 29597
rect 68100 29631 68152 29640
rect 68100 29597 68109 29631
rect 68109 29597 68143 29631
rect 68143 29597 68152 29631
rect 68100 29588 68152 29597
rect 26240 29520 26292 29572
rect 23480 29452 23532 29504
rect 25228 29452 25280 29504
rect 25504 29452 25556 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 2412 29248 2464 29300
rect 4712 29248 4764 29300
rect 7104 29291 7156 29300
rect 7104 29257 7113 29291
rect 7113 29257 7147 29291
rect 7147 29257 7156 29291
rect 7104 29248 7156 29257
rect 1952 29112 2004 29164
rect 2504 29112 2556 29164
rect 4804 29180 4856 29232
rect 2596 28976 2648 29028
rect 2688 28976 2740 29028
rect 2780 28976 2832 29028
rect 4620 29112 4672 29164
rect 7196 29180 7248 29232
rect 6644 29155 6696 29164
rect 6644 29121 6653 29155
rect 6653 29121 6687 29155
rect 6687 29121 6696 29155
rect 6644 29112 6696 29121
rect 6828 29155 6880 29164
rect 6828 29121 6837 29155
rect 6837 29121 6871 29155
rect 6871 29121 6880 29155
rect 7748 29155 7800 29164
rect 6828 29112 6880 29121
rect 7748 29121 7757 29155
rect 7757 29121 7791 29155
rect 7791 29121 7800 29155
rect 7748 29112 7800 29121
rect 8024 29155 8076 29164
rect 8024 29121 8058 29155
rect 8058 29121 8076 29155
rect 8024 29112 8076 29121
rect 9496 29112 9548 29164
rect 9772 29155 9824 29164
rect 9772 29121 9781 29155
rect 9781 29121 9815 29155
rect 9815 29121 9824 29155
rect 9772 29112 9824 29121
rect 9956 29248 10008 29300
rect 10232 29291 10284 29300
rect 10232 29257 10241 29291
rect 10241 29257 10275 29291
rect 10275 29257 10284 29291
rect 10232 29248 10284 29257
rect 12992 29248 13044 29300
rect 15200 29248 15252 29300
rect 15936 29291 15988 29300
rect 15936 29257 15945 29291
rect 15945 29257 15979 29291
rect 15979 29257 15988 29291
rect 15936 29248 15988 29257
rect 19248 29248 19300 29300
rect 10048 29112 10100 29164
rect 5448 29019 5500 29028
rect 5448 28985 5457 29019
rect 5457 28985 5491 29019
rect 5491 28985 5500 29019
rect 5448 28976 5500 28985
rect 7380 29044 7432 29096
rect 9312 29044 9364 29096
rect 12532 29180 12584 29232
rect 14464 29180 14516 29232
rect 17224 29223 17276 29232
rect 17224 29189 17233 29223
rect 17233 29189 17267 29223
rect 17267 29189 17276 29223
rect 17224 29180 17276 29189
rect 17500 29180 17552 29232
rect 12808 29112 12860 29164
rect 14648 29112 14700 29164
rect 16304 29112 16356 29164
rect 16580 29112 16632 29164
rect 17132 29155 17184 29164
rect 17132 29121 17141 29155
rect 17141 29121 17175 29155
rect 17175 29121 17184 29155
rect 17408 29155 17460 29164
rect 17132 29112 17184 29121
rect 17408 29121 17417 29155
rect 17417 29121 17451 29155
rect 17451 29121 17460 29155
rect 17408 29112 17460 29121
rect 18604 29112 18656 29164
rect 22008 29180 22060 29232
rect 24032 29180 24084 29232
rect 13820 29044 13872 29096
rect 18880 29044 18932 29096
rect 7012 28976 7064 29028
rect 9128 29019 9180 29028
rect 9128 28985 9137 29019
rect 9137 28985 9171 29019
rect 9171 28985 9180 29019
rect 19432 29155 19484 29164
rect 19432 29121 19446 29155
rect 19446 29121 19480 29155
rect 19480 29121 19484 29155
rect 19432 29112 19484 29121
rect 23848 29112 23900 29164
rect 26976 29180 27028 29232
rect 29092 29155 29144 29164
rect 29092 29121 29101 29155
rect 29101 29121 29135 29155
rect 29135 29121 29144 29155
rect 29092 29112 29144 29121
rect 9128 28976 9180 28985
rect 17960 28951 18012 28960
rect 17960 28917 17969 28951
rect 17969 28917 18003 28951
rect 18003 28917 18012 28951
rect 17960 28908 18012 28917
rect 18512 28908 18564 28960
rect 20168 28976 20220 29028
rect 23756 29019 23808 29028
rect 23756 28985 23765 29019
rect 23765 28985 23799 29019
rect 23799 28985 23808 29019
rect 23756 28976 23808 28985
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 65654 28806 65706 28858
rect 65718 28806 65770 28858
rect 65782 28806 65834 28858
rect 65846 28806 65898 28858
rect 65910 28806 65962 28858
rect 4620 28704 4672 28756
rect 8024 28704 8076 28756
rect 16396 28704 16448 28756
rect 4068 28636 4120 28688
rect 1676 28543 1728 28552
rect 1676 28509 1685 28543
rect 1685 28509 1719 28543
rect 1719 28509 1728 28543
rect 1676 28500 1728 28509
rect 2596 28500 2648 28552
rect 5632 28568 5684 28620
rect 7012 28568 7064 28620
rect 1860 28475 1912 28484
rect 1860 28441 1869 28475
rect 1869 28441 1903 28475
rect 1903 28441 1912 28475
rect 1860 28432 1912 28441
rect 3332 28432 3384 28484
rect 2044 28407 2096 28416
rect 2044 28373 2053 28407
rect 2053 28373 2087 28407
rect 2087 28373 2096 28407
rect 2044 28364 2096 28373
rect 7196 28500 7248 28552
rect 7656 28543 7708 28552
rect 7656 28509 7665 28543
rect 7665 28509 7699 28543
rect 7699 28509 7708 28543
rect 7656 28500 7708 28509
rect 7012 28432 7064 28484
rect 7380 28432 7432 28484
rect 11060 28500 11112 28552
rect 10232 28475 10284 28484
rect 10232 28441 10266 28475
rect 10266 28441 10284 28475
rect 10232 28432 10284 28441
rect 5908 28364 5960 28416
rect 6828 28364 6880 28416
rect 9404 28407 9456 28416
rect 9404 28373 9413 28407
rect 9413 28373 9447 28407
rect 9447 28373 9456 28407
rect 9404 28364 9456 28373
rect 10048 28364 10100 28416
rect 11152 28364 11204 28416
rect 12992 28543 13044 28552
rect 12992 28509 13001 28543
rect 13001 28509 13035 28543
rect 13035 28509 13044 28543
rect 12992 28500 13044 28509
rect 13360 28543 13412 28552
rect 13360 28509 13369 28543
rect 13369 28509 13403 28543
rect 13403 28509 13412 28543
rect 13360 28500 13412 28509
rect 14464 28543 14516 28552
rect 14464 28509 14473 28543
rect 14473 28509 14507 28543
rect 14507 28509 14516 28543
rect 14464 28500 14516 28509
rect 16764 28543 16816 28552
rect 16764 28509 16773 28543
rect 16773 28509 16807 28543
rect 16807 28509 16816 28543
rect 16764 28500 16816 28509
rect 16948 28543 17000 28552
rect 16948 28509 16955 28543
rect 16955 28509 17000 28543
rect 16948 28500 17000 28509
rect 21456 28611 21508 28620
rect 21456 28577 21465 28611
rect 21465 28577 21499 28611
rect 21499 28577 21508 28611
rect 21456 28568 21508 28577
rect 24032 28568 24084 28620
rect 17960 28500 18012 28552
rect 19340 28500 19392 28552
rect 20628 28500 20680 28552
rect 29000 28543 29052 28552
rect 29000 28509 29009 28543
rect 29009 28509 29043 28543
rect 29043 28509 29052 28543
rect 29000 28500 29052 28509
rect 13176 28475 13228 28484
rect 13176 28441 13185 28475
rect 13185 28441 13219 28475
rect 13219 28441 13228 28475
rect 13176 28432 13228 28441
rect 13268 28475 13320 28484
rect 13268 28441 13277 28475
rect 13277 28441 13311 28475
rect 13311 28441 13320 28475
rect 13268 28432 13320 28441
rect 16488 28432 16540 28484
rect 19064 28432 19116 28484
rect 20720 28432 20772 28484
rect 22560 28432 22612 28484
rect 25688 28432 25740 28484
rect 27712 28432 27764 28484
rect 15108 28364 15160 28416
rect 17408 28407 17460 28416
rect 17408 28373 17417 28407
rect 17417 28373 17451 28407
rect 17451 28373 17460 28407
rect 17408 28364 17460 28373
rect 19432 28364 19484 28416
rect 22008 28407 22060 28416
rect 22008 28373 22017 28407
rect 22017 28373 22051 28407
rect 22051 28373 22060 28407
rect 22008 28364 22060 28373
rect 26424 28364 26476 28416
rect 27620 28407 27672 28416
rect 27620 28373 27629 28407
rect 27629 28373 27663 28407
rect 27663 28373 27672 28407
rect 27620 28364 27672 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 1860 28160 1912 28212
rect 6828 28160 6880 28212
rect 10232 28160 10284 28212
rect 16764 28160 16816 28212
rect 20352 28160 20404 28212
rect 20720 28203 20772 28212
rect 20720 28169 20729 28203
rect 20729 28169 20763 28203
rect 20763 28169 20772 28203
rect 20720 28160 20772 28169
rect 22560 28160 22612 28212
rect 25412 28160 25464 28212
rect 26240 28160 26292 28212
rect 2044 28067 2096 28076
rect 2044 28033 2053 28067
rect 2053 28033 2087 28067
rect 2087 28033 2096 28067
rect 2044 28024 2096 28033
rect 2412 28092 2464 28144
rect 3332 28092 3384 28144
rect 5080 28092 5132 28144
rect 3148 28024 3200 28076
rect 7656 28067 7708 28076
rect 7656 28033 7665 28067
rect 7665 28033 7699 28067
rect 7699 28033 7708 28067
rect 7656 28024 7708 28033
rect 9496 28067 9548 28076
rect 9496 28033 9505 28067
rect 9505 28033 9539 28067
rect 9539 28033 9548 28067
rect 9496 28024 9548 28033
rect 9680 28067 9732 28076
rect 9680 28033 9689 28067
rect 9689 28033 9723 28067
rect 9723 28033 9732 28067
rect 9680 28024 9732 28033
rect 12440 28092 12492 28144
rect 13820 28092 13872 28144
rect 15108 28092 15160 28144
rect 2596 27956 2648 28008
rect 7012 27956 7064 28008
rect 7564 27956 7616 28008
rect 12624 28024 12676 28076
rect 9956 27956 10008 28008
rect 13360 28024 13412 28076
rect 13728 28024 13780 28076
rect 15384 28024 15436 28076
rect 16948 28092 17000 28144
rect 18972 28024 19024 28076
rect 19432 28067 19484 28076
rect 19432 28033 19441 28067
rect 19441 28033 19475 28067
rect 19475 28033 19484 28067
rect 19432 28024 19484 28033
rect 20076 28067 20128 28076
rect 13176 27956 13228 28008
rect 19340 27956 19392 28008
rect 20076 28033 20085 28067
rect 20085 28033 20119 28067
rect 20119 28033 20128 28067
rect 20076 28024 20128 28033
rect 20996 28092 21048 28144
rect 22192 28092 22244 28144
rect 21824 28024 21876 28076
rect 29000 28092 29052 28144
rect 30288 28092 30340 28144
rect 21272 27999 21324 28008
rect 21272 27965 21281 27999
rect 21281 27965 21315 27999
rect 21315 27965 21324 27999
rect 22468 28067 22520 28076
rect 22468 28033 22477 28067
rect 22477 28033 22511 28067
rect 22511 28033 22520 28067
rect 22468 28024 22520 28033
rect 25136 28067 25188 28076
rect 21272 27956 21324 27965
rect 22560 27956 22612 28008
rect 13360 27888 13412 27940
rect 20076 27888 20128 27940
rect 20536 27888 20588 27940
rect 25136 28033 25145 28067
rect 25145 28033 25179 28067
rect 25179 28033 25188 28067
rect 25136 28024 25188 28033
rect 25320 27888 25372 27940
rect 2872 27820 2924 27872
rect 7196 27863 7248 27872
rect 7196 27829 7205 27863
rect 7205 27829 7239 27863
rect 7239 27829 7248 27863
rect 7196 27820 7248 27829
rect 13452 27820 13504 27872
rect 14096 27863 14148 27872
rect 14096 27829 14105 27863
rect 14105 27829 14139 27863
rect 14139 27829 14148 27863
rect 14096 27820 14148 27829
rect 14832 27820 14884 27872
rect 15108 27820 15160 27872
rect 16212 27820 16264 27872
rect 16580 27820 16632 27872
rect 17960 27820 18012 27872
rect 19892 27820 19944 27872
rect 21272 27820 21324 27872
rect 22560 27820 22612 27872
rect 23572 27820 23624 27872
rect 24676 27820 24728 27872
rect 29184 28024 29236 28076
rect 67640 27931 67692 27940
rect 67640 27897 67649 27931
rect 67649 27897 67683 27931
rect 67683 27897 67692 27931
rect 67640 27888 67692 27897
rect 26332 27820 26384 27872
rect 29276 27863 29328 27872
rect 29276 27829 29285 27863
rect 29285 27829 29319 27863
rect 29319 27829 29328 27863
rect 29276 27820 29328 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 65654 27718 65706 27770
rect 65718 27718 65770 27770
rect 65782 27718 65834 27770
rect 65846 27718 65898 27770
rect 65910 27718 65962 27770
rect 2872 27616 2924 27668
rect 3332 27480 3384 27532
rect 9680 27616 9732 27668
rect 13452 27616 13504 27668
rect 1676 27412 1728 27464
rect 2320 27412 2372 27464
rect 2596 27412 2648 27464
rect 2136 27344 2188 27396
rect 3056 27387 3108 27396
rect 3056 27353 3065 27387
rect 3065 27353 3099 27387
rect 3099 27353 3108 27387
rect 3056 27344 3108 27353
rect 5080 27412 5132 27464
rect 5448 27455 5500 27464
rect 5448 27421 5457 27455
rect 5457 27421 5491 27455
rect 5491 27421 5500 27455
rect 5448 27412 5500 27421
rect 7748 27480 7800 27532
rect 9496 27480 9548 27532
rect 11060 27523 11112 27532
rect 11060 27489 11069 27523
rect 11069 27489 11103 27523
rect 11103 27489 11112 27523
rect 11060 27480 11112 27489
rect 7472 27455 7524 27464
rect 7472 27421 7481 27455
rect 7481 27421 7515 27455
rect 7515 27421 7524 27455
rect 7472 27412 7524 27421
rect 7564 27415 7576 27440
rect 7576 27415 7610 27440
rect 7610 27415 7616 27440
rect 7564 27388 7616 27415
rect 7656 27455 7708 27464
rect 7656 27421 7665 27455
rect 7665 27421 7699 27455
rect 7699 27421 7708 27455
rect 7656 27412 7708 27421
rect 1676 27276 1728 27328
rect 4436 27319 4488 27328
rect 4436 27285 4445 27319
rect 4445 27285 4479 27319
rect 4479 27285 4488 27319
rect 4436 27276 4488 27285
rect 6828 27319 6880 27328
rect 6828 27285 6837 27319
rect 6837 27285 6871 27319
rect 6871 27285 6880 27319
rect 9220 27344 9272 27396
rect 11152 27412 11204 27464
rect 14096 27412 14148 27464
rect 17040 27616 17092 27668
rect 17684 27616 17736 27668
rect 19892 27616 19944 27668
rect 20996 27616 21048 27668
rect 24676 27616 24728 27668
rect 25688 27659 25740 27668
rect 16304 27523 16356 27532
rect 16304 27489 16313 27523
rect 16313 27489 16347 27523
rect 16347 27489 16356 27523
rect 16304 27480 16356 27489
rect 14556 27455 14608 27464
rect 14556 27421 14565 27455
rect 14565 27421 14599 27455
rect 14599 27421 14608 27455
rect 14556 27412 14608 27421
rect 14740 27455 14792 27464
rect 14740 27421 14749 27455
rect 14749 27421 14783 27455
rect 14783 27421 14792 27455
rect 14740 27412 14792 27421
rect 15016 27412 15068 27464
rect 16488 27412 16540 27464
rect 22008 27548 22060 27600
rect 23848 27591 23900 27600
rect 19340 27523 19392 27532
rect 19340 27489 19349 27523
rect 19349 27489 19383 27523
rect 19383 27489 19392 27523
rect 19340 27480 19392 27489
rect 20352 27480 20404 27532
rect 22192 27480 22244 27532
rect 17224 27455 17276 27464
rect 17224 27421 17238 27455
rect 17238 27421 17272 27455
rect 17272 27421 17276 27455
rect 17224 27412 17276 27421
rect 18144 27412 18196 27464
rect 19064 27412 19116 27464
rect 13268 27344 13320 27396
rect 14648 27344 14700 27396
rect 17040 27387 17092 27396
rect 17040 27353 17049 27387
rect 17049 27353 17083 27387
rect 17083 27353 17092 27387
rect 17040 27344 17092 27353
rect 17132 27387 17184 27396
rect 17132 27353 17141 27387
rect 17141 27353 17175 27387
rect 17175 27353 17184 27387
rect 17132 27344 17184 27353
rect 7932 27319 7984 27328
rect 6828 27276 6880 27285
rect 7932 27285 7941 27319
rect 7941 27285 7975 27319
rect 7975 27285 7984 27319
rect 7932 27276 7984 27285
rect 12624 27276 12676 27328
rect 15936 27276 15988 27328
rect 16028 27276 16080 27328
rect 17776 27276 17828 27328
rect 18052 27344 18104 27396
rect 21824 27412 21876 27464
rect 22468 27523 22520 27532
rect 22468 27489 22477 27523
rect 22477 27489 22511 27523
rect 22511 27489 22520 27523
rect 22468 27480 22520 27489
rect 23204 27455 23256 27464
rect 23204 27421 23213 27455
rect 23213 27421 23247 27455
rect 23247 27421 23256 27455
rect 23204 27412 23256 27421
rect 23848 27557 23857 27591
rect 23857 27557 23891 27591
rect 23891 27557 23900 27591
rect 23848 27548 23900 27557
rect 24860 27548 24912 27600
rect 24952 27480 25004 27532
rect 25412 27548 25464 27600
rect 18604 27319 18656 27328
rect 18604 27285 18613 27319
rect 18613 27285 18647 27319
rect 18647 27285 18656 27319
rect 18604 27276 18656 27285
rect 23572 27455 23624 27464
rect 23572 27421 23581 27455
rect 23581 27421 23615 27455
rect 23615 27421 23624 27455
rect 23572 27412 23624 27421
rect 24216 27412 24268 27464
rect 25136 27412 25188 27464
rect 25688 27625 25697 27659
rect 25697 27625 25731 27659
rect 25731 27625 25740 27659
rect 25688 27616 25740 27625
rect 29184 27548 29236 27600
rect 27436 27480 27488 27532
rect 26056 27412 26108 27464
rect 26792 27412 26844 27464
rect 26148 27387 26200 27396
rect 23480 27276 23532 27328
rect 26148 27353 26157 27387
rect 26157 27353 26191 27387
rect 26191 27353 26200 27387
rect 26148 27344 26200 27353
rect 26424 27344 26476 27396
rect 27528 27344 27580 27396
rect 26884 27276 26936 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 2136 27115 2188 27124
rect 2136 27081 2145 27115
rect 2145 27081 2179 27115
rect 2179 27081 2188 27115
rect 2136 27072 2188 27081
rect 2320 27072 2372 27124
rect 3056 27072 3108 27124
rect 2320 26979 2372 26988
rect 2320 26945 2329 26979
rect 2329 26945 2363 26979
rect 2363 26945 2372 26979
rect 2320 26936 2372 26945
rect 3332 26979 3384 26988
rect 3332 26945 3341 26979
rect 3341 26945 3375 26979
rect 3375 26945 3384 26979
rect 3332 26936 3384 26945
rect 4436 27004 4488 27056
rect 5356 26936 5408 26988
rect 7472 27072 7524 27124
rect 14556 27072 14608 27124
rect 14648 27115 14700 27124
rect 14648 27081 14657 27115
rect 14657 27081 14691 27115
rect 14691 27081 14700 27115
rect 14648 27072 14700 27081
rect 7932 27004 7984 27056
rect 12348 27004 12400 27056
rect 12624 27047 12676 27056
rect 12624 27013 12633 27047
rect 12633 27013 12667 27047
rect 12667 27013 12676 27047
rect 12624 27004 12676 27013
rect 9588 26979 9640 26988
rect 3608 26911 3660 26920
rect 3608 26877 3617 26911
rect 3617 26877 3651 26911
rect 3651 26877 3660 26911
rect 3608 26868 3660 26877
rect 4068 26911 4120 26920
rect 4068 26877 4077 26911
rect 4077 26877 4111 26911
rect 4111 26877 4120 26911
rect 4068 26868 4120 26877
rect 9588 26945 9597 26979
rect 9597 26945 9631 26979
rect 9631 26945 9640 26979
rect 9588 26936 9640 26945
rect 7104 26868 7156 26920
rect 7472 26732 7524 26784
rect 9220 26868 9272 26920
rect 12992 26936 13044 26988
rect 13360 27004 13412 27056
rect 14280 27004 14332 27056
rect 9588 26800 9640 26852
rect 9680 26800 9732 26852
rect 13728 26936 13780 26988
rect 15384 27072 15436 27124
rect 17500 27072 17552 27124
rect 18972 27115 19024 27124
rect 18972 27081 18981 27115
rect 18981 27081 19015 27115
rect 19015 27081 19024 27115
rect 18972 27072 19024 27081
rect 19064 27072 19116 27124
rect 15568 27004 15620 27056
rect 15108 26936 15160 26988
rect 15752 26979 15804 26988
rect 15752 26945 15761 26979
rect 15761 26945 15795 26979
rect 15795 26945 15804 26979
rect 15752 26936 15804 26945
rect 16304 27004 16356 27056
rect 17960 27004 18012 27056
rect 21824 27072 21876 27124
rect 23480 27115 23532 27124
rect 23480 27081 23489 27115
rect 23489 27081 23523 27115
rect 23523 27081 23532 27115
rect 23480 27072 23532 27081
rect 25320 27072 25372 27124
rect 26332 27115 26384 27124
rect 26332 27081 26341 27115
rect 26341 27081 26375 27115
rect 26375 27081 26384 27115
rect 26332 27072 26384 27081
rect 27528 27072 27580 27124
rect 27712 27072 27764 27124
rect 15936 26979 15988 26988
rect 15936 26945 15945 26979
rect 15945 26945 15979 26979
rect 15979 26945 15988 26979
rect 15936 26936 15988 26945
rect 16120 26979 16172 26988
rect 16120 26945 16129 26979
rect 16129 26945 16163 26979
rect 16163 26945 16172 26979
rect 16672 26979 16724 26988
rect 16120 26936 16172 26945
rect 16672 26945 16681 26979
rect 16681 26945 16715 26979
rect 16715 26945 16724 26979
rect 16672 26936 16724 26945
rect 17500 26979 17552 26988
rect 15200 26868 15252 26920
rect 17500 26945 17509 26979
rect 17509 26945 17543 26979
rect 17543 26945 17552 26979
rect 17500 26936 17552 26945
rect 18052 26936 18104 26988
rect 18604 26936 18656 26988
rect 19340 26979 19392 26988
rect 19340 26945 19349 26979
rect 19349 26945 19383 26979
rect 19383 26945 19392 26979
rect 19340 26936 19392 26945
rect 22560 27004 22612 27056
rect 23756 27004 23808 27056
rect 19984 26936 20036 26988
rect 20352 26979 20404 26988
rect 20352 26945 20361 26979
rect 20361 26945 20395 26979
rect 20395 26945 20404 26979
rect 20352 26936 20404 26945
rect 23204 26936 23256 26988
rect 25504 26936 25556 26988
rect 26792 26936 26844 26988
rect 26148 26868 26200 26920
rect 27344 26979 27396 26988
rect 27344 26945 27353 26979
rect 27353 26945 27387 26979
rect 27387 26945 27396 26979
rect 27344 26936 27396 26945
rect 27528 26936 27580 26988
rect 29184 26936 29236 26988
rect 27436 26868 27488 26920
rect 16948 26800 17000 26852
rect 19248 26800 19300 26852
rect 22008 26800 22060 26852
rect 23572 26800 23624 26852
rect 26332 26800 26384 26852
rect 27068 26800 27120 26852
rect 8208 26732 8260 26784
rect 13912 26732 13964 26784
rect 15476 26732 15528 26784
rect 15660 26732 15712 26784
rect 17408 26732 17460 26784
rect 18420 26732 18472 26784
rect 67640 26775 67692 26784
rect 67640 26741 67649 26775
rect 67649 26741 67683 26775
rect 67683 26741 67692 26775
rect 67640 26732 67692 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 65654 26630 65706 26682
rect 65718 26630 65770 26682
rect 65782 26630 65834 26682
rect 65846 26630 65898 26682
rect 65910 26630 65962 26682
rect 5816 26571 5868 26580
rect 5816 26537 5825 26571
rect 5825 26537 5859 26571
rect 5859 26537 5868 26571
rect 5816 26528 5868 26537
rect 9680 26528 9732 26580
rect 14096 26528 14148 26580
rect 15200 26528 15252 26580
rect 15476 26528 15528 26580
rect 16120 26528 16172 26580
rect 27068 26528 27120 26580
rect 2596 26435 2648 26444
rect 2596 26401 2605 26435
rect 2605 26401 2639 26435
rect 2639 26401 2648 26435
rect 2596 26392 2648 26401
rect 7012 26435 7064 26444
rect 7012 26401 7021 26435
rect 7021 26401 7055 26435
rect 7055 26401 7064 26435
rect 7012 26392 7064 26401
rect 7472 26392 7524 26444
rect 9220 26392 9272 26444
rect 13728 26392 13780 26444
rect 14924 26460 14976 26512
rect 16672 26460 16724 26512
rect 17408 26503 17460 26512
rect 17408 26469 17417 26503
rect 17417 26469 17451 26503
rect 17451 26469 17460 26503
rect 17408 26460 17460 26469
rect 20352 26460 20404 26512
rect 3884 26367 3936 26376
rect 3884 26333 3893 26367
rect 3893 26333 3927 26367
rect 3927 26333 3936 26367
rect 3884 26324 3936 26333
rect 4252 26324 4304 26376
rect 5448 26324 5500 26376
rect 7288 26367 7340 26376
rect 7288 26333 7297 26367
rect 7297 26333 7331 26367
rect 7331 26333 7340 26367
rect 7288 26324 7340 26333
rect 7932 26367 7984 26376
rect 7932 26333 7941 26367
rect 7941 26333 7975 26367
rect 7975 26333 7984 26367
rect 7932 26324 7984 26333
rect 3056 26256 3108 26308
rect 8852 26324 8904 26376
rect 11796 26367 11848 26376
rect 11796 26333 11805 26367
rect 11805 26333 11839 26367
rect 11839 26333 11848 26367
rect 11796 26324 11848 26333
rect 13820 26324 13872 26376
rect 14096 26367 14148 26376
rect 14096 26333 14105 26367
rect 14105 26333 14139 26367
rect 14139 26333 14148 26367
rect 14096 26324 14148 26333
rect 14740 26324 14792 26376
rect 15108 26324 15160 26376
rect 15384 26324 15436 26376
rect 7472 26188 7524 26240
rect 8392 26256 8444 26308
rect 9312 26256 9364 26308
rect 12900 26256 12952 26308
rect 12992 26256 13044 26308
rect 14280 26299 14332 26308
rect 14280 26265 14289 26299
rect 14289 26265 14323 26299
rect 14323 26265 14332 26299
rect 14280 26256 14332 26265
rect 14372 26299 14424 26308
rect 14372 26265 14381 26299
rect 14381 26265 14415 26299
rect 14415 26265 14424 26299
rect 14372 26256 14424 26265
rect 15016 26256 15068 26308
rect 15660 26367 15712 26376
rect 15660 26333 15669 26367
rect 15669 26333 15703 26367
rect 15703 26333 15712 26367
rect 19340 26392 19392 26444
rect 30288 26392 30340 26444
rect 15660 26324 15712 26333
rect 17040 26367 17092 26376
rect 17040 26333 17049 26367
rect 17049 26333 17083 26367
rect 17083 26333 17092 26367
rect 17040 26324 17092 26333
rect 17224 26367 17276 26376
rect 17224 26333 17238 26367
rect 17238 26333 17272 26367
rect 17272 26333 17276 26367
rect 17224 26324 17276 26333
rect 8484 26188 8536 26240
rect 10416 26231 10468 26240
rect 10416 26197 10425 26231
rect 10425 26197 10459 26231
rect 10459 26197 10468 26231
rect 10416 26188 10468 26197
rect 13820 26188 13872 26240
rect 14740 26188 14792 26240
rect 14924 26188 14976 26240
rect 15200 26231 15252 26240
rect 15200 26197 15209 26231
rect 15209 26197 15243 26231
rect 15243 26197 15252 26231
rect 15200 26188 15252 26197
rect 15292 26188 15344 26240
rect 17132 26299 17184 26308
rect 17132 26265 17141 26299
rect 17141 26265 17175 26299
rect 17175 26265 17184 26299
rect 17132 26256 17184 26265
rect 16672 26188 16724 26240
rect 17776 26324 17828 26376
rect 18144 26367 18196 26376
rect 18144 26333 18153 26367
rect 18153 26333 18187 26367
rect 18187 26333 18196 26367
rect 18144 26324 18196 26333
rect 19248 26324 19300 26376
rect 20352 26324 20404 26376
rect 22744 26367 22796 26376
rect 22744 26333 22753 26367
rect 22753 26333 22787 26367
rect 22787 26333 22796 26367
rect 22744 26324 22796 26333
rect 26240 26324 26292 26376
rect 22468 26299 22520 26308
rect 22468 26265 22486 26299
rect 22486 26265 22520 26299
rect 22468 26256 22520 26265
rect 23204 26256 23256 26308
rect 23572 26256 23624 26308
rect 18696 26188 18748 26240
rect 19064 26188 19116 26240
rect 23848 26231 23900 26240
rect 23848 26197 23857 26231
rect 23857 26197 23891 26231
rect 23891 26197 23900 26231
rect 23848 26188 23900 26197
rect 24860 26256 24912 26308
rect 25964 26256 26016 26308
rect 27620 26324 27672 26376
rect 26976 26256 27028 26308
rect 27528 26256 27580 26308
rect 30748 26256 30800 26308
rect 31576 26188 31628 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 14096 25984 14148 26036
rect 14464 25984 14516 26036
rect 5816 25916 5868 25968
rect 8392 25916 8444 25968
rect 1676 25848 1728 25900
rect 2964 25848 3016 25900
rect 4252 25891 4304 25900
rect 4252 25857 4261 25891
rect 4261 25857 4295 25891
rect 4295 25857 4304 25891
rect 4252 25848 4304 25857
rect 8300 25848 8352 25900
rect 9404 25916 9456 25968
rect 15200 25916 15252 25968
rect 20628 25984 20680 26036
rect 22468 26027 22520 26036
rect 22468 25993 22477 26027
rect 22477 25993 22511 26027
rect 22511 25993 22520 26027
rect 22468 25984 22520 25993
rect 24860 26027 24912 26036
rect 24860 25993 24869 26027
rect 24869 25993 24903 26027
rect 24903 25993 24912 26027
rect 24860 25984 24912 25993
rect 26056 25984 26108 26036
rect 20352 25916 20404 25968
rect 9036 25848 9088 25900
rect 11796 25891 11848 25900
rect 11796 25857 11805 25891
rect 11805 25857 11839 25891
rect 11839 25857 11848 25891
rect 11796 25848 11848 25857
rect 14648 25891 14700 25900
rect 14648 25857 14657 25891
rect 14657 25857 14691 25891
rect 14691 25857 14700 25891
rect 14648 25848 14700 25857
rect 15568 25891 15620 25900
rect 15568 25857 15577 25891
rect 15577 25857 15611 25891
rect 15611 25857 15620 25891
rect 15568 25848 15620 25857
rect 17040 25848 17092 25900
rect 17316 25848 17368 25900
rect 18144 25848 18196 25900
rect 18696 25891 18748 25900
rect 18696 25857 18705 25891
rect 18705 25857 18739 25891
rect 18739 25857 18748 25891
rect 18696 25848 18748 25857
rect 18880 25891 18932 25900
rect 18880 25857 18889 25891
rect 18889 25857 18923 25891
rect 18923 25857 18932 25891
rect 18880 25848 18932 25857
rect 20536 25848 20588 25900
rect 22008 25891 22060 25900
rect 22008 25857 22017 25891
rect 22017 25857 22051 25891
rect 22051 25857 22060 25891
rect 22008 25848 22060 25857
rect 23848 25916 23900 25968
rect 30288 25984 30340 26036
rect 30748 26027 30800 26036
rect 30748 25993 30757 26027
rect 30757 25993 30791 26027
rect 30791 25993 30800 26027
rect 30748 25984 30800 25993
rect 22192 25891 22244 25900
rect 22192 25857 22201 25891
rect 22201 25857 22235 25891
rect 22235 25857 22244 25891
rect 22192 25848 22244 25857
rect 24216 25891 24268 25900
rect 24216 25857 24225 25891
rect 24225 25857 24259 25891
rect 24259 25857 24268 25891
rect 24216 25848 24268 25857
rect 14096 25780 14148 25832
rect 14924 25780 14976 25832
rect 16672 25823 16724 25832
rect 16672 25789 16681 25823
rect 16681 25789 16715 25823
rect 16715 25789 16724 25823
rect 16672 25780 16724 25789
rect 23756 25780 23808 25832
rect 24584 25891 24636 25900
rect 24584 25857 24613 25891
rect 24613 25857 24636 25891
rect 24584 25848 24636 25857
rect 25412 25848 25464 25900
rect 26792 25848 26844 25900
rect 27252 25891 27304 25900
rect 27252 25857 27261 25891
rect 27261 25857 27295 25891
rect 27295 25857 27304 25891
rect 27252 25848 27304 25857
rect 24952 25780 25004 25832
rect 27528 25848 27580 25900
rect 31576 25916 31628 25968
rect 30104 25891 30156 25900
rect 30104 25857 30113 25891
rect 30113 25857 30147 25891
rect 30147 25857 30156 25891
rect 30104 25848 30156 25857
rect 30288 25891 30340 25900
rect 30288 25857 30297 25891
rect 30297 25857 30331 25891
rect 30331 25857 30340 25891
rect 30288 25848 30340 25857
rect 2412 25644 2464 25696
rect 2872 25687 2924 25696
rect 2872 25653 2881 25687
rect 2881 25653 2915 25687
rect 2915 25653 2924 25687
rect 2872 25644 2924 25653
rect 9128 25644 9180 25696
rect 17132 25712 17184 25764
rect 27436 25712 27488 25764
rect 29828 25712 29880 25764
rect 30564 25848 30616 25900
rect 31024 25848 31076 25900
rect 13176 25644 13228 25696
rect 14740 25644 14792 25696
rect 19708 25644 19760 25696
rect 21732 25644 21784 25696
rect 23664 25687 23716 25696
rect 23664 25653 23673 25687
rect 23673 25653 23707 25687
rect 23707 25653 23716 25687
rect 23664 25644 23716 25653
rect 24584 25644 24636 25696
rect 26884 25644 26936 25696
rect 27160 25644 27212 25696
rect 30288 25644 30340 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 65654 25542 65706 25594
rect 65718 25542 65770 25594
rect 65782 25542 65834 25594
rect 65846 25542 65898 25594
rect 65910 25542 65962 25594
rect 2964 25483 3016 25492
rect 2964 25449 2973 25483
rect 2973 25449 3007 25483
rect 3007 25449 3016 25483
rect 2964 25440 3016 25449
rect 2872 25372 2924 25424
rect 7932 25440 7984 25492
rect 9036 25440 9088 25492
rect 12900 25483 12952 25492
rect 12900 25449 12909 25483
rect 12909 25449 12943 25483
rect 12943 25449 12952 25483
rect 12900 25440 12952 25449
rect 14372 25372 14424 25424
rect 2320 25279 2372 25288
rect 2320 25245 2329 25279
rect 2329 25245 2363 25279
rect 2363 25245 2372 25279
rect 2320 25236 2372 25245
rect 1676 25100 1728 25152
rect 2504 25100 2556 25152
rect 5448 25236 5500 25288
rect 8300 25304 8352 25356
rect 14096 25347 14148 25356
rect 14096 25313 14105 25347
rect 14105 25313 14139 25347
rect 14139 25313 14148 25347
rect 14096 25304 14148 25313
rect 7012 25168 7064 25220
rect 7564 25236 7616 25288
rect 7748 25279 7800 25288
rect 7748 25245 7757 25279
rect 7757 25245 7791 25279
rect 7791 25245 7800 25279
rect 7748 25236 7800 25245
rect 7912 25279 7964 25288
rect 7912 25245 7920 25279
rect 7920 25245 7954 25279
rect 7954 25245 7964 25279
rect 7912 25236 7964 25245
rect 8011 25276 8063 25285
rect 8011 25242 8020 25276
rect 8020 25242 8054 25276
rect 8054 25242 8063 25276
rect 8011 25233 8063 25242
rect 8208 25236 8260 25288
rect 8852 25236 8904 25288
rect 9128 25279 9180 25288
rect 9128 25245 9137 25279
rect 9137 25245 9171 25279
rect 9171 25245 9180 25279
rect 9128 25236 9180 25245
rect 13176 25279 13228 25288
rect 13176 25245 13199 25279
rect 13199 25245 13228 25279
rect 13176 25236 13228 25245
rect 8484 25168 8536 25220
rect 12992 25168 13044 25220
rect 13360 25279 13412 25288
rect 13360 25245 13374 25279
rect 13374 25245 13408 25279
rect 13408 25245 13412 25279
rect 13360 25236 13412 25245
rect 13912 25236 13964 25288
rect 14372 25279 14424 25288
rect 14372 25245 14381 25279
rect 14381 25245 14415 25279
rect 14415 25245 14424 25279
rect 14372 25236 14424 25245
rect 16948 25236 17000 25288
rect 18880 25440 18932 25492
rect 27252 25440 27304 25492
rect 27528 25440 27580 25492
rect 30564 25440 30616 25492
rect 19248 25372 19300 25424
rect 17224 25304 17276 25356
rect 17316 25279 17368 25288
rect 17316 25245 17325 25279
rect 17325 25245 17359 25279
rect 17359 25245 17368 25279
rect 17316 25236 17368 25245
rect 17776 25304 17828 25356
rect 18604 25279 18656 25288
rect 18604 25245 18613 25279
rect 18613 25245 18647 25279
rect 18647 25245 18656 25279
rect 18604 25236 18656 25245
rect 19432 25236 19484 25288
rect 20536 25372 20588 25424
rect 26884 25372 26936 25424
rect 19708 25279 19760 25288
rect 19708 25245 19717 25279
rect 19717 25245 19751 25279
rect 19751 25245 19760 25279
rect 19708 25236 19760 25245
rect 20352 25304 20404 25356
rect 20536 25236 20588 25288
rect 22744 25236 22796 25288
rect 15016 25168 15068 25220
rect 17408 25211 17460 25220
rect 17408 25177 17417 25211
rect 17417 25177 17451 25211
rect 17451 25177 17460 25211
rect 17408 25168 17460 25177
rect 23480 25168 23532 25220
rect 26148 25168 26200 25220
rect 26700 25236 26752 25288
rect 27160 25279 27212 25288
rect 27160 25245 27169 25279
rect 27169 25245 27203 25279
rect 27203 25245 27212 25279
rect 27160 25236 27212 25245
rect 29460 25236 29512 25288
rect 30104 25236 30156 25288
rect 26976 25211 27028 25220
rect 26976 25177 26985 25211
rect 26985 25177 27019 25211
rect 27019 25177 27028 25211
rect 26976 25168 27028 25177
rect 33968 25236 34020 25288
rect 68100 25279 68152 25288
rect 68100 25245 68109 25279
rect 68109 25245 68143 25279
rect 68143 25245 68152 25279
rect 68100 25236 68152 25245
rect 31392 25168 31444 25220
rect 7932 25100 7984 25152
rect 9864 25143 9916 25152
rect 9864 25109 9873 25143
rect 9873 25109 9907 25143
rect 9907 25109 9916 25143
rect 9864 25100 9916 25109
rect 15384 25100 15436 25152
rect 15936 25143 15988 25152
rect 15936 25109 15945 25143
rect 15945 25109 15979 25143
rect 15979 25109 15988 25143
rect 15936 25100 15988 25109
rect 17684 25143 17736 25152
rect 17684 25109 17693 25143
rect 17693 25109 17727 25143
rect 17727 25109 17736 25143
rect 17684 25100 17736 25109
rect 23296 25100 23348 25152
rect 25688 25100 25740 25152
rect 26332 25143 26384 25152
rect 26332 25109 26341 25143
rect 26341 25109 26375 25143
rect 26375 25109 26384 25143
rect 26332 25100 26384 25109
rect 31116 25100 31168 25152
rect 31668 25100 31720 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 7564 24896 7616 24948
rect 8208 24896 8260 24948
rect 9864 24896 9916 24948
rect 12624 24939 12676 24948
rect 12624 24905 12633 24939
rect 12633 24905 12667 24939
rect 12667 24905 12676 24939
rect 12624 24896 12676 24905
rect 15936 24896 15988 24948
rect 16120 24896 16172 24948
rect 22192 24896 22244 24948
rect 23480 24939 23532 24948
rect 23480 24905 23489 24939
rect 23489 24905 23523 24939
rect 23523 24905 23532 24939
rect 23480 24896 23532 24905
rect 26056 24896 26108 24948
rect 31116 24939 31168 24948
rect 31116 24905 31125 24939
rect 31125 24905 31159 24939
rect 31159 24905 31168 24939
rect 31116 24896 31168 24905
rect 1676 24828 1728 24880
rect 3240 24828 3292 24880
rect 2412 24803 2464 24812
rect 2412 24769 2421 24803
rect 2421 24769 2455 24803
rect 2455 24769 2464 24803
rect 2412 24760 2464 24769
rect 2504 24803 2556 24812
rect 2504 24769 2513 24803
rect 2513 24769 2547 24803
rect 2547 24769 2556 24803
rect 2504 24760 2556 24769
rect 3700 24760 3752 24812
rect 5448 24828 5500 24880
rect 5540 24828 5592 24880
rect 4068 24803 4120 24812
rect 4068 24769 4102 24803
rect 4102 24769 4120 24803
rect 4068 24760 4120 24769
rect 7748 24760 7800 24812
rect 8484 24803 8536 24812
rect 8484 24769 8493 24803
rect 8493 24769 8527 24803
rect 8527 24769 8536 24803
rect 8484 24760 8536 24769
rect 8668 24803 8720 24812
rect 8668 24769 8677 24803
rect 8677 24769 8711 24803
rect 8711 24769 8720 24803
rect 8668 24760 8720 24769
rect 2320 24692 2372 24744
rect 3056 24692 3108 24744
rect 6276 24692 6328 24744
rect 8024 24692 8076 24744
rect 8576 24692 8628 24744
rect 10416 24760 10468 24812
rect 12072 24803 12124 24812
rect 12072 24769 12081 24803
rect 12081 24769 12115 24803
rect 12115 24769 12124 24803
rect 12072 24760 12124 24769
rect 9404 24692 9456 24744
rect 13176 24828 13228 24880
rect 16028 24828 16080 24880
rect 16212 24828 16264 24880
rect 18604 24828 18656 24880
rect 13728 24760 13780 24812
rect 14372 24760 14424 24812
rect 15476 24760 15528 24812
rect 19708 24803 19760 24812
rect 19708 24769 19726 24803
rect 19726 24769 19760 24803
rect 19708 24760 19760 24769
rect 20628 24760 20680 24812
rect 22284 24760 22336 24812
rect 23756 24803 23808 24812
rect 23756 24769 23765 24803
rect 23765 24769 23799 24803
rect 23799 24769 23808 24803
rect 23756 24760 23808 24769
rect 14280 24692 14332 24744
rect 23664 24692 23716 24744
rect 23940 24803 23992 24812
rect 23940 24769 23954 24803
rect 23954 24769 23988 24803
rect 23988 24769 23992 24803
rect 23940 24760 23992 24769
rect 24216 24760 24268 24812
rect 24584 24760 24636 24812
rect 24860 24760 24912 24812
rect 25412 24760 25464 24812
rect 25688 24760 25740 24812
rect 26332 24828 26384 24880
rect 29000 24760 29052 24812
rect 29828 24828 29880 24880
rect 29460 24803 29512 24812
rect 29460 24769 29469 24803
rect 29469 24769 29503 24803
rect 29503 24769 29512 24803
rect 29460 24760 29512 24769
rect 30012 24760 30064 24812
rect 31024 24828 31076 24880
rect 31668 24760 31720 24812
rect 10968 24599 11020 24608
rect 10968 24565 10977 24599
rect 10977 24565 11011 24599
rect 11011 24565 11020 24599
rect 14740 24599 14792 24608
rect 10968 24556 11020 24565
rect 14740 24565 14749 24599
rect 14749 24565 14783 24599
rect 14783 24565 14792 24599
rect 14740 24556 14792 24565
rect 26056 24624 26108 24676
rect 17040 24556 17092 24608
rect 18236 24556 18288 24608
rect 20536 24599 20588 24608
rect 20536 24565 20545 24599
rect 20545 24565 20579 24599
rect 20579 24565 20588 24599
rect 20536 24556 20588 24565
rect 21824 24599 21876 24608
rect 21824 24565 21833 24599
rect 21833 24565 21867 24599
rect 21867 24565 21876 24599
rect 21824 24556 21876 24565
rect 26148 24556 26200 24608
rect 26608 24556 26660 24608
rect 27068 24556 27120 24608
rect 28816 24599 28868 24608
rect 28816 24565 28825 24599
rect 28825 24565 28859 24599
rect 28859 24565 28868 24599
rect 28816 24556 28868 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 65654 24454 65706 24506
rect 65718 24454 65770 24506
rect 65782 24454 65834 24506
rect 65846 24454 65898 24506
rect 65910 24454 65962 24506
rect 3700 24352 3752 24404
rect 7012 24395 7064 24404
rect 7012 24361 7021 24395
rect 7021 24361 7055 24395
rect 7055 24361 7064 24395
rect 7012 24352 7064 24361
rect 7104 24352 7156 24404
rect 8116 24352 8168 24404
rect 8852 24352 8904 24404
rect 9036 24352 9088 24404
rect 10968 24352 11020 24404
rect 13360 24352 13412 24404
rect 2504 24284 2556 24336
rect 3332 24284 3384 24336
rect 7380 24284 7432 24336
rect 3608 24216 3660 24268
rect 3976 24216 4028 24268
rect 1676 24080 1728 24132
rect 5172 24148 5224 24200
rect 1952 24055 2004 24064
rect 1952 24021 1961 24055
rect 1961 24021 1995 24055
rect 1995 24021 2004 24055
rect 1952 24012 2004 24021
rect 2780 24012 2832 24064
rect 3884 24080 3936 24132
rect 6276 24123 6328 24132
rect 6276 24089 6285 24123
rect 6285 24089 6319 24123
rect 6319 24089 6328 24123
rect 6276 24080 6328 24089
rect 7012 24080 7064 24132
rect 7472 24191 7524 24200
rect 7472 24157 7486 24191
rect 7486 24157 7520 24191
rect 7520 24157 7524 24191
rect 7472 24148 7524 24157
rect 7748 24148 7800 24200
rect 8116 24191 8168 24200
rect 8116 24157 8125 24191
rect 8125 24157 8159 24191
rect 8159 24157 8168 24191
rect 8116 24148 8168 24157
rect 9404 24191 9456 24200
rect 9404 24157 9413 24191
rect 9413 24157 9447 24191
rect 9447 24157 9456 24191
rect 9404 24148 9456 24157
rect 10692 24148 10744 24200
rect 8852 24080 8904 24132
rect 5724 24055 5776 24064
rect 5724 24021 5733 24055
rect 5733 24021 5767 24055
rect 5767 24021 5776 24055
rect 5724 24012 5776 24021
rect 7196 24012 7248 24064
rect 7656 24012 7708 24064
rect 9312 24012 9364 24064
rect 15568 24284 15620 24336
rect 19708 24352 19760 24404
rect 23940 24352 23992 24404
rect 26240 24352 26292 24404
rect 26976 24352 27028 24404
rect 27344 24352 27396 24404
rect 12624 24216 12676 24268
rect 12072 24148 12124 24200
rect 14280 24191 14332 24200
rect 14280 24157 14289 24191
rect 14289 24157 14323 24191
rect 14323 24157 14332 24191
rect 14280 24148 14332 24157
rect 15108 24148 15160 24200
rect 13820 24080 13872 24132
rect 17224 24284 17276 24336
rect 22284 24284 22336 24336
rect 26148 24284 26200 24336
rect 27436 24284 27488 24336
rect 18328 24216 18380 24268
rect 17040 24191 17092 24200
rect 17040 24157 17049 24191
rect 17049 24157 17083 24191
rect 17083 24157 17092 24191
rect 17040 24148 17092 24157
rect 17132 24191 17184 24200
rect 17132 24157 17146 24191
rect 17146 24157 17180 24191
rect 17180 24157 17184 24191
rect 17132 24148 17184 24157
rect 17592 24148 17644 24200
rect 18236 24191 18288 24200
rect 18236 24157 18245 24191
rect 18245 24157 18279 24191
rect 18279 24157 18288 24191
rect 18236 24148 18288 24157
rect 19340 24148 19392 24200
rect 17408 24080 17460 24132
rect 17500 24080 17552 24132
rect 12532 24012 12584 24064
rect 13360 24012 13412 24064
rect 16580 24012 16632 24064
rect 17776 24012 17828 24064
rect 18144 24080 18196 24132
rect 19984 24148 20036 24200
rect 20352 24080 20404 24132
rect 22376 24148 22428 24200
rect 23296 24148 23348 24200
rect 27804 24148 27856 24200
rect 21916 24080 21968 24132
rect 21824 24012 21876 24064
rect 23204 24080 23256 24132
rect 23756 24080 23808 24132
rect 24860 24012 24912 24064
rect 27252 24080 27304 24132
rect 29000 24148 29052 24200
rect 29460 24148 29512 24200
rect 31392 24191 31444 24200
rect 31392 24157 31401 24191
rect 31401 24157 31435 24191
rect 31435 24157 31444 24191
rect 31392 24148 31444 24157
rect 33968 24191 34020 24200
rect 33968 24157 33977 24191
rect 33977 24157 34011 24191
rect 34011 24157 34020 24191
rect 33968 24148 34020 24157
rect 68100 24191 68152 24200
rect 68100 24157 68109 24191
rect 68109 24157 68143 24191
rect 68143 24157 68152 24191
rect 68100 24148 68152 24157
rect 28356 24055 28408 24064
rect 28356 24021 28365 24055
rect 28365 24021 28399 24055
rect 28399 24021 28408 24055
rect 28356 24012 28408 24021
rect 31208 24012 31260 24064
rect 32588 24055 32640 24064
rect 32588 24021 32597 24055
rect 32597 24021 32631 24055
rect 32631 24021 32640 24055
rect 32588 24012 32640 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 4068 23808 4120 23860
rect 5356 23808 5408 23860
rect 3240 23715 3292 23724
rect 3240 23681 3249 23715
rect 3249 23681 3283 23715
rect 3283 23681 3292 23715
rect 3240 23672 3292 23681
rect 3332 23715 3384 23724
rect 3332 23681 3341 23715
rect 3341 23681 3375 23715
rect 3375 23681 3384 23715
rect 3332 23672 3384 23681
rect 5540 23740 5592 23792
rect 5724 23672 5776 23724
rect 6828 23740 6880 23792
rect 7932 23740 7984 23792
rect 8576 23808 8628 23860
rect 8852 23851 8904 23860
rect 8852 23817 8861 23851
rect 8861 23817 8895 23851
rect 8895 23817 8904 23851
rect 8852 23808 8904 23817
rect 9864 23808 9916 23860
rect 12900 23808 12952 23860
rect 15016 23808 15068 23860
rect 15476 23851 15528 23860
rect 15476 23817 15485 23851
rect 15485 23817 15519 23851
rect 15519 23817 15528 23851
rect 15476 23808 15528 23817
rect 15568 23808 15620 23860
rect 6920 23715 6972 23724
rect 6920 23681 6929 23715
rect 6929 23681 6963 23715
rect 6963 23681 6972 23715
rect 6920 23672 6972 23681
rect 7288 23672 7340 23724
rect 7380 23672 7432 23724
rect 2320 23647 2372 23656
rect 2320 23613 2329 23647
rect 2329 23613 2363 23647
rect 2363 23613 2372 23647
rect 2320 23604 2372 23613
rect 2780 23604 2832 23656
rect 6460 23604 6512 23656
rect 8024 23604 8076 23656
rect 8300 23672 8352 23724
rect 3700 23536 3752 23588
rect 7012 23536 7064 23588
rect 3884 23468 3936 23520
rect 7932 23468 7984 23520
rect 13360 23740 13412 23792
rect 18604 23808 18656 23860
rect 20444 23808 20496 23860
rect 27804 23808 27856 23860
rect 12532 23672 12584 23724
rect 12992 23672 13044 23724
rect 13544 23715 13596 23724
rect 13544 23681 13553 23715
rect 13553 23681 13587 23715
rect 13587 23681 13596 23715
rect 13544 23672 13596 23681
rect 13912 23715 13964 23724
rect 13912 23681 13921 23715
rect 13921 23681 13955 23715
rect 13955 23681 13964 23715
rect 13912 23672 13964 23681
rect 15016 23715 15068 23724
rect 15016 23681 15025 23715
rect 15025 23681 15059 23715
rect 15059 23681 15068 23715
rect 15016 23672 15068 23681
rect 18328 23740 18380 23792
rect 21916 23740 21968 23792
rect 25596 23740 25648 23792
rect 27252 23740 27304 23792
rect 29092 23808 29144 23860
rect 29276 23808 29328 23860
rect 31208 23808 31260 23860
rect 28816 23783 28868 23792
rect 28816 23749 28850 23783
rect 28850 23749 28868 23783
rect 28816 23740 28868 23749
rect 15660 23672 15712 23724
rect 17316 23715 17368 23724
rect 17316 23681 17323 23715
rect 17323 23681 17368 23715
rect 17316 23672 17368 23681
rect 17408 23715 17460 23724
rect 17408 23681 17417 23715
rect 17417 23681 17451 23715
rect 17451 23681 17460 23715
rect 17408 23672 17460 23681
rect 17592 23715 17644 23724
rect 17592 23681 17606 23715
rect 17606 23681 17640 23715
rect 17640 23681 17644 23715
rect 17592 23672 17644 23681
rect 18144 23672 18196 23724
rect 16212 23604 16264 23656
rect 19340 23604 19392 23656
rect 19616 23647 19668 23656
rect 19616 23613 19625 23647
rect 19625 23613 19659 23647
rect 19659 23613 19668 23647
rect 19616 23604 19668 23613
rect 17500 23536 17552 23588
rect 19248 23536 19300 23588
rect 21824 23672 21876 23724
rect 23112 23672 23164 23724
rect 24584 23715 24636 23724
rect 24584 23681 24593 23715
rect 24593 23681 24627 23715
rect 24627 23681 24636 23715
rect 24584 23672 24636 23681
rect 26884 23672 26936 23724
rect 31024 23672 31076 23724
rect 31300 23672 31352 23724
rect 32588 23672 32640 23724
rect 23664 23604 23716 23656
rect 24952 23604 25004 23656
rect 13268 23511 13320 23520
rect 13268 23477 13277 23511
rect 13277 23477 13311 23511
rect 13311 23477 13320 23511
rect 13268 23468 13320 23477
rect 17224 23468 17276 23520
rect 22744 23536 22796 23588
rect 26148 23604 26200 23656
rect 26976 23536 27028 23588
rect 22100 23468 22152 23520
rect 25412 23468 25464 23520
rect 26332 23468 26384 23520
rect 30012 23468 30064 23520
rect 30656 23468 30708 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 65654 23366 65706 23418
rect 65718 23366 65770 23418
rect 65782 23366 65834 23418
rect 65846 23366 65898 23418
rect 65910 23366 65962 23418
rect 2412 23264 2464 23316
rect 2596 23264 2648 23316
rect 6920 23264 6972 23316
rect 8300 23264 8352 23316
rect 8668 23264 8720 23316
rect 12992 23307 13044 23316
rect 12992 23273 13001 23307
rect 13001 23273 13035 23307
rect 13035 23273 13044 23307
rect 12992 23264 13044 23273
rect 15016 23264 15068 23316
rect 15660 23307 15712 23316
rect 15660 23273 15669 23307
rect 15669 23273 15703 23307
rect 15703 23273 15712 23307
rect 15660 23264 15712 23273
rect 15752 23264 15804 23316
rect 21916 23307 21968 23316
rect 5632 23239 5684 23248
rect 5632 23205 5641 23239
rect 5641 23205 5675 23239
rect 5675 23205 5684 23239
rect 5632 23196 5684 23205
rect 13544 23239 13596 23248
rect 13544 23205 13553 23239
rect 13553 23205 13587 23239
rect 13587 23205 13596 23239
rect 13544 23196 13596 23205
rect 17500 23196 17552 23248
rect 17592 23196 17644 23248
rect 21916 23273 21925 23307
rect 21925 23273 21959 23307
rect 21959 23273 21968 23307
rect 21916 23264 21968 23273
rect 25596 23307 25648 23316
rect 25596 23273 25605 23307
rect 25605 23273 25639 23307
rect 25639 23273 25648 23307
rect 25596 23264 25648 23273
rect 1952 23128 2004 23180
rect 1860 23103 1912 23112
rect 1860 23069 1869 23103
rect 1869 23069 1903 23103
rect 1903 23069 1912 23103
rect 1860 23060 1912 23069
rect 2320 23103 2372 23112
rect 2320 23069 2329 23103
rect 2329 23069 2363 23103
rect 2363 23069 2372 23103
rect 2320 23060 2372 23069
rect 3332 23128 3384 23180
rect 2044 22992 2096 23044
rect 2872 23060 2924 23112
rect 6368 23060 6420 23112
rect 7288 23060 7340 23112
rect 9312 23128 9364 23180
rect 9404 23128 9456 23180
rect 14280 23128 14332 23180
rect 8944 23103 8996 23112
rect 8944 23069 8953 23103
rect 8953 23069 8987 23103
rect 8987 23069 8996 23103
rect 8944 23060 8996 23069
rect 9036 23060 9088 23112
rect 12440 23060 12492 23112
rect 13820 23060 13872 23112
rect 6092 22992 6144 23044
rect 3056 22924 3108 22976
rect 3884 22924 3936 22976
rect 5172 22967 5224 22976
rect 5172 22933 5181 22967
rect 5181 22933 5215 22967
rect 5215 22933 5224 22967
rect 5172 22924 5224 22933
rect 9036 22924 9088 22976
rect 9496 22992 9548 23044
rect 13268 22992 13320 23044
rect 13912 22992 13964 23044
rect 14740 23060 14792 23112
rect 19340 23128 19392 23180
rect 17592 23103 17644 23112
rect 17592 23069 17601 23103
rect 17601 23069 17635 23103
rect 17635 23069 17644 23103
rect 17592 23060 17644 23069
rect 19432 23103 19484 23112
rect 19432 23069 19441 23103
rect 19441 23069 19475 23103
rect 19475 23069 19484 23103
rect 19432 23060 19484 23069
rect 19616 23103 19668 23112
rect 19616 23069 19625 23103
rect 19625 23069 19659 23103
rect 19659 23069 19668 23103
rect 19616 23060 19668 23069
rect 20352 23128 20404 23180
rect 14924 22992 14976 23044
rect 15384 23035 15436 23044
rect 15384 23001 15393 23035
rect 15393 23001 15427 23035
rect 15427 23001 15436 23035
rect 15384 22992 15436 23001
rect 16028 22992 16080 23044
rect 17040 22992 17092 23044
rect 20076 23060 20128 23112
rect 20628 23060 20680 23112
rect 22652 23103 22704 23112
rect 22652 23069 22661 23103
rect 22661 23069 22695 23103
rect 22695 23069 22704 23103
rect 22652 23060 22704 23069
rect 22836 23103 22888 23112
rect 22836 23069 22845 23103
rect 22845 23069 22879 23103
rect 22879 23069 22888 23103
rect 22836 23060 22888 23069
rect 23756 23196 23808 23248
rect 26976 23171 27028 23180
rect 26976 23137 26985 23171
rect 26985 23137 27019 23171
rect 27019 23137 27028 23171
rect 26976 23128 27028 23137
rect 29828 23171 29880 23180
rect 29828 23137 29837 23171
rect 29837 23137 29871 23171
rect 29871 23137 29880 23171
rect 29828 23128 29880 23137
rect 30472 23128 30524 23180
rect 31392 23128 31444 23180
rect 15016 22924 15068 22976
rect 15108 22924 15160 22976
rect 15844 22924 15896 22976
rect 28356 23060 28408 23112
rect 28908 23060 28960 23112
rect 29920 23060 29972 23112
rect 30932 23060 30984 23112
rect 23112 22992 23164 23044
rect 28080 22992 28132 23044
rect 31116 22992 31168 23044
rect 23296 22967 23348 22976
rect 23296 22933 23305 22967
rect 23305 22933 23339 22967
rect 23339 22933 23348 22967
rect 23296 22924 23348 22933
rect 23756 22967 23808 22976
rect 23756 22933 23765 22967
rect 23765 22933 23799 22967
rect 23799 22933 23808 22967
rect 23756 22924 23808 22933
rect 29000 22967 29052 22976
rect 29000 22933 29009 22967
rect 29009 22933 29043 22967
rect 29043 22933 29052 22967
rect 29000 22924 29052 22933
rect 31024 22967 31076 22976
rect 31024 22933 31033 22967
rect 31033 22933 31067 22967
rect 31067 22933 31076 22967
rect 31024 22924 31076 22933
rect 32956 22967 33008 22976
rect 32956 22933 32965 22967
rect 32965 22933 32999 22967
rect 32999 22933 33008 22967
rect 32956 22924 33008 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 2504 22720 2556 22772
rect 9496 22763 9548 22772
rect 2320 22652 2372 22704
rect 3976 22652 4028 22704
rect 1952 22627 2004 22636
rect 1952 22593 1961 22627
rect 1961 22593 1995 22627
rect 1995 22593 2004 22627
rect 1952 22584 2004 22593
rect 2044 22627 2096 22636
rect 2044 22593 2053 22627
rect 2053 22593 2087 22627
rect 2087 22593 2096 22627
rect 2044 22584 2096 22593
rect 2504 22584 2556 22636
rect 2872 22627 2924 22636
rect 2872 22593 2881 22627
rect 2881 22593 2915 22627
rect 2915 22593 2924 22627
rect 2872 22584 2924 22593
rect 6920 22652 6972 22704
rect 5172 22627 5224 22636
rect 5172 22593 5181 22627
rect 5181 22593 5215 22627
rect 5215 22593 5224 22627
rect 5356 22627 5408 22636
rect 5172 22584 5224 22593
rect 5356 22593 5365 22627
rect 5365 22593 5399 22627
rect 5399 22593 5408 22627
rect 5356 22584 5408 22593
rect 8024 22652 8076 22704
rect 8484 22652 8536 22704
rect 8116 22627 8168 22636
rect 8116 22593 8125 22627
rect 8125 22593 8159 22627
rect 8159 22593 8168 22627
rect 8116 22584 8168 22593
rect 8208 22584 8260 22636
rect 8852 22627 8904 22636
rect 8852 22593 8861 22627
rect 8861 22593 8895 22627
rect 8895 22593 8904 22627
rect 8852 22584 8904 22593
rect 9036 22627 9088 22636
rect 9036 22593 9045 22627
rect 9045 22593 9079 22627
rect 9079 22593 9088 22627
rect 9036 22584 9088 22593
rect 9496 22729 9505 22763
rect 9505 22729 9539 22763
rect 9539 22729 9548 22763
rect 9496 22720 9548 22729
rect 13820 22695 13872 22704
rect 13820 22661 13829 22695
rect 13829 22661 13863 22695
rect 13863 22661 13872 22695
rect 13820 22652 13872 22661
rect 13912 22695 13964 22704
rect 13912 22661 13921 22695
rect 13921 22661 13955 22695
rect 13955 22661 13964 22695
rect 13912 22652 13964 22661
rect 4620 22448 4672 22500
rect 7380 22448 7432 22500
rect 7472 22448 7524 22500
rect 8576 22516 8628 22568
rect 12992 22584 13044 22636
rect 22652 22720 22704 22772
rect 28080 22763 28132 22772
rect 15016 22695 15068 22704
rect 15016 22661 15025 22695
rect 15025 22661 15059 22695
rect 15059 22661 15068 22695
rect 15016 22652 15068 22661
rect 14924 22627 14976 22636
rect 14280 22516 14332 22568
rect 14924 22593 14933 22627
rect 14933 22593 14967 22627
rect 14967 22593 14976 22627
rect 14924 22584 14976 22593
rect 15844 22627 15896 22636
rect 15844 22593 15853 22627
rect 15853 22593 15887 22627
rect 15887 22593 15896 22627
rect 15844 22584 15896 22593
rect 17500 22584 17552 22636
rect 18880 22627 18932 22636
rect 18880 22593 18889 22627
rect 18889 22593 18923 22627
rect 18923 22593 18932 22627
rect 18880 22584 18932 22593
rect 19340 22652 19392 22704
rect 23296 22652 23348 22704
rect 25228 22652 25280 22704
rect 28080 22729 28089 22763
rect 28089 22729 28123 22763
rect 28123 22729 28132 22763
rect 28080 22720 28132 22729
rect 31116 22720 31168 22772
rect 19064 22627 19116 22636
rect 19064 22593 19073 22627
rect 19073 22593 19107 22627
rect 19107 22593 19116 22627
rect 19064 22584 19116 22593
rect 4712 22423 4764 22432
rect 4712 22389 4721 22423
rect 4721 22389 4755 22423
rect 4755 22389 4764 22423
rect 4712 22380 4764 22389
rect 6920 22380 6972 22432
rect 15292 22423 15344 22432
rect 15292 22389 15301 22423
rect 15301 22389 15335 22423
rect 15335 22389 15344 22423
rect 15292 22380 15344 22389
rect 15936 22423 15988 22432
rect 15936 22389 15945 22423
rect 15945 22389 15979 22423
rect 15979 22389 15988 22423
rect 15936 22380 15988 22389
rect 16396 22380 16448 22432
rect 18512 22380 18564 22432
rect 19432 22584 19484 22636
rect 21640 22516 21692 22568
rect 26240 22627 26292 22636
rect 26240 22593 26249 22627
rect 26249 22593 26283 22627
rect 26283 22593 26292 22627
rect 26240 22584 26292 22593
rect 27436 22627 27488 22636
rect 19984 22448 20036 22500
rect 24584 22559 24636 22568
rect 24584 22525 24593 22559
rect 24593 22525 24627 22559
rect 24627 22525 24636 22559
rect 24584 22516 24636 22525
rect 26792 22516 26844 22568
rect 26976 22516 27028 22568
rect 25228 22448 25280 22500
rect 27436 22593 27445 22627
rect 27445 22593 27479 22627
rect 27479 22593 27488 22627
rect 27436 22584 27488 22593
rect 28908 22652 28960 22704
rect 29000 22652 29052 22704
rect 29552 22652 29604 22704
rect 27804 22627 27856 22636
rect 27804 22593 27813 22627
rect 27813 22593 27847 22627
rect 27847 22593 27856 22627
rect 27804 22584 27856 22593
rect 29092 22584 29144 22636
rect 29920 22584 29972 22636
rect 30196 22627 30248 22636
rect 30196 22593 30205 22627
rect 30205 22593 30239 22627
rect 30239 22593 30248 22627
rect 30196 22584 30248 22593
rect 30380 22627 30432 22636
rect 30380 22593 30389 22627
rect 30389 22593 30423 22627
rect 30423 22593 30432 22627
rect 30380 22584 30432 22593
rect 30472 22627 30524 22636
rect 30472 22593 30481 22627
rect 30481 22593 30515 22627
rect 30515 22593 30524 22627
rect 30472 22584 30524 22593
rect 30656 22584 30708 22636
rect 31484 22627 31536 22636
rect 31484 22593 31493 22627
rect 31493 22593 31527 22627
rect 31527 22593 31536 22627
rect 31484 22584 31536 22593
rect 29460 22448 29512 22500
rect 31116 22448 31168 22500
rect 67640 22491 67692 22500
rect 67640 22457 67649 22491
rect 67649 22457 67683 22491
rect 67683 22457 67692 22491
rect 67640 22448 67692 22457
rect 20076 22380 20128 22432
rect 22928 22380 22980 22432
rect 29000 22380 29052 22432
rect 29184 22380 29236 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 65654 22278 65706 22330
rect 65718 22278 65770 22330
rect 65782 22278 65834 22330
rect 65846 22278 65898 22330
rect 65910 22278 65962 22330
rect 1952 22176 2004 22228
rect 5172 22176 5224 22228
rect 7288 22176 7340 22228
rect 15936 22176 15988 22228
rect 19064 22176 19116 22228
rect 22836 22176 22888 22228
rect 23112 22176 23164 22228
rect 23756 22176 23808 22228
rect 27804 22176 27856 22228
rect 30380 22219 30432 22228
rect 30380 22185 30389 22219
rect 30389 22185 30423 22219
rect 30423 22185 30432 22219
rect 30380 22176 30432 22185
rect 14280 22108 14332 22160
rect 3056 22083 3108 22092
rect 3056 22049 3065 22083
rect 3065 22049 3099 22083
rect 3099 22049 3108 22083
rect 3056 22040 3108 22049
rect 5264 22040 5316 22092
rect 1676 22015 1728 22024
rect 1676 21981 1685 22015
rect 1685 21981 1719 22015
rect 1719 21981 1728 22015
rect 1676 21972 1728 21981
rect 4620 21972 4672 22024
rect 6276 22040 6328 22092
rect 7104 22040 7156 22092
rect 8116 22040 8168 22092
rect 8852 21972 8904 22024
rect 5816 21904 5868 21956
rect 9036 21904 9088 21956
rect 9312 21947 9364 21956
rect 9312 21913 9321 21947
rect 9321 21913 9355 21947
rect 9355 21913 9364 21947
rect 9312 21904 9364 21913
rect 10968 21904 11020 21956
rect 11152 22040 11204 22092
rect 14832 21972 14884 22024
rect 15844 22108 15896 22160
rect 2504 21879 2556 21888
rect 2504 21845 2513 21879
rect 2513 21845 2547 21879
rect 2547 21845 2556 21879
rect 2504 21836 2556 21845
rect 3884 21836 3936 21888
rect 6092 21836 6144 21888
rect 6552 21836 6604 21888
rect 6828 21836 6880 21888
rect 8300 21836 8352 21888
rect 10140 21836 10192 21888
rect 12808 21836 12860 21888
rect 14372 21879 14424 21888
rect 14372 21845 14381 21879
rect 14381 21845 14415 21879
rect 14415 21845 14424 21879
rect 14372 21836 14424 21845
rect 14740 21904 14792 21956
rect 15108 21947 15160 21956
rect 15108 21913 15117 21947
rect 15117 21913 15151 21947
rect 15151 21913 15160 21947
rect 15108 21904 15160 21913
rect 18052 22040 18104 22092
rect 21640 22083 21692 22092
rect 21640 22049 21649 22083
rect 21649 22049 21683 22083
rect 21683 22049 21692 22083
rect 21640 22040 21692 22049
rect 22652 22040 22704 22092
rect 28540 22108 28592 22160
rect 26240 22083 26292 22092
rect 17592 21972 17644 22024
rect 18328 22015 18380 22024
rect 18328 21981 18337 22015
rect 18337 21981 18371 22015
rect 18371 21981 18380 22015
rect 18328 21972 18380 21981
rect 18512 22015 18564 22024
rect 18512 21981 18521 22015
rect 18521 21981 18555 22015
rect 18555 21981 18564 22015
rect 18512 21972 18564 21981
rect 20260 21972 20312 22024
rect 21916 22015 21968 22024
rect 21916 21981 21925 22015
rect 21925 21981 21959 22015
rect 21959 21981 21968 22015
rect 21916 21972 21968 21981
rect 22376 22015 22428 22024
rect 22376 21981 22385 22015
rect 22385 21981 22419 22015
rect 22419 21981 22428 22015
rect 22376 21972 22428 21981
rect 26240 22049 26249 22083
rect 26249 22049 26283 22083
rect 26283 22049 26292 22083
rect 26240 22040 26292 22049
rect 30932 22083 30984 22092
rect 30932 22049 30941 22083
rect 30941 22049 30975 22083
rect 30975 22049 30984 22083
rect 30932 22040 30984 22049
rect 23572 21972 23624 22024
rect 16580 21947 16632 21956
rect 16580 21913 16589 21947
rect 16589 21913 16623 21947
rect 16623 21913 16632 21947
rect 16580 21904 16632 21913
rect 17960 21904 18012 21956
rect 22836 21904 22888 21956
rect 25872 21972 25924 22024
rect 26516 22015 26568 22024
rect 26516 21981 26525 22015
rect 26525 21981 26559 22015
rect 26559 21981 26568 22015
rect 26516 21972 26568 21981
rect 31024 21972 31076 22024
rect 17224 21836 17276 21888
rect 18880 21836 18932 21888
rect 25320 21836 25372 21888
rect 27344 21904 27396 21956
rect 29828 21904 29880 21956
rect 32956 21972 33008 22024
rect 34152 22015 34204 22024
rect 34152 21981 34161 22015
rect 34161 21981 34195 22015
rect 34195 21981 34204 22015
rect 34152 21972 34204 21981
rect 31208 21947 31260 21956
rect 31208 21913 31242 21947
rect 31242 21913 31260 21947
rect 31208 21904 31260 21913
rect 33600 21904 33652 21956
rect 28080 21836 28132 21888
rect 32128 21836 32180 21888
rect 32312 21879 32364 21888
rect 32312 21845 32321 21879
rect 32321 21845 32355 21879
rect 32355 21845 32364 21879
rect 32312 21836 32364 21845
rect 32772 21879 32824 21888
rect 32772 21845 32781 21879
rect 32781 21845 32815 21879
rect 32815 21845 32824 21879
rect 32772 21836 32824 21845
rect 35900 21879 35952 21888
rect 35900 21845 35909 21879
rect 35909 21845 35943 21879
rect 35943 21845 35952 21879
rect 35900 21836 35952 21845
rect 37648 21879 37700 21888
rect 37648 21845 37657 21879
rect 37657 21845 37691 21879
rect 37691 21845 37700 21879
rect 37648 21836 37700 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 3148 21632 3200 21684
rect 3976 21632 4028 21684
rect 7288 21632 7340 21684
rect 8024 21632 8076 21684
rect 9312 21632 9364 21684
rect 2872 21564 2924 21616
rect 4712 21607 4764 21616
rect 4712 21573 4746 21607
rect 4746 21573 4764 21607
rect 4712 21564 4764 21573
rect 3332 21496 3384 21548
rect 3884 21496 3936 21548
rect 4068 21496 4120 21548
rect 6368 21539 6420 21548
rect 6368 21505 6377 21539
rect 6377 21505 6411 21539
rect 6411 21505 6420 21539
rect 6368 21496 6420 21505
rect 6552 21539 6604 21548
rect 6552 21505 6561 21539
rect 6561 21505 6595 21539
rect 6595 21505 6604 21539
rect 6552 21496 6604 21505
rect 7748 21496 7800 21548
rect 6644 21428 6696 21480
rect 5816 21403 5868 21412
rect 5816 21369 5825 21403
rect 5825 21369 5859 21403
rect 5859 21369 5868 21403
rect 5816 21360 5868 21369
rect 1860 21292 1912 21344
rect 2596 21292 2648 21344
rect 3240 21292 3292 21344
rect 5724 21292 5776 21344
rect 11152 21564 11204 21616
rect 11612 21607 11664 21616
rect 11612 21573 11621 21607
rect 11621 21573 11655 21607
rect 11655 21573 11664 21607
rect 11612 21564 11664 21573
rect 15016 21632 15068 21684
rect 16580 21632 16632 21684
rect 17684 21632 17736 21684
rect 18052 21632 18104 21684
rect 22376 21632 22428 21684
rect 9680 21496 9732 21548
rect 12440 21539 12492 21548
rect 12440 21505 12449 21539
rect 12449 21505 12483 21539
rect 12483 21505 12492 21539
rect 12440 21496 12492 21505
rect 12716 21539 12768 21548
rect 12716 21505 12750 21539
rect 12750 21505 12768 21539
rect 12716 21496 12768 21505
rect 14372 21496 14424 21548
rect 15844 21496 15896 21548
rect 16948 21539 17000 21548
rect 16948 21505 16957 21539
rect 16957 21505 16991 21539
rect 16991 21505 17000 21539
rect 16948 21496 17000 21505
rect 17592 21496 17644 21548
rect 19800 21539 19852 21548
rect 19800 21505 19818 21539
rect 19818 21505 19852 21539
rect 19800 21496 19852 21505
rect 20076 21539 20128 21548
rect 20076 21505 20085 21539
rect 20085 21505 20119 21539
rect 20119 21505 20128 21539
rect 20076 21496 20128 21505
rect 21088 21539 21140 21548
rect 21088 21505 21097 21539
rect 21097 21505 21131 21539
rect 21131 21505 21140 21539
rect 21088 21496 21140 21505
rect 23112 21496 23164 21548
rect 23664 21539 23716 21548
rect 9220 21428 9272 21480
rect 20720 21428 20772 21480
rect 10968 21403 11020 21412
rect 10968 21369 10977 21403
rect 10977 21369 11011 21403
rect 11011 21369 11020 21403
rect 10968 21360 11020 21369
rect 20076 21360 20128 21412
rect 9036 21335 9088 21344
rect 9036 21301 9045 21335
rect 9045 21301 9079 21335
rect 9079 21301 9088 21335
rect 9036 21292 9088 21301
rect 11796 21292 11848 21344
rect 18880 21292 18932 21344
rect 23664 21505 23673 21539
rect 23673 21505 23707 21539
rect 23707 21505 23716 21539
rect 23664 21496 23716 21505
rect 26700 21632 26752 21684
rect 28908 21632 28960 21684
rect 31208 21632 31260 21684
rect 23572 21428 23624 21480
rect 25412 21539 25464 21548
rect 25412 21505 25421 21539
rect 25421 21505 25455 21539
rect 25455 21505 25464 21539
rect 25412 21496 25464 21505
rect 25504 21428 25556 21480
rect 25872 21496 25924 21548
rect 26424 21360 26476 21412
rect 27528 21496 27580 21548
rect 28540 21539 28592 21548
rect 28540 21505 28549 21539
rect 28549 21505 28583 21539
rect 28583 21505 28592 21539
rect 28540 21496 28592 21505
rect 28724 21539 28776 21548
rect 28724 21505 28733 21539
rect 28733 21505 28767 21539
rect 28767 21505 28776 21539
rect 28724 21496 28776 21505
rect 27712 21428 27764 21480
rect 32772 21564 32824 21616
rect 33968 21564 34020 21616
rect 30196 21496 30248 21548
rect 30656 21539 30708 21548
rect 30656 21505 30665 21539
rect 30665 21505 30699 21539
rect 30699 21505 30708 21539
rect 30656 21496 30708 21505
rect 30840 21539 30892 21548
rect 30840 21505 30849 21539
rect 30849 21505 30883 21539
rect 30883 21505 30892 21539
rect 30840 21496 30892 21505
rect 33416 21496 33468 21548
rect 27436 21360 27488 21412
rect 31392 21428 31444 21480
rect 32128 21428 32180 21480
rect 35624 21496 35676 21548
rect 37648 21564 37700 21616
rect 26056 21292 26108 21344
rect 27068 21292 27120 21344
rect 33140 21292 33192 21344
rect 34796 21292 34848 21344
rect 67640 21335 67692 21344
rect 67640 21301 67649 21335
rect 67649 21301 67683 21335
rect 67683 21301 67692 21335
rect 67640 21292 67692 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 65654 21190 65706 21242
rect 65718 21190 65770 21242
rect 65782 21190 65834 21242
rect 65846 21190 65898 21242
rect 65910 21190 65962 21242
rect 5724 21088 5776 21140
rect 8116 21088 8168 21140
rect 9680 21088 9732 21140
rect 12716 21088 12768 21140
rect 16948 21088 17000 21140
rect 17684 21088 17736 21140
rect 19800 21088 19852 21140
rect 4068 20952 4120 21004
rect 6644 20995 6696 21004
rect 6644 20961 6653 20995
rect 6653 20961 6687 20995
rect 6687 20961 6696 20995
rect 6644 20952 6696 20961
rect 2320 20927 2372 20936
rect 2320 20893 2329 20927
rect 2329 20893 2363 20927
rect 2363 20893 2372 20927
rect 2320 20884 2372 20893
rect 2780 20884 2832 20936
rect 8392 20884 8444 20936
rect 10600 21020 10652 21072
rect 17040 21063 17092 21072
rect 10140 20952 10192 21004
rect 10324 20884 10376 20936
rect 17040 21029 17049 21063
rect 17049 21029 17083 21063
rect 17083 21029 17092 21063
rect 17040 21020 17092 21029
rect 18236 21020 18288 21072
rect 19984 21020 20036 21072
rect 20444 21020 20496 21072
rect 21088 21020 21140 21072
rect 21732 21088 21784 21140
rect 22468 21088 22520 21140
rect 22744 21088 22796 21140
rect 6920 20859 6972 20868
rect 6920 20825 6954 20859
rect 6954 20825 6972 20859
rect 6920 20816 6972 20825
rect 7564 20816 7616 20868
rect 8116 20816 8168 20868
rect 9588 20816 9640 20868
rect 3332 20748 3384 20800
rect 6368 20748 6420 20800
rect 7840 20748 7892 20800
rect 11796 20816 11848 20868
rect 12164 20884 12216 20936
rect 15476 20927 15528 20936
rect 15476 20893 15485 20927
rect 15485 20893 15519 20927
rect 15519 20893 15528 20927
rect 15476 20884 15528 20893
rect 14372 20816 14424 20868
rect 12164 20748 12216 20800
rect 15016 20748 15068 20800
rect 15384 20816 15436 20868
rect 16304 20816 16356 20868
rect 17592 20859 17644 20868
rect 17592 20825 17601 20859
rect 17601 20825 17635 20859
rect 17635 20825 17644 20859
rect 17592 20816 17644 20825
rect 18328 20859 18380 20868
rect 18328 20825 18337 20859
rect 18337 20825 18371 20859
rect 18371 20825 18380 20859
rect 18328 20816 18380 20825
rect 18880 20816 18932 20868
rect 19156 20884 19208 20936
rect 20076 20952 20128 21004
rect 20628 20952 20680 21004
rect 19616 20927 19668 20936
rect 19616 20893 19625 20927
rect 19625 20893 19659 20927
rect 19659 20893 19668 20927
rect 19616 20884 19668 20893
rect 22376 20884 22428 20936
rect 22652 20884 22704 20936
rect 22744 20927 22796 20936
rect 22744 20893 22753 20927
rect 22753 20893 22787 20927
rect 22787 20893 22796 20927
rect 22744 20884 22796 20893
rect 20628 20816 20680 20868
rect 20260 20748 20312 20800
rect 20720 20748 20772 20800
rect 21548 20816 21600 20868
rect 23388 20952 23440 21004
rect 24860 21020 24912 21072
rect 25872 21020 25924 21072
rect 26792 20995 26844 21004
rect 23480 20927 23532 20936
rect 23480 20893 23489 20927
rect 23489 20893 23523 20927
rect 23523 20893 23532 20927
rect 23480 20884 23532 20893
rect 23664 20884 23716 20936
rect 23388 20859 23440 20868
rect 23388 20825 23397 20859
rect 23397 20825 23431 20859
rect 23431 20825 23440 20859
rect 23388 20816 23440 20825
rect 25412 20884 25464 20936
rect 26792 20961 26801 20995
rect 26801 20961 26835 20995
rect 26835 20961 26844 20995
rect 26792 20952 26844 20961
rect 28540 20952 28592 21004
rect 29092 21088 29144 21140
rect 30656 21088 30708 21140
rect 33600 21131 33652 21140
rect 33600 21097 33609 21131
rect 33609 21097 33643 21131
rect 33643 21097 33652 21131
rect 33600 21088 33652 21097
rect 35624 21131 35676 21140
rect 35624 21097 35633 21131
rect 35633 21097 35667 21131
rect 35667 21097 35676 21131
rect 35624 21088 35676 21097
rect 37648 21088 37700 21140
rect 27068 20927 27120 20936
rect 27068 20893 27102 20927
rect 27102 20893 27120 20927
rect 27068 20884 27120 20893
rect 27344 20884 27396 20936
rect 28816 20927 28868 20936
rect 28816 20893 28825 20927
rect 28825 20893 28859 20927
rect 28859 20893 28868 20927
rect 28816 20884 28868 20893
rect 30288 20884 30340 20936
rect 33140 20927 33192 20936
rect 24860 20748 24912 20800
rect 25136 20748 25188 20800
rect 29000 20816 29052 20868
rect 30104 20816 30156 20868
rect 32312 20816 32364 20868
rect 28080 20748 28132 20800
rect 28264 20748 28316 20800
rect 30840 20791 30892 20800
rect 30840 20757 30849 20791
rect 30849 20757 30883 20791
rect 30883 20757 30892 20791
rect 30840 20748 30892 20757
rect 33140 20893 33149 20927
rect 33149 20893 33183 20927
rect 33183 20893 33192 20927
rect 33140 20884 33192 20893
rect 34520 20952 34572 21004
rect 34796 20952 34848 21004
rect 34980 20927 35032 20936
rect 34980 20893 34989 20927
rect 34989 20893 35023 20927
rect 35023 20893 35032 20927
rect 34980 20884 35032 20893
rect 38200 20952 38252 21004
rect 33508 20816 33560 20868
rect 37464 20884 37516 20936
rect 35440 20816 35492 20868
rect 35716 20816 35768 20868
rect 34796 20748 34848 20800
rect 34980 20748 35032 20800
rect 36636 20791 36688 20800
rect 36636 20757 36645 20791
rect 36645 20757 36679 20791
rect 36679 20757 36688 20791
rect 36636 20748 36688 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 2872 20476 2924 20528
rect 6736 20544 6788 20596
rect 7472 20544 7524 20596
rect 7748 20587 7800 20596
rect 7748 20553 7757 20587
rect 7757 20553 7791 20587
rect 7791 20553 7800 20587
rect 7748 20544 7800 20553
rect 5632 20476 5684 20528
rect 1952 20451 2004 20460
rect 1952 20417 1961 20451
rect 1961 20417 1995 20451
rect 1995 20417 2004 20451
rect 1952 20408 2004 20417
rect 2136 20451 2188 20460
rect 2136 20417 2145 20451
rect 2145 20417 2179 20451
rect 2179 20417 2188 20451
rect 2136 20408 2188 20417
rect 3056 20451 3108 20460
rect 3056 20417 3090 20451
rect 3090 20417 3108 20451
rect 3056 20408 3108 20417
rect 4712 20408 4764 20460
rect 15384 20544 15436 20596
rect 8300 20408 8352 20460
rect 8852 20408 8904 20460
rect 10324 20451 10376 20460
rect 10324 20417 10333 20451
rect 10333 20417 10367 20451
rect 10367 20417 10376 20451
rect 10324 20408 10376 20417
rect 10600 20451 10652 20460
rect 10600 20417 10609 20451
rect 10609 20417 10643 20451
rect 10643 20417 10652 20451
rect 10600 20408 10652 20417
rect 11060 20408 11112 20460
rect 11612 20408 11664 20460
rect 15752 20451 15804 20460
rect 4160 20315 4212 20324
rect 4160 20281 4169 20315
rect 4169 20281 4203 20315
rect 4203 20281 4212 20315
rect 4160 20272 4212 20281
rect 5264 20272 5316 20324
rect 7932 20272 7984 20324
rect 8760 20340 8812 20392
rect 12440 20383 12492 20392
rect 12440 20349 12449 20383
rect 12449 20349 12483 20383
rect 12483 20349 12492 20383
rect 12440 20340 12492 20349
rect 15752 20417 15761 20451
rect 15761 20417 15795 20451
rect 15795 20417 15804 20451
rect 15752 20408 15804 20417
rect 16028 20476 16080 20528
rect 16396 20544 16448 20596
rect 20076 20544 20128 20596
rect 20720 20544 20772 20596
rect 22284 20544 22336 20596
rect 22928 20544 22980 20596
rect 24584 20544 24636 20596
rect 25504 20544 25556 20596
rect 27712 20587 27764 20596
rect 27712 20553 27721 20587
rect 27721 20553 27755 20587
rect 27755 20553 27764 20587
rect 27712 20544 27764 20553
rect 28540 20587 28592 20596
rect 28540 20553 28549 20587
rect 28549 20553 28583 20587
rect 28583 20553 28592 20587
rect 28540 20544 28592 20553
rect 35716 20587 35768 20596
rect 15568 20340 15620 20392
rect 16948 20451 17000 20460
rect 16948 20417 16957 20451
rect 16957 20417 16991 20451
rect 16991 20417 17000 20451
rect 16948 20408 17000 20417
rect 16396 20340 16448 20392
rect 17592 20408 17644 20460
rect 18328 20476 18380 20528
rect 23480 20519 23532 20528
rect 23480 20485 23489 20519
rect 23489 20485 23523 20519
rect 23523 20485 23532 20519
rect 23480 20476 23532 20485
rect 23572 20519 23624 20528
rect 23572 20485 23581 20519
rect 23581 20485 23615 20519
rect 23615 20485 23624 20519
rect 23572 20476 23624 20485
rect 18052 20408 18104 20460
rect 18236 20408 18288 20460
rect 19156 20340 19208 20392
rect 19340 20340 19392 20392
rect 21088 20408 21140 20460
rect 23204 20408 23256 20460
rect 21272 20340 21324 20392
rect 2044 20204 2096 20256
rect 4620 20204 4672 20256
rect 7288 20204 7340 20256
rect 15844 20272 15896 20324
rect 20720 20272 20772 20324
rect 23664 20272 23716 20324
rect 25228 20408 25280 20460
rect 30932 20519 30984 20528
rect 30932 20485 30941 20519
rect 30941 20485 30975 20519
rect 30975 20485 30984 20519
rect 30932 20476 30984 20485
rect 35716 20553 35725 20587
rect 35725 20553 35759 20587
rect 35759 20553 35768 20587
rect 35716 20544 35768 20553
rect 25688 20451 25740 20460
rect 25688 20417 25697 20451
rect 25697 20417 25731 20451
rect 25731 20417 25740 20451
rect 25688 20408 25740 20417
rect 25780 20451 25832 20460
rect 25780 20417 25825 20451
rect 25825 20417 25832 20451
rect 25780 20408 25832 20417
rect 29000 20408 29052 20460
rect 29276 20451 29328 20460
rect 29276 20417 29285 20451
rect 29285 20417 29319 20451
rect 29319 20417 29328 20451
rect 29276 20408 29328 20417
rect 29920 20408 29972 20460
rect 31760 20408 31812 20460
rect 33416 20408 33468 20460
rect 34704 20408 34756 20460
rect 34796 20408 34848 20460
rect 36636 20476 36688 20528
rect 28264 20340 28316 20392
rect 35532 20408 35584 20460
rect 38200 20451 38252 20460
rect 38200 20417 38209 20451
rect 38209 20417 38243 20451
rect 38243 20417 38252 20451
rect 38200 20408 38252 20417
rect 38292 20408 38344 20460
rect 24676 20272 24728 20324
rect 26884 20272 26936 20324
rect 12808 20204 12860 20256
rect 15752 20204 15804 20256
rect 16212 20204 16264 20256
rect 16672 20247 16724 20256
rect 16672 20213 16681 20247
rect 16681 20213 16715 20247
rect 16715 20213 16724 20247
rect 16672 20204 16724 20213
rect 18972 20204 19024 20256
rect 19432 20204 19484 20256
rect 19892 20247 19944 20256
rect 19892 20213 19901 20247
rect 19901 20213 19935 20247
rect 19935 20213 19944 20247
rect 19892 20204 19944 20213
rect 21548 20204 21600 20256
rect 23940 20204 23992 20256
rect 25504 20204 25556 20256
rect 31116 20272 31168 20324
rect 34152 20272 34204 20324
rect 35348 20272 35400 20324
rect 35440 20272 35492 20324
rect 37464 20315 37516 20324
rect 37464 20281 37473 20315
rect 37473 20281 37507 20315
rect 37507 20281 37516 20315
rect 37464 20272 37516 20281
rect 38200 20272 38252 20324
rect 30472 20204 30524 20256
rect 37648 20204 37700 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 65654 20102 65706 20154
rect 65718 20102 65770 20154
rect 65782 20102 65834 20154
rect 65846 20102 65898 20154
rect 65910 20102 65962 20154
rect 3056 20000 3108 20052
rect 3148 20000 3200 20052
rect 8392 20000 8444 20052
rect 12440 20000 12492 20052
rect 16028 20000 16080 20052
rect 16120 20000 16172 20052
rect 2320 19932 2372 19984
rect 4344 19932 4396 19984
rect 5356 19932 5408 19984
rect 2780 19864 2832 19916
rect 3056 19864 3108 19916
rect 4068 19864 4120 19916
rect 1860 19839 1912 19848
rect 1860 19805 1869 19839
rect 1869 19805 1903 19839
rect 1903 19805 1912 19839
rect 1860 19796 1912 19805
rect 2044 19839 2096 19848
rect 2044 19805 2053 19839
rect 2053 19805 2087 19839
rect 2087 19805 2096 19839
rect 2044 19796 2096 19805
rect 2412 19796 2464 19848
rect 4344 19839 4396 19848
rect 4344 19805 4353 19839
rect 4353 19805 4387 19839
rect 4387 19805 4396 19839
rect 4344 19796 4396 19805
rect 4528 19839 4580 19848
rect 4528 19805 4537 19839
rect 4537 19805 4571 19839
rect 4571 19805 4580 19839
rect 4528 19796 4580 19805
rect 5080 19796 5132 19848
rect 8300 19796 8352 19848
rect 9220 19839 9272 19848
rect 9220 19805 9229 19839
rect 9229 19805 9263 19839
rect 9263 19805 9272 19839
rect 9220 19796 9272 19805
rect 7288 19728 7340 19780
rect 7564 19771 7616 19780
rect 7564 19737 7573 19771
rect 7573 19737 7607 19771
rect 7607 19737 7616 19771
rect 7564 19728 7616 19737
rect 8024 19771 8076 19780
rect 8024 19737 8033 19771
rect 8033 19737 8067 19771
rect 8067 19737 8076 19771
rect 8024 19728 8076 19737
rect 2228 19660 2280 19712
rect 6736 19660 6788 19712
rect 8484 19660 8536 19712
rect 9128 19728 9180 19780
rect 16488 19932 16540 19984
rect 25688 20000 25740 20052
rect 26424 20000 26476 20052
rect 27528 20000 27580 20052
rect 30196 20000 30248 20052
rect 31760 20043 31812 20052
rect 31760 20009 31769 20043
rect 31769 20009 31803 20043
rect 31803 20009 31812 20043
rect 31760 20000 31812 20009
rect 19892 19932 19944 19984
rect 15476 19864 15528 19916
rect 19156 19864 19208 19916
rect 11336 19839 11388 19848
rect 11336 19805 11345 19839
rect 11345 19805 11379 19839
rect 11379 19805 11388 19839
rect 11336 19796 11388 19805
rect 12348 19796 12400 19848
rect 15016 19796 15068 19848
rect 16212 19839 16264 19848
rect 16212 19805 16221 19839
rect 16221 19805 16255 19839
rect 16255 19805 16264 19839
rect 16212 19796 16264 19805
rect 16672 19796 16724 19848
rect 19432 19839 19484 19848
rect 19432 19805 19441 19839
rect 19441 19805 19475 19839
rect 19475 19805 19484 19839
rect 19432 19796 19484 19805
rect 19524 19839 19576 19848
rect 19524 19805 19533 19839
rect 19533 19805 19567 19839
rect 19567 19805 19576 19839
rect 19800 19839 19852 19848
rect 19524 19796 19576 19805
rect 19800 19805 19809 19839
rect 19809 19805 19843 19839
rect 19843 19805 19852 19839
rect 19800 19796 19852 19805
rect 20260 19839 20312 19848
rect 20260 19805 20269 19839
rect 20269 19805 20303 19839
rect 20303 19805 20312 19839
rect 20260 19796 20312 19805
rect 20444 19839 20496 19848
rect 20444 19805 20453 19839
rect 20453 19805 20487 19839
rect 20487 19805 20496 19839
rect 20444 19796 20496 19805
rect 22928 19864 22980 19916
rect 14924 19728 14976 19780
rect 17592 19728 17644 19780
rect 19156 19728 19208 19780
rect 20076 19728 20128 19780
rect 21180 19796 21232 19848
rect 21272 19796 21324 19848
rect 24768 19864 24820 19916
rect 25136 19864 25188 19916
rect 25504 19864 25556 19916
rect 22652 19728 22704 19780
rect 18144 19660 18196 19712
rect 20536 19660 20588 19712
rect 22376 19660 22428 19712
rect 23664 19796 23716 19848
rect 24492 19796 24544 19848
rect 25228 19839 25280 19848
rect 25228 19805 25232 19839
rect 25232 19805 25266 19839
rect 25266 19805 25280 19839
rect 25228 19796 25280 19805
rect 25412 19839 25464 19848
rect 25412 19805 25421 19839
rect 25421 19805 25455 19839
rect 25455 19805 25464 19839
rect 25412 19796 25464 19805
rect 24952 19728 25004 19780
rect 25688 19839 25740 19848
rect 25688 19805 25697 19839
rect 25697 19805 25731 19839
rect 25731 19805 25740 19839
rect 26424 19839 26476 19848
rect 25688 19796 25740 19805
rect 26424 19805 26433 19839
rect 26433 19805 26467 19839
rect 26467 19805 26476 19839
rect 26424 19796 26476 19805
rect 26608 19839 26660 19848
rect 26608 19805 26617 19839
rect 26617 19805 26651 19839
rect 26651 19805 26660 19839
rect 26608 19796 26660 19805
rect 27436 19864 27488 19916
rect 24676 19660 24728 19712
rect 25044 19703 25096 19712
rect 25044 19669 25053 19703
rect 25053 19669 25087 19703
rect 25087 19669 25096 19703
rect 25044 19660 25096 19669
rect 25964 19728 26016 19780
rect 26148 19728 26200 19780
rect 27528 19796 27580 19848
rect 28540 19839 28592 19848
rect 28540 19805 28549 19839
rect 28549 19805 28583 19839
rect 28583 19805 28592 19839
rect 28540 19796 28592 19805
rect 29000 19932 29052 19984
rect 30288 19932 30340 19984
rect 27068 19703 27120 19712
rect 27068 19669 27077 19703
rect 27077 19669 27111 19703
rect 27111 19669 27120 19703
rect 27068 19660 27120 19669
rect 29092 19796 29144 19848
rect 30288 19839 30340 19848
rect 30288 19805 30297 19839
rect 30297 19805 30331 19839
rect 30331 19805 30340 19839
rect 30288 19796 30340 19805
rect 30196 19728 30248 19780
rect 30472 19771 30524 19780
rect 30472 19737 30481 19771
rect 30481 19737 30515 19771
rect 30515 19737 30524 19771
rect 30472 19728 30524 19737
rect 31392 19839 31444 19848
rect 31392 19805 31401 19839
rect 31401 19805 31435 19839
rect 31435 19805 31444 19839
rect 31392 19796 31444 19805
rect 29184 19660 29236 19712
rect 30380 19660 30432 19712
rect 35348 19796 35400 19848
rect 39028 19796 39080 19848
rect 68100 19839 68152 19848
rect 68100 19805 68109 19839
rect 68109 19805 68143 19839
rect 68143 19805 68152 19839
rect 68100 19796 68152 19805
rect 34704 19771 34756 19780
rect 34704 19737 34713 19771
rect 34713 19737 34747 19771
rect 34747 19737 34756 19771
rect 34704 19728 34756 19737
rect 35808 19728 35860 19780
rect 37464 19771 37516 19780
rect 37464 19737 37473 19771
rect 37473 19737 37507 19771
rect 37507 19737 37516 19771
rect 37464 19728 37516 19737
rect 37648 19771 37700 19780
rect 37648 19737 37657 19771
rect 37657 19737 37691 19771
rect 37691 19737 37700 19771
rect 37648 19728 37700 19737
rect 34796 19660 34848 19712
rect 35256 19660 35308 19712
rect 37740 19660 37792 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 2412 19456 2464 19508
rect 2688 19456 2740 19508
rect 5632 19456 5684 19508
rect 8484 19456 8536 19508
rect 9128 19499 9180 19508
rect 9128 19465 9137 19499
rect 9137 19465 9171 19499
rect 9171 19465 9180 19499
rect 9128 19456 9180 19465
rect 2228 19388 2280 19440
rect 1860 19320 1912 19372
rect 2320 19363 2372 19372
rect 2320 19329 2329 19363
rect 2329 19329 2363 19363
rect 2363 19329 2372 19363
rect 2320 19320 2372 19329
rect 3240 19320 3292 19372
rect 3424 19363 3476 19372
rect 3424 19329 3433 19363
rect 3433 19329 3467 19363
rect 3467 19329 3476 19363
rect 3424 19320 3476 19329
rect 4068 19320 4120 19372
rect 7104 19320 7156 19372
rect 8484 19363 8536 19372
rect 8484 19329 8493 19363
rect 8493 19329 8527 19363
rect 8527 19329 8536 19363
rect 8484 19320 8536 19329
rect 9220 19388 9272 19440
rect 10324 19388 10376 19440
rect 12164 19388 12216 19440
rect 14924 19431 14976 19440
rect 8760 19363 8812 19372
rect 8760 19329 8769 19363
rect 8769 19329 8803 19363
rect 8803 19329 8812 19363
rect 14924 19397 14933 19431
rect 14933 19397 14967 19431
rect 14967 19397 14976 19431
rect 14924 19388 14976 19397
rect 8760 19320 8812 19329
rect 7012 19295 7064 19304
rect 7012 19261 7021 19295
rect 7021 19261 7055 19295
rect 7055 19261 7064 19295
rect 7012 19252 7064 19261
rect 7472 19252 7524 19304
rect 8392 19252 8444 19304
rect 14464 19320 14516 19372
rect 16856 19456 16908 19508
rect 17500 19456 17552 19508
rect 20260 19456 20312 19508
rect 16488 19388 16540 19440
rect 20628 19388 20680 19440
rect 22744 19456 22796 19508
rect 26148 19456 26200 19508
rect 28540 19456 28592 19508
rect 29460 19456 29512 19508
rect 30196 19456 30248 19508
rect 35808 19499 35860 19508
rect 35808 19465 35817 19499
rect 35817 19465 35851 19499
rect 35851 19465 35860 19499
rect 35808 19456 35860 19465
rect 38292 19456 38344 19508
rect 9036 19184 9088 19236
rect 12992 19184 13044 19236
rect 15568 19252 15620 19304
rect 16396 19320 16448 19372
rect 18972 19363 19024 19372
rect 18972 19329 18981 19363
rect 18981 19329 19015 19363
rect 19015 19329 19024 19363
rect 18972 19320 19024 19329
rect 19156 19363 19208 19372
rect 19156 19329 19165 19363
rect 19165 19329 19199 19363
rect 19199 19329 19208 19363
rect 19156 19320 19208 19329
rect 19432 19320 19484 19372
rect 20536 19363 20588 19372
rect 17316 19295 17368 19304
rect 17316 19261 17325 19295
rect 17325 19261 17359 19295
rect 17359 19261 17368 19295
rect 17316 19252 17368 19261
rect 18052 19252 18104 19304
rect 20536 19329 20545 19363
rect 20545 19329 20579 19363
rect 20579 19329 20588 19363
rect 20536 19320 20588 19329
rect 26976 19363 27028 19372
rect 26976 19329 26985 19363
rect 26985 19329 27019 19363
rect 27019 19329 27028 19363
rect 26976 19320 27028 19329
rect 27068 19320 27120 19372
rect 30932 19388 30984 19440
rect 31116 19388 31168 19440
rect 29184 19320 29236 19372
rect 20444 19252 20496 19304
rect 21180 19295 21232 19304
rect 21180 19261 21189 19295
rect 21189 19261 21223 19295
rect 21223 19261 21232 19295
rect 21180 19252 21232 19261
rect 21364 19252 21416 19304
rect 25136 19252 25188 19304
rect 33508 19388 33560 19440
rect 33876 19320 33928 19372
rect 34796 19320 34848 19372
rect 35164 19363 35216 19372
rect 35164 19329 35173 19363
rect 35173 19329 35207 19363
rect 35207 19329 35216 19363
rect 35164 19320 35216 19329
rect 35256 19320 35308 19372
rect 35716 19320 35768 19372
rect 37556 19363 37608 19372
rect 37556 19329 37565 19363
rect 37565 19329 37599 19363
rect 37599 19329 37608 19363
rect 37556 19320 37608 19329
rect 37740 19363 37792 19372
rect 37740 19329 37749 19363
rect 37749 19329 37783 19363
rect 37783 19329 37792 19363
rect 37740 19320 37792 19329
rect 33140 19252 33192 19304
rect 37372 19252 37424 19304
rect 38200 19320 38252 19372
rect 39212 19320 39264 19372
rect 39028 19252 39080 19304
rect 16396 19184 16448 19236
rect 22836 19184 22888 19236
rect 33692 19184 33744 19236
rect 35348 19184 35400 19236
rect 5172 19116 5224 19168
rect 13084 19159 13136 19168
rect 13084 19125 13093 19159
rect 13093 19125 13127 19159
rect 13127 19125 13136 19159
rect 13084 19116 13136 19125
rect 15384 19159 15436 19168
rect 15384 19125 15393 19159
rect 15393 19125 15427 19159
rect 15427 19125 15436 19159
rect 15384 19116 15436 19125
rect 20628 19116 20680 19168
rect 23664 19116 23716 19168
rect 28356 19159 28408 19168
rect 28356 19125 28365 19159
rect 28365 19125 28399 19159
rect 28399 19125 28408 19159
rect 28356 19116 28408 19125
rect 33324 19159 33376 19168
rect 33324 19125 33333 19159
rect 33333 19125 33367 19159
rect 33367 19125 33376 19159
rect 33324 19116 33376 19125
rect 35164 19116 35216 19168
rect 35624 19116 35676 19168
rect 37924 19116 37976 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 65654 19014 65706 19066
rect 65718 19014 65770 19066
rect 65782 19014 65834 19066
rect 65846 19014 65898 19066
rect 65910 19014 65962 19066
rect 2320 18912 2372 18964
rect 3240 18912 3292 18964
rect 7012 18912 7064 18964
rect 12992 18912 13044 18964
rect 15844 18912 15896 18964
rect 20720 18912 20772 18964
rect 21272 18912 21324 18964
rect 24492 18912 24544 18964
rect 26608 18912 26660 18964
rect 29460 18912 29512 18964
rect 34520 18912 34572 18964
rect 37096 18912 37148 18964
rect 38936 18912 38988 18964
rect 39212 18955 39264 18964
rect 39212 18921 39221 18955
rect 39221 18921 39255 18955
rect 39255 18921 39264 18955
rect 39212 18912 39264 18921
rect 14372 18844 14424 18896
rect 18328 18844 18380 18896
rect 19156 18844 19208 18896
rect 7104 18776 7156 18828
rect 9680 18776 9732 18828
rect 2136 18751 2188 18760
rect 2136 18717 2145 18751
rect 2145 18717 2179 18751
rect 2179 18717 2188 18751
rect 2136 18708 2188 18717
rect 4988 18708 5040 18760
rect 5172 18640 5224 18692
rect 7840 18708 7892 18760
rect 7932 18708 7984 18760
rect 8760 18708 8812 18760
rect 10968 18751 11020 18760
rect 8852 18640 8904 18692
rect 10968 18717 10977 18751
rect 10977 18717 11011 18751
rect 11011 18717 11020 18751
rect 10968 18708 11020 18717
rect 12440 18708 12492 18760
rect 15476 18751 15528 18760
rect 15476 18717 15485 18751
rect 15485 18717 15519 18751
rect 15519 18717 15528 18751
rect 15476 18708 15528 18717
rect 11520 18640 11572 18692
rect 9036 18572 9088 18624
rect 10508 18572 10560 18624
rect 12624 18640 12676 18692
rect 13176 18615 13228 18624
rect 13176 18581 13185 18615
rect 13185 18581 13219 18615
rect 13219 18581 13228 18615
rect 13176 18572 13228 18581
rect 14464 18572 14516 18624
rect 15384 18640 15436 18692
rect 16396 18751 16448 18760
rect 16396 18717 16405 18751
rect 16405 18717 16439 18751
rect 16439 18717 16448 18751
rect 16396 18708 16448 18717
rect 16672 18751 16724 18760
rect 16672 18717 16681 18751
rect 16681 18717 16715 18751
rect 16715 18717 16724 18751
rect 16672 18708 16724 18717
rect 16764 18751 16816 18760
rect 16764 18717 16773 18751
rect 16773 18717 16807 18751
rect 16807 18717 16816 18751
rect 16764 18708 16816 18717
rect 17316 18708 17368 18760
rect 17500 18751 17552 18760
rect 17500 18717 17509 18751
rect 17509 18717 17543 18751
rect 17543 18717 17552 18751
rect 17500 18708 17552 18717
rect 18052 18708 18104 18760
rect 18328 18751 18380 18760
rect 18328 18717 18337 18751
rect 18337 18717 18371 18751
rect 18371 18717 18380 18751
rect 18328 18708 18380 18717
rect 18696 18776 18748 18828
rect 19432 18776 19484 18828
rect 34612 18844 34664 18896
rect 35716 18844 35768 18896
rect 37280 18844 37332 18896
rect 20260 18776 20312 18828
rect 15752 18640 15804 18692
rect 19340 18708 19392 18760
rect 19984 18708 20036 18760
rect 20444 18708 20496 18760
rect 21364 18776 21416 18828
rect 21640 18776 21692 18828
rect 21180 18708 21232 18760
rect 26976 18776 27028 18828
rect 22008 18708 22060 18760
rect 22100 18751 22152 18760
rect 22100 18717 22109 18751
rect 22109 18717 22143 18751
rect 22143 18717 22152 18751
rect 22100 18708 22152 18717
rect 22468 18708 22520 18760
rect 24952 18708 25004 18760
rect 28356 18708 28408 18760
rect 28816 18751 28868 18760
rect 28816 18717 28825 18751
rect 28825 18717 28859 18751
rect 28859 18717 28868 18751
rect 28816 18708 28868 18717
rect 29552 18708 29604 18760
rect 30196 18708 30248 18760
rect 35348 18776 35400 18828
rect 39028 18776 39080 18828
rect 32956 18708 33008 18760
rect 33140 18751 33192 18760
rect 33140 18717 33149 18751
rect 33149 18717 33183 18751
rect 33183 18717 33192 18751
rect 33140 18708 33192 18717
rect 33600 18708 33652 18760
rect 37556 18708 37608 18760
rect 37832 18708 37884 18760
rect 24124 18640 24176 18692
rect 16948 18615 17000 18624
rect 16948 18581 16957 18615
rect 16957 18581 16991 18615
rect 16991 18581 17000 18615
rect 16948 18572 17000 18581
rect 17408 18572 17460 18624
rect 20812 18572 20864 18624
rect 20904 18572 20956 18624
rect 24584 18615 24636 18624
rect 24584 18581 24593 18615
rect 24593 18581 24627 18615
rect 24627 18581 24636 18615
rect 24584 18572 24636 18581
rect 28172 18572 28224 18624
rect 28816 18572 28868 18624
rect 29000 18572 29052 18624
rect 31484 18640 31536 18692
rect 31944 18640 31996 18692
rect 38108 18640 38160 18692
rect 31024 18572 31076 18624
rect 35900 18615 35952 18624
rect 35900 18581 35909 18615
rect 35909 18581 35943 18615
rect 35943 18581 35952 18615
rect 35900 18572 35952 18581
rect 37372 18572 37424 18624
rect 38936 18751 38988 18760
rect 38936 18717 38945 18751
rect 38945 18717 38979 18751
rect 38979 18717 38988 18751
rect 38936 18708 38988 18717
rect 68100 18751 68152 18760
rect 68100 18717 68109 18751
rect 68109 18717 68143 18751
rect 68143 18717 68152 18751
rect 68100 18708 68152 18717
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 8024 18368 8076 18420
rect 11520 18411 11572 18420
rect 11520 18377 11529 18411
rect 11529 18377 11563 18411
rect 11563 18377 11572 18411
rect 11520 18368 11572 18377
rect 1860 18275 1912 18284
rect 1860 18241 1869 18275
rect 1869 18241 1903 18275
rect 1903 18241 1912 18275
rect 1860 18232 1912 18241
rect 2044 18275 2096 18284
rect 2044 18241 2048 18275
rect 2048 18241 2082 18275
rect 2082 18241 2096 18275
rect 2044 18232 2096 18241
rect 2136 18275 2188 18284
rect 2136 18241 2145 18275
rect 2145 18241 2179 18275
rect 2179 18241 2188 18275
rect 2136 18232 2188 18241
rect 2688 18232 2740 18284
rect 3424 18300 3476 18352
rect 8852 18343 8904 18352
rect 8852 18309 8861 18343
rect 8861 18309 8895 18343
rect 8895 18309 8904 18343
rect 8852 18300 8904 18309
rect 16672 18368 16724 18420
rect 6920 18232 6972 18284
rect 8024 18232 8076 18284
rect 8300 18232 8352 18284
rect 9680 18275 9732 18284
rect 9680 18241 9689 18275
rect 9689 18241 9723 18275
rect 9723 18241 9732 18275
rect 11796 18275 11848 18284
rect 9680 18232 9732 18241
rect 11796 18241 11805 18275
rect 11805 18241 11839 18275
rect 11839 18241 11848 18275
rect 11796 18232 11848 18241
rect 13176 18300 13228 18352
rect 15844 18343 15896 18352
rect 15844 18309 15853 18343
rect 15853 18309 15887 18343
rect 15887 18309 15896 18343
rect 15844 18300 15896 18309
rect 16120 18300 16172 18352
rect 12164 18275 12216 18284
rect 10600 18164 10652 18216
rect 12164 18241 12173 18275
rect 12173 18241 12207 18275
rect 12207 18241 12216 18275
rect 12164 18232 12216 18241
rect 12256 18232 12308 18284
rect 15292 18232 15344 18284
rect 16488 18232 16540 18284
rect 16948 18300 17000 18352
rect 17132 18232 17184 18284
rect 17316 18275 17368 18284
rect 17316 18241 17325 18275
rect 17325 18241 17359 18275
rect 17359 18241 17368 18275
rect 17316 18232 17368 18241
rect 4620 18028 4672 18080
rect 6368 18071 6420 18080
rect 6368 18037 6377 18071
rect 6377 18037 6411 18071
rect 6411 18037 6420 18071
rect 6368 18028 6420 18037
rect 9496 18028 9548 18080
rect 12440 18164 12492 18216
rect 16396 18164 16448 18216
rect 20904 18368 20956 18420
rect 21916 18368 21968 18420
rect 22284 18368 22336 18420
rect 28724 18368 28776 18420
rect 28816 18368 28868 18420
rect 38108 18411 38160 18420
rect 21088 18300 21140 18352
rect 21180 18300 21232 18352
rect 18696 18275 18748 18284
rect 18696 18241 18705 18275
rect 18705 18241 18739 18275
rect 18739 18241 18748 18275
rect 18696 18232 18748 18241
rect 20076 18232 20128 18284
rect 20536 18275 20588 18284
rect 16764 18096 16816 18148
rect 19432 18096 19484 18148
rect 20536 18241 20544 18275
rect 20544 18241 20578 18275
rect 20578 18241 20588 18275
rect 20536 18232 20588 18241
rect 20628 18275 20680 18284
rect 20628 18241 20637 18275
rect 20637 18241 20671 18275
rect 20671 18241 20680 18275
rect 21272 18275 21324 18284
rect 20628 18232 20680 18241
rect 21272 18241 21281 18275
rect 21281 18241 21315 18275
rect 21315 18241 21324 18275
rect 21272 18232 21324 18241
rect 12716 18028 12768 18080
rect 17132 18028 17184 18080
rect 19984 18071 20036 18080
rect 19984 18037 19993 18071
rect 19993 18037 20027 18071
rect 20027 18037 20036 18071
rect 19984 18028 20036 18037
rect 20720 18096 20772 18148
rect 24124 18343 24176 18352
rect 24124 18309 24142 18343
rect 24142 18309 24176 18343
rect 24124 18300 24176 18309
rect 28448 18300 28500 18352
rect 26332 18275 26384 18284
rect 26332 18241 26341 18275
rect 26341 18241 26375 18275
rect 26375 18241 26384 18275
rect 38108 18377 38117 18411
rect 38117 18377 38151 18411
rect 38151 18377 38160 18411
rect 38108 18368 38160 18377
rect 30288 18300 30340 18352
rect 26332 18232 26384 18241
rect 31024 18275 31076 18284
rect 31024 18241 31033 18275
rect 31033 18241 31067 18275
rect 31067 18241 31076 18275
rect 31024 18232 31076 18241
rect 33324 18300 33376 18352
rect 37464 18300 37516 18352
rect 24400 18207 24452 18216
rect 24400 18173 24409 18207
rect 24409 18173 24443 18207
rect 24443 18173 24452 18207
rect 24400 18164 24452 18173
rect 25228 18164 25280 18216
rect 27620 18164 27672 18216
rect 28172 18164 28224 18216
rect 28724 18164 28776 18216
rect 29736 18207 29788 18216
rect 28448 18096 28500 18148
rect 29736 18173 29745 18207
rect 29745 18173 29779 18207
rect 29779 18173 29788 18207
rect 29736 18164 29788 18173
rect 31116 18164 31168 18216
rect 33508 18164 33560 18216
rect 29184 18139 29236 18148
rect 29184 18105 29193 18139
rect 29193 18105 29227 18139
rect 29227 18105 29236 18139
rect 29184 18096 29236 18105
rect 30288 18096 30340 18148
rect 31392 18096 31444 18148
rect 34704 18232 34756 18284
rect 35348 18275 35400 18284
rect 35348 18241 35357 18275
rect 35357 18241 35391 18275
rect 35391 18241 35400 18275
rect 35348 18232 35400 18241
rect 35440 18232 35492 18284
rect 37924 18275 37976 18284
rect 37924 18241 37933 18275
rect 37933 18241 37967 18275
rect 37967 18241 37976 18275
rect 37924 18232 37976 18241
rect 38660 18232 38712 18284
rect 39028 18207 39080 18216
rect 39028 18173 39037 18207
rect 39037 18173 39071 18207
rect 39071 18173 39080 18207
rect 39028 18164 39080 18173
rect 31024 18028 31076 18080
rect 33416 18028 33468 18080
rect 36728 18071 36780 18080
rect 36728 18037 36737 18071
rect 36737 18037 36771 18071
rect 36771 18037 36780 18071
rect 36728 18028 36780 18037
rect 40408 18071 40460 18080
rect 40408 18037 40417 18071
rect 40417 18037 40451 18071
rect 40451 18037 40460 18071
rect 40408 18028 40460 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 65654 17926 65706 17978
rect 65718 17926 65770 17978
rect 65782 17926 65834 17978
rect 65846 17926 65898 17978
rect 65910 17926 65962 17978
rect 2688 17867 2740 17876
rect 2688 17833 2697 17867
rect 2697 17833 2731 17867
rect 2731 17833 2740 17867
rect 2688 17824 2740 17833
rect 12256 17824 12308 17876
rect 20536 17824 20588 17876
rect 22284 17824 22336 17876
rect 24768 17867 24820 17876
rect 24768 17833 24777 17867
rect 24777 17833 24811 17867
rect 24811 17833 24820 17867
rect 24768 17824 24820 17833
rect 26976 17824 27028 17876
rect 2044 17688 2096 17740
rect 7104 17688 7156 17740
rect 7380 17688 7432 17740
rect 8208 17688 8260 17740
rect 4620 17620 4672 17672
rect 5356 17620 5408 17672
rect 9404 17663 9456 17672
rect 4804 17552 4856 17604
rect 7104 17552 7156 17604
rect 9404 17629 9413 17663
rect 9413 17629 9447 17663
rect 9447 17629 9456 17663
rect 9404 17620 9456 17629
rect 9496 17620 9548 17672
rect 9680 17663 9732 17672
rect 9680 17629 9689 17663
rect 9689 17629 9723 17663
rect 9723 17629 9732 17663
rect 9680 17620 9732 17629
rect 12440 17688 12492 17740
rect 16028 17620 16080 17672
rect 16856 17663 16908 17672
rect 16856 17629 16865 17663
rect 16865 17629 16899 17663
rect 16899 17629 16908 17663
rect 16856 17620 16908 17629
rect 17408 17688 17460 17740
rect 17040 17663 17092 17672
rect 17040 17629 17049 17663
rect 17049 17629 17083 17663
rect 17083 17629 17092 17663
rect 17040 17620 17092 17629
rect 17316 17620 17368 17672
rect 18144 17663 18196 17672
rect 18144 17629 18153 17663
rect 18153 17629 18187 17663
rect 18187 17629 18196 17663
rect 18144 17620 18196 17629
rect 18328 17663 18380 17672
rect 18328 17629 18337 17663
rect 18337 17629 18371 17663
rect 18371 17629 18380 17663
rect 18328 17620 18380 17629
rect 18696 17620 18748 17672
rect 20904 17756 20956 17808
rect 20076 17620 20128 17672
rect 24308 17688 24360 17740
rect 27988 17824 28040 17876
rect 33876 17867 33928 17876
rect 29736 17688 29788 17740
rect 31760 17688 31812 17740
rect 33140 17688 33192 17740
rect 33876 17833 33885 17867
rect 33885 17833 33919 17867
rect 33919 17833 33928 17867
rect 33876 17824 33928 17833
rect 35440 17824 35492 17876
rect 37280 17867 37332 17876
rect 37280 17833 37289 17867
rect 37289 17833 37323 17867
rect 37323 17833 37332 17867
rect 37280 17824 37332 17833
rect 33784 17756 33836 17808
rect 34612 17688 34664 17740
rect 37372 17756 37424 17808
rect 7932 17552 7984 17604
rect 8300 17595 8352 17604
rect 8300 17561 8309 17595
rect 8309 17561 8343 17595
rect 8343 17561 8352 17595
rect 8300 17552 8352 17561
rect 12624 17552 12676 17604
rect 6644 17484 6696 17536
rect 8116 17484 8168 17536
rect 11796 17484 11848 17536
rect 13544 17484 13596 17536
rect 15936 17527 15988 17536
rect 15936 17493 15945 17527
rect 15945 17493 15979 17527
rect 15979 17493 15988 17527
rect 15936 17484 15988 17493
rect 16028 17484 16080 17536
rect 19432 17552 19484 17604
rect 18696 17527 18748 17536
rect 18696 17493 18705 17527
rect 18705 17493 18739 17527
rect 18739 17493 18748 17527
rect 18696 17484 18748 17493
rect 18972 17484 19024 17536
rect 20628 17552 20680 17604
rect 20812 17663 20864 17672
rect 20812 17629 20821 17663
rect 20821 17629 20855 17663
rect 20855 17629 20864 17663
rect 24584 17663 24636 17672
rect 20812 17620 20864 17629
rect 24584 17629 24593 17663
rect 24593 17629 24627 17663
rect 24627 17629 24636 17663
rect 24584 17620 24636 17629
rect 25136 17620 25188 17672
rect 21180 17552 21232 17604
rect 21364 17595 21416 17604
rect 21364 17561 21373 17595
rect 21373 17561 21407 17595
rect 21407 17561 21416 17595
rect 21364 17552 21416 17561
rect 24492 17552 24544 17604
rect 24676 17552 24728 17604
rect 25872 17595 25924 17604
rect 25872 17561 25881 17595
rect 25881 17561 25915 17595
rect 25915 17561 25924 17595
rect 25872 17552 25924 17561
rect 27068 17552 27120 17604
rect 27252 17552 27304 17604
rect 27344 17552 27396 17604
rect 21272 17484 21324 17536
rect 23204 17527 23256 17536
rect 23204 17493 23213 17527
rect 23213 17493 23247 17527
rect 23247 17493 23256 17527
rect 23204 17484 23256 17493
rect 26516 17527 26568 17536
rect 26516 17493 26525 17527
rect 26525 17493 26559 17527
rect 26559 17493 26568 17527
rect 26516 17484 26568 17493
rect 26608 17484 26660 17536
rect 27988 17484 28040 17536
rect 29184 17620 29236 17672
rect 29276 17620 29328 17672
rect 30840 17620 30892 17672
rect 31392 17620 31444 17672
rect 32312 17620 32364 17672
rect 33232 17663 33284 17672
rect 33232 17629 33241 17663
rect 33241 17629 33275 17663
rect 33275 17629 33284 17663
rect 33232 17620 33284 17629
rect 33416 17663 33468 17672
rect 33416 17629 33425 17663
rect 33425 17629 33459 17663
rect 33459 17629 33468 17663
rect 33416 17620 33468 17629
rect 33508 17663 33560 17672
rect 33508 17629 33517 17663
rect 33517 17629 33551 17663
rect 33551 17629 33560 17663
rect 33508 17620 33560 17629
rect 34796 17620 34848 17672
rect 29092 17484 29144 17536
rect 31392 17484 31444 17536
rect 33968 17484 34020 17536
rect 34704 17484 34756 17536
rect 35532 17552 35584 17604
rect 35624 17484 35676 17536
rect 35808 17663 35860 17672
rect 35808 17629 35817 17663
rect 35817 17629 35851 17663
rect 35851 17629 35860 17663
rect 35808 17620 35860 17629
rect 37464 17620 37516 17672
rect 37832 17663 37884 17672
rect 37832 17629 37841 17663
rect 37841 17629 37875 17663
rect 37875 17629 37884 17663
rect 37832 17620 37884 17629
rect 38016 17663 38068 17672
rect 38016 17629 38025 17663
rect 38025 17629 38059 17663
rect 38059 17629 38068 17663
rect 38016 17620 38068 17629
rect 38292 17824 38344 17876
rect 38660 17824 38712 17876
rect 38752 17620 38804 17672
rect 40408 17620 40460 17672
rect 36636 17595 36688 17604
rect 36636 17561 36645 17595
rect 36645 17561 36679 17595
rect 36679 17561 36688 17595
rect 36636 17552 36688 17561
rect 37740 17552 37792 17604
rect 38844 17552 38896 17604
rect 39304 17595 39356 17604
rect 39304 17561 39313 17595
rect 39313 17561 39347 17595
rect 39347 17561 39356 17595
rect 39304 17552 39356 17561
rect 35808 17484 35860 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 2412 17280 2464 17332
rect 2320 17212 2372 17264
rect 1860 17187 1912 17196
rect 1860 17153 1869 17187
rect 1869 17153 1903 17187
rect 1903 17153 1912 17187
rect 1860 17144 1912 17153
rect 5080 17144 5132 17196
rect 6920 17280 6972 17332
rect 6368 17212 6420 17264
rect 6644 17212 6696 17264
rect 14556 17280 14608 17332
rect 4988 17076 5040 17128
rect 6276 17144 6328 17196
rect 6920 17144 6972 17196
rect 7104 17144 7156 17196
rect 7380 17187 7432 17196
rect 7380 17153 7389 17187
rect 7389 17153 7423 17187
rect 7423 17153 7432 17187
rect 7380 17144 7432 17153
rect 2228 16983 2280 16992
rect 2228 16949 2237 16983
rect 2237 16949 2271 16983
rect 2271 16949 2280 16983
rect 2228 16940 2280 16949
rect 7564 17187 7616 17196
rect 7564 17153 7573 17187
rect 7573 17153 7607 17187
rect 7607 17153 7616 17187
rect 7564 17144 7616 17153
rect 8024 17144 8076 17196
rect 10968 17212 11020 17264
rect 10508 17187 10560 17196
rect 10508 17153 10517 17187
rect 10517 17153 10551 17187
rect 10551 17153 10560 17187
rect 10508 17144 10560 17153
rect 12440 17212 12492 17264
rect 12900 17212 12952 17264
rect 13452 17212 13504 17264
rect 11612 17144 11664 17196
rect 13268 17144 13320 17196
rect 13544 17187 13596 17196
rect 13544 17153 13553 17187
rect 13553 17153 13587 17187
rect 13587 17153 13596 17187
rect 13544 17144 13596 17153
rect 15844 17280 15896 17332
rect 17040 17323 17092 17332
rect 17040 17289 17049 17323
rect 17049 17289 17083 17323
rect 17083 17289 17092 17323
rect 17040 17280 17092 17289
rect 24492 17280 24544 17332
rect 25320 17280 25372 17332
rect 27344 17323 27396 17332
rect 27344 17289 27353 17323
rect 27353 17289 27387 17323
rect 27387 17289 27396 17323
rect 27344 17280 27396 17289
rect 15936 17212 15988 17264
rect 18788 17212 18840 17264
rect 15844 17187 15896 17196
rect 12716 17076 12768 17128
rect 15844 17153 15853 17187
rect 15853 17153 15887 17187
rect 15887 17153 15896 17187
rect 15844 17144 15896 17153
rect 16672 17187 16724 17196
rect 16672 17153 16681 17187
rect 16681 17153 16715 17187
rect 16715 17153 16724 17187
rect 16672 17144 16724 17153
rect 18880 17187 18932 17196
rect 18880 17153 18889 17187
rect 18889 17153 18923 17187
rect 18923 17153 18932 17187
rect 18880 17144 18932 17153
rect 26516 17212 26568 17264
rect 27712 17280 27764 17332
rect 27804 17280 27856 17332
rect 29276 17280 29328 17332
rect 31944 17280 31996 17332
rect 27896 17212 27948 17264
rect 28632 17255 28684 17264
rect 28632 17221 28641 17255
rect 28641 17221 28675 17255
rect 28675 17221 28684 17255
rect 28632 17212 28684 17221
rect 29644 17255 29696 17264
rect 29644 17221 29653 17255
rect 29653 17221 29687 17255
rect 29687 17221 29696 17255
rect 29644 17212 29696 17221
rect 31392 17212 31444 17264
rect 31760 17212 31812 17264
rect 37740 17280 37792 17332
rect 38844 17280 38896 17332
rect 16856 17076 16908 17128
rect 18328 17076 18380 17128
rect 7840 16940 7892 16992
rect 9864 16940 9916 16992
rect 10416 16940 10468 16992
rect 20076 17144 20128 17196
rect 20812 17187 20864 17196
rect 20812 17153 20821 17187
rect 20821 17153 20855 17187
rect 20855 17153 20864 17187
rect 20812 17144 20864 17153
rect 20904 17187 20956 17196
rect 20904 17153 20949 17187
rect 20949 17153 20956 17187
rect 20904 17144 20956 17153
rect 22100 17144 22152 17196
rect 24492 17187 24544 17196
rect 24492 17153 24501 17187
rect 24501 17153 24535 17187
rect 24535 17153 24544 17187
rect 24492 17144 24544 17153
rect 25136 17187 25188 17196
rect 25136 17153 25145 17187
rect 25145 17153 25179 17187
rect 25179 17153 25188 17187
rect 25136 17144 25188 17153
rect 23572 17119 23624 17128
rect 23572 17085 23581 17119
rect 23581 17085 23615 17119
rect 23615 17085 23624 17119
rect 23572 17076 23624 17085
rect 24308 17076 24360 17128
rect 27528 17144 27580 17196
rect 27804 17187 27856 17196
rect 27804 17153 27813 17187
rect 27813 17153 27847 17187
rect 27847 17153 27856 17187
rect 27804 17144 27856 17153
rect 20904 17008 20956 17060
rect 25688 17008 25740 17060
rect 26608 17008 26660 17060
rect 26792 17008 26844 17060
rect 29092 17144 29144 17196
rect 29552 17187 29604 17196
rect 29552 17153 29561 17187
rect 29561 17153 29595 17187
rect 29595 17153 29604 17187
rect 29552 17144 29604 17153
rect 28908 17076 28960 17128
rect 30012 17144 30064 17196
rect 31024 17187 31076 17196
rect 31024 17153 31033 17187
rect 31033 17153 31067 17187
rect 31067 17153 31076 17187
rect 31024 17144 31076 17153
rect 31116 17187 31168 17196
rect 31116 17153 31125 17187
rect 31125 17153 31159 17187
rect 31159 17153 31168 17187
rect 31116 17144 31168 17153
rect 31484 17144 31536 17196
rect 30932 17076 30984 17128
rect 14004 16983 14056 16992
rect 14004 16949 14013 16983
rect 14013 16949 14047 16983
rect 14047 16949 14056 16983
rect 14004 16940 14056 16949
rect 20628 16940 20680 16992
rect 26240 16940 26292 16992
rect 29368 16983 29420 16992
rect 29368 16949 29377 16983
rect 29377 16949 29411 16983
rect 29411 16949 29420 16983
rect 29368 16940 29420 16949
rect 29736 17008 29788 17060
rect 32956 17212 33008 17264
rect 33140 17144 33192 17196
rect 35348 17144 35400 17196
rect 35624 17144 35676 17196
rect 37372 17144 37424 17196
rect 37832 17187 37884 17196
rect 37832 17153 37841 17187
rect 37841 17153 37875 17187
rect 37875 17153 37884 17187
rect 37832 17144 37884 17153
rect 38384 17144 38436 17196
rect 39028 17144 39080 17196
rect 38108 17008 38160 17060
rect 67640 17051 67692 17060
rect 67640 17017 67649 17051
rect 67649 17017 67683 17051
rect 67683 17017 67692 17051
rect 67640 17008 67692 17017
rect 31024 16940 31076 16992
rect 32496 16983 32548 16992
rect 32496 16949 32505 16983
rect 32505 16949 32539 16983
rect 32539 16949 32548 16983
rect 32496 16940 32548 16949
rect 37280 16983 37332 16992
rect 37280 16949 37289 16983
rect 37289 16949 37323 16983
rect 37323 16949 37332 16983
rect 37280 16940 37332 16949
rect 40592 16983 40644 16992
rect 40592 16949 40601 16983
rect 40601 16949 40635 16983
rect 40635 16949 40644 16983
rect 40592 16940 40644 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 65654 16838 65706 16890
rect 65718 16838 65770 16890
rect 65782 16838 65834 16890
rect 65846 16838 65898 16890
rect 65910 16838 65962 16890
rect 3240 16779 3292 16788
rect 3240 16745 3249 16779
rect 3249 16745 3283 16779
rect 3283 16745 3292 16779
rect 3240 16736 3292 16745
rect 5080 16736 5132 16788
rect 7380 16736 7432 16788
rect 10784 16736 10836 16788
rect 2044 16575 2096 16584
rect 2044 16541 2053 16575
rect 2053 16541 2087 16575
rect 2087 16541 2096 16575
rect 2044 16532 2096 16541
rect 2228 16575 2280 16584
rect 2228 16541 2232 16575
rect 2232 16541 2266 16575
rect 2266 16541 2280 16575
rect 2228 16532 2280 16541
rect 3240 16532 3292 16584
rect 3792 16575 3844 16584
rect 3792 16541 3801 16575
rect 3801 16541 3835 16575
rect 3835 16541 3844 16575
rect 3792 16532 3844 16541
rect 6644 16600 6696 16652
rect 7656 16668 7708 16720
rect 8116 16600 8168 16652
rect 8760 16600 8812 16652
rect 9404 16600 9456 16652
rect 6368 16532 6420 16584
rect 6552 16532 6604 16584
rect 10416 16575 10468 16584
rect 10416 16541 10425 16575
rect 10425 16541 10459 16575
rect 10459 16541 10468 16575
rect 10416 16532 10468 16541
rect 10508 16575 10560 16584
rect 10508 16541 10517 16575
rect 10517 16541 10551 16575
rect 10551 16541 10560 16575
rect 10508 16532 10560 16541
rect 10784 16532 10836 16584
rect 15200 16736 15252 16788
rect 16028 16736 16080 16788
rect 22100 16779 22152 16788
rect 22100 16745 22109 16779
rect 22109 16745 22143 16779
rect 22143 16745 22152 16779
rect 22100 16736 22152 16745
rect 23572 16736 23624 16788
rect 24400 16736 24452 16788
rect 16672 16668 16724 16720
rect 19432 16668 19484 16720
rect 19616 16668 19668 16720
rect 20444 16668 20496 16720
rect 21088 16668 21140 16720
rect 21364 16668 21416 16720
rect 24492 16668 24544 16720
rect 15844 16600 15896 16652
rect 16212 16600 16264 16652
rect 6276 16464 6328 16516
rect 2320 16396 2372 16448
rect 5264 16396 5316 16448
rect 6920 16464 6972 16516
rect 7564 16464 7616 16516
rect 9864 16464 9916 16516
rect 11612 16464 11664 16516
rect 13268 16532 13320 16584
rect 14004 16532 14056 16584
rect 13084 16464 13136 16516
rect 13544 16464 13596 16516
rect 17040 16532 17092 16584
rect 17316 16600 17368 16652
rect 18236 16532 18288 16584
rect 19616 16575 19668 16584
rect 17408 16464 17460 16516
rect 19616 16541 19625 16575
rect 19625 16541 19659 16575
rect 19659 16541 19668 16575
rect 19616 16532 19668 16541
rect 22652 16600 22704 16652
rect 31024 16736 31076 16788
rect 33232 16736 33284 16788
rect 34796 16779 34848 16788
rect 34796 16745 34805 16779
rect 34805 16745 34839 16779
rect 34839 16745 34848 16779
rect 34796 16736 34848 16745
rect 37280 16736 37332 16788
rect 38108 16779 38160 16788
rect 38108 16745 38117 16779
rect 38117 16745 38151 16779
rect 38151 16745 38160 16779
rect 38108 16736 38160 16745
rect 29552 16668 29604 16720
rect 29000 16600 29052 16652
rect 30840 16600 30892 16652
rect 7012 16439 7064 16448
rect 7012 16405 7021 16439
rect 7021 16405 7055 16439
rect 7055 16405 7064 16439
rect 7012 16396 7064 16405
rect 16764 16396 16816 16448
rect 18052 16439 18104 16448
rect 18052 16405 18061 16439
rect 18061 16405 18095 16439
rect 18095 16405 18104 16439
rect 18052 16396 18104 16405
rect 19432 16507 19484 16516
rect 19432 16473 19441 16507
rect 19441 16473 19475 16507
rect 19475 16473 19484 16507
rect 19432 16464 19484 16473
rect 21272 16464 21324 16516
rect 21640 16396 21692 16448
rect 21824 16575 21876 16584
rect 21824 16541 21833 16575
rect 21833 16541 21867 16575
rect 21867 16541 21876 16575
rect 21824 16532 21876 16541
rect 28172 16532 28224 16584
rect 32956 16600 33008 16652
rect 31576 16532 31628 16584
rect 32864 16532 32916 16584
rect 33416 16532 33468 16584
rect 38384 16668 38436 16720
rect 36636 16643 36688 16652
rect 36636 16609 36645 16643
rect 36645 16609 36679 16643
rect 36679 16609 36688 16643
rect 36636 16600 36688 16609
rect 25780 16464 25832 16516
rect 28908 16464 28960 16516
rect 31116 16507 31168 16516
rect 31116 16473 31125 16507
rect 31125 16473 31159 16507
rect 31159 16473 31168 16507
rect 31116 16464 31168 16473
rect 31208 16507 31260 16516
rect 31208 16473 31217 16507
rect 31217 16473 31251 16507
rect 31251 16473 31260 16507
rect 31208 16464 31260 16473
rect 32128 16464 32180 16516
rect 34520 16464 34572 16516
rect 37740 16507 37792 16516
rect 37740 16473 37749 16507
rect 37749 16473 37783 16507
rect 37783 16473 37792 16507
rect 37740 16464 37792 16473
rect 37832 16464 37884 16516
rect 40592 16464 40644 16516
rect 24308 16396 24360 16448
rect 26332 16439 26384 16448
rect 26332 16405 26341 16439
rect 26341 16405 26375 16439
rect 26375 16405 26384 16439
rect 26332 16396 26384 16405
rect 27344 16396 27396 16448
rect 31484 16396 31536 16448
rect 32588 16396 32640 16448
rect 34060 16396 34112 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 6828 16192 6880 16244
rect 11336 16192 11388 16244
rect 14372 16235 14424 16244
rect 14372 16201 14381 16235
rect 14381 16201 14415 16235
rect 14415 16201 14424 16235
rect 14372 16192 14424 16201
rect 17040 16235 17092 16244
rect 17040 16201 17049 16235
rect 17049 16201 17083 16235
rect 17083 16201 17092 16235
rect 17040 16192 17092 16201
rect 18236 16192 18288 16244
rect 21824 16235 21876 16244
rect 21824 16201 21833 16235
rect 21833 16201 21867 16235
rect 21867 16201 21876 16235
rect 21824 16192 21876 16201
rect 23112 16192 23164 16244
rect 25780 16235 25832 16244
rect 5172 16167 5224 16176
rect 5172 16133 5181 16167
rect 5181 16133 5215 16167
rect 5215 16133 5224 16167
rect 5172 16124 5224 16133
rect 2044 16099 2096 16108
rect 2044 16065 2053 16099
rect 2053 16065 2087 16099
rect 2087 16065 2096 16099
rect 2044 16056 2096 16065
rect 2228 16099 2280 16108
rect 2228 16065 2237 16099
rect 2237 16065 2271 16099
rect 2271 16065 2280 16099
rect 2228 16056 2280 16065
rect 2320 16099 2372 16108
rect 2320 16065 2329 16099
rect 2329 16065 2363 16099
rect 2363 16065 2372 16099
rect 2320 16056 2372 16065
rect 2688 16056 2740 16108
rect 4988 16056 5040 16108
rect 4896 15920 4948 15972
rect 6552 16099 6604 16108
rect 6552 16065 6561 16099
rect 6561 16065 6595 16099
rect 6595 16065 6604 16099
rect 6552 16056 6604 16065
rect 10324 16124 10376 16176
rect 13912 16124 13964 16176
rect 16672 16167 16724 16176
rect 16672 16133 16681 16167
rect 16681 16133 16715 16167
rect 16715 16133 16724 16167
rect 16672 16124 16724 16133
rect 19432 16124 19484 16176
rect 19800 16124 19852 16176
rect 25780 16201 25789 16235
rect 25789 16201 25823 16235
rect 25823 16201 25832 16235
rect 25780 16192 25832 16201
rect 7564 16099 7616 16108
rect 7564 16065 7573 16099
rect 7573 16065 7607 16099
rect 7607 16065 7616 16099
rect 7564 16056 7616 16065
rect 12440 16056 12492 16108
rect 12624 16099 12676 16108
rect 12624 16065 12633 16099
rect 12633 16065 12667 16099
rect 12667 16065 12676 16099
rect 12624 16056 12676 16065
rect 15016 16099 15068 16108
rect 15016 16065 15025 16099
rect 15025 16065 15059 16099
rect 15059 16065 15068 16099
rect 15016 16056 15068 16065
rect 7012 15988 7064 16040
rect 7748 15988 7800 16040
rect 5264 15920 5316 15972
rect 5448 15963 5500 15972
rect 5448 15929 5457 15963
rect 5457 15929 5491 15963
rect 5491 15929 5500 15963
rect 5448 15920 5500 15929
rect 6368 15920 6420 15972
rect 7564 15920 7616 15972
rect 15292 15988 15344 16040
rect 17960 16056 18012 16108
rect 18696 16056 18748 16108
rect 19708 16099 19760 16108
rect 19708 16065 19718 16099
rect 19718 16065 19752 16099
rect 19752 16065 19760 16099
rect 19708 16056 19760 16065
rect 20076 16099 20128 16108
rect 20076 16065 20090 16099
rect 20090 16065 20124 16099
rect 20124 16065 20128 16099
rect 20076 16056 20128 16065
rect 15384 15920 15436 15972
rect 15752 15988 15804 16040
rect 16396 15988 16448 16040
rect 20260 15988 20312 16040
rect 21824 15988 21876 16040
rect 22928 16056 22980 16108
rect 25136 16124 25188 16176
rect 25320 16124 25372 16176
rect 25964 16056 26016 16108
rect 26332 16124 26384 16176
rect 24860 15988 24912 16040
rect 25780 15988 25832 16040
rect 26240 16099 26292 16108
rect 26240 16065 26249 16099
rect 26249 16065 26283 16099
rect 26283 16065 26292 16099
rect 28908 16192 28960 16244
rect 29920 16235 29972 16244
rect 29920 16201 29929 16235
rect 29929 16201 29963 16235
rect 29963 16201 29972 16235
rect 29920 16192 29972 16201
rect 33140 16192 33192 16244
rect 34520 16235 34572 16244
rect 34520 16201 34529 16235
rect 34529 16201 34563 16235
rect 34563 16201 34572 16235
rect 34520 16192 34572 16201
rect 37740 16192 37792 16244
rect 28632 16167 28684 16176
rect 28632 16133 28641 16167
rect 28641 16133 28675 16167
rect 28675 16133 28684 16167
rect 28632 16124 28684 16133
rect 26240 16056 26292 16065
rect 26792 16056 26844 16108
rect 28816 16056 28868 16108
rect 30840 16056 30892 16108
rect 31208 16099 31260 16108
rect 31208 16065 31217 16099
rect 31217 16065 31251 16099
rect 31251 16065 31260 16099
rect 31208 16056 31260 16065
rect 31668 16056 31720 16108
rect 27712 15988 27764 16040
rect 28540 15988 28592 16040
rect 19432 15920 19484 15972
rect 20352 15920 20404 15972
rect 32864 16124 32916 16176
rect 32312 16099 32364 16108
rect 32312 16065 32321 16099
rect 32321 16065 32355 16099
rect 32355 16065 32364 16099
rect 32312 16056 32364 16065
rect 32496 16099 32548 16108
rect 32496 16065 32505 16099
rect 32505 16065 32539 16099
rect 32539 16065 32548 16099
rect 32496 16056 32548 16065
rect 32680 16099 32732 16108
rect 32680 16065 32689 16099
rect 32689 16065 32723 16099
rect 32723 16065 32732 16099
rect 32680 16056 32732 16065
rect 33600 16056 33652 16108
rect 34060 16099 34112 16108
rect 34060 16065 34069 16099
rect 34069 16065 34103 16099
rect 34103 16065 34112 16099
rect 34060 16056 34112 16065
rect 32956 15988 33008 16040
rect 33692 15988 33744 16040
rect 37648 16124 37700 16176
rect 2688 15895 2740 15904
rect 2688 15861 2697 15895
rect 2697 15861 2731 15895
rect 2731 15861 2740 15895
rect 2688 15852 2740 15861
rect 6460 15895 6512 15904
rect 6460 15861 6469 15895
rect 6469 15861 6503 15895
rect 6503 15861 6512 15895
rect 6460 15852 6512 15861
rect 7196 15895 7248 15904
rect 7196 15861 7205 15895
rect 7205 15861 7239 15895
rect 7239 15861 7248 15895
rect 7196 15852 7248 15861
rect 12164 15895 12216 15904
rect 12164 15861 12173 15895
rect 12173 15861 12207 15895
rect 12207 15861 12216 15895
rect 12164 15852 12216 15861
rect 13084 15852 13136 15904
rect 13544 15895 13596 15904
rect 13544 15861 13553 15895
rect 13553 15861 13587 15895
rect 13587 15861 13596 15895
rect 13544 15852 13596 15861
rect 20444 15852 20496 15904
rect 20904 15895 20956 15904
rect 20904 15861 20913 15895
rect 20913 15861 20947 15895
rect 20947 15861 20956 15895
rect 20904 15852 20956 15861
rect 25504 15852 25556 15904
rect 25596 15852 25648 15904
rect 31392 15852 31444 15904
rect 37464 16056 37516 16108
rect 37648 15988 37700 16040
rect 38200 16056 38252 16108
rect 38844 16056 38896 16108
rect 41236 15988 41288 16040
rect 36544 15852 36596 15904
rect 38660 15852 38712 15904
rect 67640 15895 67692 15904
rect 67640 15861 67649 15895
rect 67649 15861 67683 15895
rect 67683 15861 67692 15895
rect 67640 15852 67692 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 65654 15750 65706 15802
rect 65718 15750 65770 15802
rect 65782 15750 65834 15802
rect 65846 15750 65898 15802
rect 65910 15750 65962 15802
rect 2228 15691 2280 15700
rect 2228 15657 2237 15691
rect 2237 15657 2271 15691
rect 2271 15657 2280 15691
rect 2228 15648 2280 15657
rect 6920 15648 6972 15700
rect 11336 15648 11388 15700
rect 15660 15648 15712 15700
rect 19708 15648 19760 15700
rect 19800 15648 19852 15700
rect 20812 15648 20864 15700
rect 21824 15691 21876 15700
rect 21824 15657 21833 15691
rect 21833 15657 21867 15691
rect 21867 15657 21876 15691
rect 21824 15648 21876 15657
rect 25596 15648 25648 15700
rect 27344 15691 27396 15700
rect 2688 15512 2740 15564
rect 7012 15580 7064 15632
rect 10784 15580 10836 15632
rect 1860 15487 1912 15496
rect 1860 15453 1869 15487
rect 1869 15453 1903 15487
rect 1903 15453 1912 15487
rect 1860 15444 1912 15453
rect 3148 15444 3200 15496
rect 3792 15487 3844 15496
rect 3792 15453 3801 15487
rect 3801 15453 3835 15487
rect 3835 15453 3844 15487
rect 3792 15444 3844 15453
rect 6368 15512 6420 15564
rect 8024 15512 8076 15564
rect 12716 15512 12768 15564
rect 7288 15444 7340 15496
rect 7840 15487 7892 15496
rect 7840 15453 7849 15487
rect 7849 15453 7883 15487
rect 7883 15453 7892 15487
rect 7840 15444 7892 15453
rect 5080 15376 5132 15428
rect 7748 15376 7800 15428
rect 5264 15308 5316 15360
rect 6276 15308 6328 15360
rect 6920 15308 6972 15360
rect 9680 15444 9732 15496
rect 12164 15487 12216 15496
rect 12164 15453 12173 15487
rect 12173 15453 12207 15487
rect 12207 15453 12216 15487
rect 12164 15444 12216 15453
rect 13084 15487 13136 15496
rect 13084 15453 13093 15487
rect 13093 15453 13127 15487
rect 13127 15453 13136 15487
rect 13084 15444 13136 15453
rect 13268 15487 13320 15496
rect 13268 15453 13277 15487
rect 13277 15453 13311 15487
rect 13311 15453 13320 15487
rect 13268 15444 13320 15453
rect 14188 15444 14240 15496
rect 14372 15444 14424 15496
rect 25412 15580 25464 15632
rect 16488 15444 16540 15496
rect 18052 15444 18104 15496
rect 19432 15487 19484 15496
rect 19432 15453 19441 15487
rect 19441 15453 19475 15487
rect 19475 15453 19484 15487
rect 19432 15444 19484 15453
rect 19800 15512 19852 15564
rect 13360 15376 13412 15428
rect 13544 15376 13596 15428
rect 15476 15376 15528 15428
rect 17960 15376 18012 15428
rect 20076 15444 20128 15496
rect 20720 15512 20772 15564
rect 24860 15512 24912 15564
rect 27344 15657 27353 15691
rect 27353 15657 27387 15691
rect 27387 15657 27396 15691
rect 27344 15648 27396 15657
rect 28632 15648 28684 15700
rect 37096 15648 37148 15700
rect 37740 15648 37792 15700
rect 38844 15691 38896 15700
rect 20352 15444 20404 15496
rect 22008 15487 22060 15496
rect 22008 15453 22017 15487
rect 22017 15453 22051 15487
rect 22051 15453 22060 15487
rect 22008 15444 22060 15453
rect 22100 15487 22152 15496
rect 22100 15453 22109 15487
rect 22109 15453 22143 15487
rect 22143 15453 22152 15487
rect 22284 15487 22336 15496
rect 22100 15444 22152 15453
rect 22284 15453 22293 15487
rect 22293 15453 22327 15487
rect 22327 15453 22336 15487
rect 22284 15444 22336 15453
rect 25872 15444 25924 15496
rect 26056 15487 26108 15496
rect 26056 15453 26065 15487
rect 26065 15453 26099 15487
rect 26099 15453 26108 15487
rect 26056 15444 26108 15453
rect 32864 15580 32916 15632
rect 33692 15623 33744 15632
rect 33692 15589 33701 15623
rect 33701 15589 33735 15623
rect 33735 15589 33744 15623
rect 33692 15580 33744 15589
rect 37648 15580 37700 15632
rect 38844 15657 38853 15691
rect 38853 15657 38887 15691
rect 38887 15657 38896 15691
rect 38844 15648 38896 15657
rect 27160 15487 27212 15496
rect 27160 15453 27169 15487
rect 27169 15453 27203 15487
rect 27203 15453 27212 15487
rect 27160 15444 27212 15453
rect 28172 15444 28224 15496
rect 29736 15512 29788 15564
rect 32496 15512 32548 15564
rect 25136 15376 25188 15428
rect 27252 15376 27304 15428
rect 29000 15444 29052 15496
rect 32312 15444 32364 15496
rect 35808 15512 35860 15564
rect 12624 15351 12676 15360
rect 12624 15317 12633 15351
rect 12633 15317 12667 15351
rect 12667 15317 12676 15351
rect 12624 15308 12676 15317
rect 20076 15351 20128 15360
rect 20076 15317 20085 15351
rect 20085 15317 20119 15351
rect 20119 15317 20128 15351
rect 20076 15308 20128 15317
rect 25228 15351 25280 15360
rect 25228 15317 25237 15351
rect 25237 15317 25271 15351
rect 25271 15317 25280 15351
rect 25228 15308 25280 15317
rect 28080 15351 28132 15360
rect 28080 15317 28089 15351
rect 28089 15317 28123 15351
rect 28123 15317 28132 15351
rect 28080 15308 28132 15317
rect 29460 15376 29512 15428
rect 29552 15376 29604 15428
rect 28632 15308 28684 15360
rect 31024 15308 31076 15360
rect 32588 15308 32640 15360
rect 32772 15308 32824 15360
rect 32956 15308 33008 15360
rect 35348 15376 35400 15428
rect 35992 15487 36044 15496
rect 35992 15453 36001 15487
rect 36001 15453 36035 15487
rect 36035 15453 36044 15487
rect 35992 15444 36044 15453
rect 37280 15444 37332 15496
rect 33232 15351 33284 15360
rect 33232 15317 33241 15351
rect 33241 15317 33275 15351
rect 33275 15317 33284 15351
rect 33232 15308 33284 15317
rect 33324 15308 33376 15360
rect 35716 15308 35768 15360
rect 36268 15308 36320 15360
rect 37464 15376 37516 15428
rect 41236 15555 41288 15564
rect 41236 15521 41245 15555
rect 41245 15521 41279 15555
rect 41279 15521 41288 15555
rect 41236 15512 41288 15521
rect 38476 15419 38528 15428
rect 38476 15385 38485 15419
rect 38485 15385 38519 15419
rect 38519 15385 38528 15419
rect 38476 15376 38528 15385
rect 38660 15419 38712 15428
rect 38660 15385 38669 15419
rect 38669 15385 38703 15419
rect 38703 15385 38712 15419
rect 38660 15376 38712 15385
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 3792 15104 3844 15156
rect 4804 15036 4856 15088
rect 5356 15079 5408 15088
rect 5356 15045 5365 15079
rect 5365 15045 5399 15079
rect 5399 15045 5408 15079
rect 5356 15036 5408 15045
rect 6828 15036 6880 15088
rect 4068 14968 4120 15020
rect 5080 15011 5132 15020
rect 5080 14977 5089 15011
rect 5089 14977 5123 15011
rect 5123 14977 5132 15011
rect 5080 14968 5132 14977
rect 5264 15011 5316 15020
rect 5264 14977 5273 15011
rect 5273 14977 5307 15011
rect 5307 14977 5316 15011
rect 5264 14968 5316 14977
rect 6552 14968 6604 15020
rect 7748 14968 7800 15020
rect 10140 15104 10192 15156
rect 10324 15147 10376 15156
rect 10324 15113 10333 15147
rect 10333 15113 10367 15147
rect 10367 15113 10376 15147
rect 10324 15104 10376 15113
rect 12532 15104 12584 15156
rect 15200 15104 15252 15156
rect 10232 15036 10284 15088
rect 11060 15036 11112 15088
rect 12440 15036 12492 15088
rect 12624 15036 12676 15088
rect 9036 14968 9088 15020
rect 9220 15011 9272 15020
rect 9220 14977 9254 15011
rect 9254 14977 9272 15011
rect 11888 15011 11940 15020
rect 9220 14968 9272 14977
rect 11888 14977 11897 15011
rect 11897 14977 11931 15011
rect 11931 14977 11940 15011
rect 11888 14968 11940 14977
rect 14372 15011 14424 15020
rect 14372 14977 14381 15011
rect 14381 14977 14415 15011
rect 14415 14977 14424 15011
rect 14372 14968 14424 14977
rect 17960 15104 18012 15156
rect 22008 15104 22060 15156
rect 28908 15147 28960 15156
rect 17592 15036 17644 15088
rect 18972 15036 19024 15088
rect 16488 14968 16540 15020
rect 16764 14968 16816 15020
rect 20996 15036 21048 15088
rect 24860 15036 24912 15088
rect 28908 15113 28917 15147
rect 28917 15113 28951 15147
rect 28951 15113 28960 15147
rect 28908 15104 28960 15113
rect 29552 15147 29604 15156
rect 29552 15113 29561 15147
rect 29561 15113 29595 15147
rect 29595 15113 29604 15147
rect 29552 15104 29604 15113
rect 32496 15147 32548 15156
rect 20720 15011 20772 15020
rect 20720 14977 20729 15011
rect 20729 14977 20763 15011
rect 20763 14977 20772 15011
rect 20720 14968 20772 14977
rect 22008 15011 22060 15020
rect 22008 14977 22017 15011
rect 22017 14977 22051 15011
rect 22051 14977 22060 15011
rect 22008 14968 22060 14977
rect 22284 15011 22336 15020
rect 22284 14977 22293 15011
rect 22293 14977 22327 15011
rect 22327 14977 22336 15011
rect 22284 14968 22336 14977
rect 24952 14968 25004 15020
rect 25320 14968 25372 15020
rect 6828 14900 6880 14952
rect 7196 14900 7248 14952
rect 12532 14943 12584 14952
rect 12532 14909 12541 14943
rect 12541 14909 12575 14943
rect 12575 14909 12584 14943
rect 12532 14900 12584 14909
rect 22192 14943 22244 14952
rect 22192 14909 22201 14943
rect 22201 14909 22235 14943
rect 22235 14909 22244 14943
rect 22192 14900 22244 14909
rect 24308 14943 24360 14952
rect 24308 14909 24317 14943
rect 24317 14909 24351 14943
rect 24351 14909 24360 14943
rect 24308 14900 24360 14909
rect 25228 14900 25280 14952
rect 26240 14968 26292 15020
rect 29000 14968 29052 15020
rect 5632 14875 5684 14884
rect 5632 14841 5641 14875
rect 5641 14841 5675 14875
rect 5675 14841 5684 14875
rect 5632 14832 5684 14841
rect 5724 14832 5776 14884
rect 8208 14832 8260 14884
rect 13912 14875 13964 14884
rect 13912 14841 13921 14875
rect 13921 14841 13955 14875
rect 13955 14841 13964 14875
rect 13912 14832 13964 14841
rect 22928 14875 22980 14884
rect 1952 14764 2004 14816
rect 4068 14764 4120 14816
rect 10508 14764 10560 14816
rect 11980 14764 12032 14816
rect 22376 14764 22428 14816
rect 22928 14841 22937 14875
rect 22937 14841 22971 14875
rect 22971 14841 22980 14875
rect 22928 14832 22980 14841
rect 25780 14832 25832 14884
rect 25872 14832 25924 14884
rect 29276 15036 29328 15088
rect 29644 14968 29696 15020
rect 31116 15036 31168 15088
rect 32496 15113 32505 15147
rect 32505 15113 32539 15147
rect 32539 15113 32548 15147
rect 32496 15104 32548 15113
rect 32128 15079 32180 15088
rect 32128 15045 32137 15079
rect 32137 15045 32171 15079
rect 32171 15045 32180 15079
rect 32128 15036 32180 15045
rect 32312 15079 32364 15088
rect 32312 15045 32321 15079
rect 32321 15045 32355 15079
rect 32355 15045 32364 15079
rect 35992 15104 36044 15156
rect 32312 15036 32364 15045
rect 33232 15036 33284 15088
rect 36268 15079 36320 15088
rect 36268 15045 36277 15079
rect 36277 15045 36311 15079
rect 36311 15045 36320 15079
rect 37372 15104 37424 15156
rect 38476 15104 38528 15156
rect 36268 15036 36320 15045
rect 38660 15036 38712 15088
rect 30012 15011 30064 15020
rect 30012 14977 30021 15011
rect 30021 14977 30055 15011
rect 30055 14977 30064 15011
rect 30012 14968 30064 14977
rect 31392 14968 31444 15020
rect 31484 15011 31536 15020
rect 31484 14977 31493 15011
rect 31493 14977 31527 15011
rect 31527 14977 31536 15011
rect 31484 14968 31536 14977
rect 30932 14900 30984 14952
rect 34428 14943 34480 14952
rect 34428 14909 34437 14943
rect 34437 14909 34471 14943
rect 34471 14909 34480 14943
rect 34428 14900 34480 14909
rect 35256 15011 35308 15020
rect 35256 14977 35265 15011
rect 35265 14977 35299 15011
rect 35299 14977 35308 15011
rect 35256 14968 35308 14977
rect 35440 15011 35492 15020
rect 35440 14977 35449 15011
rect 35449 14977 35483 15011
rect 35483 14977 35492 15011
rect 35440 14968 35492 14977
rect 35808 14968 35860 15020
rect 36452 15011 36504 15020
rect 36452 14977 36461 15011
rect 36461 14977 36495 15011
rect 36495 14977 36504 15011
rect 36452 14968 36504 14977
rect 37556 14968 37608 15020
rect 37740 14968 37792 15020
rect 36728 14900 36780 14952
rect 29368 14764 29420 14816
rect 36912 14832 36964 14884
rect 38016 14832 38068 14884
rect 37464 14764 37516 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 65654 14662 65706 14714
rect 65718 14662 65770 14714
rect 65782 14662 65834 14714
rect 65846 14662 65898 14714
rect 65910 14662 65962 14714
rect 9220 14560 9272 14612
rect 9772 14560 9824 14612
rect 10784 14560 10836 14612
rect 11888 14560 11940 14612
rect 17224 14603 17276 14612
rect 2136 14492 2188 14544
rect 2228 14492 2280 14544
rect 7472 14492 7524 14544
rect 1768 14399 1820 14408
rect 1768 14365 1777 14399
rect 1777 14365 1811 14399
rect 1811 14365 1820 14399
rect 1768 14356 1820 14365
rect 1952 14399 2004 14408
rect 1952 14365 1961 14399
rect 1961 14365 1995 14399
rect 1995 14365 2004 14399
rect 1952 14356 2004 14365
rect 2228 14356 2280 14408
rect 3792 14399 3844 14408
rect 3792 14365 3801 14399
rect 3801 14365 3835 14399
rect 3835 14365 3844 14399
rect 3792 14356 3844 14365
rect 4896 14356 4948 14408
rect 5264 14399 5316 14408
rect 5264 14365 5273 14399
rect 5273 14365 5307 14399
rect 5307 14365 5316 14399
rect 5264 14356 5316 14365
rect 6460 14424 6512 14476
rect 5724 14356 5776 14408
rect 6828 14399 6880 14408
rect 6828 14365 6837 14399
rect 6837 14365 6871 14399
rect 6871 14365 6880 14399
rect 6828 14356 6880 14365
rect 7840 14424 7892 14476
rect 7472 14356 7524 14408
rect 7656 14356 7708 14408
rect 9036 14424 9088 14476
rect 17224 14569 17233 14603
rect 17233 14569 17267 14603
rect 17267 14569 17276 14603
rect 17224 14560 17276 14569
rect 20168 14560 20220 14612
rect 24952 14560 25004 14612
rect 22468 14492 22520 14544
rect 25320 14492 25372 14544
rect 7196 14288 7248 14340
rect 8208 14356 8260 14408
rect 9220 14356 9272 14408
rect 14096 14356 14148 14408
rect 14464 14356 14516 14408
rect 9128 14331 9180 14340
rect 9128 14297 9137 14331
rect 9137 14297 9171 14331
rect 9171 14297 9180 14331
rect 9128 14288 9180 14297
rect 11244 14288 11296 14340
rect 11336 14288 11388 14340
rect 12256 14288 12308 14340
rect 14372 14288 14424 14340
rect 15384 14424 15436 14476
rect 16120 14424 16172 14476
rect 22376 14467 22428 14476
rect 22376 14433 22385 14467
rect 22385 14433 22419 14467
rect 22419 14433 22428 14467
rect 22376 14424 22428 14433
rect 15292 14356 15344 14408
rect 2780 14220 2832 14272
rect 5724 14263 5776 14272
rect 5724 14229 5733 14263
rect 5733 14229 5767 14263
rect 5767 14229 5776 14263
rect 5724 14220 5776 14229
rect 7012 14220 7064 14272
rect 8024 14220 8076 14272
rect 8116 14220 8168 14272
rect 8392 14263 8444 14272
rect 8392 14229 8401 14263
rect 8401 14229 8435 14263
rect 8435 14229 8444 14263
rect 8392 14220 8444 14229
rect 12624 14220 12676 14272
rect 13360 14263 13412 14272
rect 13360 14229 13369 14263
rect 13369 14229 13403 14263
rect 13403 14229 13412 14263
rect 13360 14220 13412 14229
rect 15936 14399 15988 14408
rect 15936 14365 15946 14399
rect 15946 14365 15980 14399
rect 15980 14365 15988 14399
rect 15936 14356 15988 14365
rect 17132 14399 17184 14408
rect 17132 14365 17141 14399
rect 17141 14365 17175 14399
rect 17175 14365 17184 14399
rect 17132 14356 17184 14365
rect 20168 14356 20220 14408
rect 20720 14399 20772 14408
rect 20720 14365 20729 14399
rect 20729 14365 20763 14399
rect 20763 14365 20772 14399
rect 20720 14356 20772 14365
rect 23940 14356 23992 14408
rect 25320 14399 25372 14408
rect 25320 14365 25329 14399
rect 25329 14365 25363 14399
rect 25363 14365 25372 14399
rect 25320 14356 25372 14365
rect 25780 14424 25832 14476
rect 25504 14399 25556 14408
rect 25504 14365 25513 14399
rect 25513 14365 25547 14399
rect 25547 14365 25556 14399
rect 25504 14356 25556 14365
rect 15752 14288 15804 14340
rect 27252 14492 27304 14544
rect 27988 14356 28040 14408
rect 28172 14492 28224 14544
rect 28908 14560 28960 14612
rect 29736 14492 29788 14544
rect 30012 14492 30064 14544
rect 30564 14492 30616 14544
rect 30932 14535 30984 14544
rect 30932 14501 30941 14535
rect 30941 14501 30975 14535
rect 30975 14501 30984 14535
rect 30932 14492 30984 14501
rect 32312 14492 32364 14544
rect 28356 14356 28408 14408
rect 30564 14356 30616 14408
rect 31576 14356 31628 14408
rect 31668 14399 31720 14408
rect 31668 14365 31677 14399
rect 31677 14365 31711 14399
rect 31711 14365 31720 14399
rect 31668 14356 31720 14365
rect 26240 14331 26292 14340
rect 26240 14297 26249 14331
rect 26249 14297 26283 14331
rect 26283 14297 26292 14331
rect 26240 14288 26292 14297
rect 27712 14288 27764 14340
rect 28632 14288 28684 14340
rect 29092 14288 29144 14340
rect 29736 14331 29788 14340
rect 29736 14297 29745 14331
rect 29745 14297 29779 14331
rect 29779 14297 29788 14331
rect 29736 14288 29788 14297
rect 31024 14288 31076 14340
rect 16396 14220 16448 14272
rect 16672 14220 16724 14272
rect 17132 14220 17184 14272
rect 18788 14220 18840 14272
rect 20720 14220 20772 14272
rect 22928 14220 22980 14272
rect 24952 14220 25004 14272
rect 27344 14220 27396 14272
rect 29644 14220 29696 14272
rect 31484 14220 31536 14272
rect 33140 14356 33192 14408
rect 37648 14492 37700 14544
rect 37924 14492 37976 14544
rect 34244 14356 34296 14408
rect 37280 14356 37332 14408
rect 37464 14356 37516 14408
rect 38016 14399 38068 14408
rect 38016 14365 38045 14399
rect 38045 14365 38068 14399
rect 38936 14399 38988 14408
rect 38016 14356 38068 14365
rect 38936 14365 38945 14399
rect 38945 14365 38979 14399
rect 38979 14365 38988 14399
rect 38936 14356 38988 14365
rect 68100 14399 68152 14408
rect 68100 14365 68109 14399
rect 68109 14365 68143 14399
rect 68143 14365 68152 14399
rect 68100 14356 68152 14365
rect 35900 14288 35952 14340
rect 36820 14331 36872 14340
rect 36820 14297 36829 14331
rect 36829 14297 36863 14331
rect 36863 14297 36872 14331
rect 36820 14288 36872 14297
rect 32956 14263 33008 14272
rect 32956 14229 32965 14263
rect 32965 14229 32999 14263
rect 32999 14229 33008 14263
rect 32956 14220 33008 14229
rect 34428 14220 34480 14272
rect 36636 14220 36688 14272
rect 37740 14220 37792 14272
rect 38844 14288 38896 14340
rect 38292 14263 38344 14272
rect 38292 14229 38301 14263
rect 38301 14229 38335 14263
rect 38335 14229 38344 14263
rect 38292 14220 38344 14229
rect 39120 14263 39172 14272
rect 39120 14229 39129 14263
rect 39129 14229 39163 14263
rect 39163 14229 39172 14263
rect 39120 14220 39172 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 4068 14059 4120 14068
rect 4068 14025 4077 14059
rect 4077 14025 4111 14059
rect 4111 14025 4120 14059
rect 4068 14016 4120 14025
rect 6644 14016 6696 14068
rect 7288 14016 7340 14068
rect 8116 14016 8168 14068
rect 9128 14016 9180 14068
rect 11152 14016 11204 14068
rect 11244 14016 11296 14068
rect 14188 14016 14240 14068
rect 3148 13948 3200 14000
rect 2780 13880 2832 13932
rect 4620 13948 4672 14000
rect 8392 13948 8444 14000
rect 4804 13923 4856 13932
rect 4804 13889 4813 13923
rect 4813 13889 4847 13923
rect 4847 13889 4856 13923
rect 4804 13880 4856 13889
rect 1768 13812 1820 13864
rect 6828 13880 6880 13932
rect 7748 13880 7800 13932
rect 9036 13880 9088 13932
rect 11796 13923 11848 13932
rect 3056 13676 3108 13728
rect 5908 13676 5960 13728
rect 8300 13744 8352 13796
rect 9036 13744 9088 13796
rect 11796 13889 11805 13923
rect 11805 13889 11839 13923
rect 11839 13889 11848 13923
rect 11796 13880 11848 13889
rect 11980 13923 12032 13932
rect 11980 13889 11989 13923
rect 11989 13889 12023 13923
rect 12023 13889 12032 13923
rect 11980 13880 12032 13889
rect 13268 13948 13320 14000
rect 12624 13880 12676 13932
rect 14096 13923 14148 13932
rect 14096 13889 14105 13923
rect 14105 13889 14139 13923
rect 14139 13889 14148 13923
rect 14096 13880 14148 13889
rect 15568 13923 15620 13932
rect 15568 13889 15577 13923
rect 15577 13889 15611 13923
rect 15611 13889 15620 13923
rect 15568 13880 15620 13889
rect 16120 13948 16172 14000
rect 16672 13923 16724 13932
rect 12716 13812 12768 13864
rect 11888 13744 11940 13796
rect 13636 13812 13688 13864
rect 15200 13812 15252 13864
rect 16672 13889 16681 13923
rect 16681 13889 16715 13923
rect 16715 13889 16724 13923
rect 16672 13880 16724 13889
rect 20168 14016 20220 14068
rect 18144 13880 18196 13932
rect 23388 13948 23440 14000
rect 25320 13948 25372 14000
rect 32496 14016 32548 14068
rect 32772 14016 32824 14068
rect 30564 13948 30616 14000
rect 19984 13880 20036 13932
rect 20168 13923 20220 13932
rect 20168 13889 20202 13923
rect 20202 13889 20220 13923
rect 22284 13923 22336 13932
rect 20168 13880 20220 13889
rect 22284 13889 22293 13923
rect 22293 13889 22327 13923
rect 22327 13889 22336 13923
rect 22284 13880 22336 13889
rect 22652 13880 22704 13932
rect 23572 13923 23624 13932
rect 23572 13889 23581 13923
rect 23581 13889 23615 13923
rect 23615 13889 23624 13923
rect 23572 13880 23624 13889
rect 24492 13880 24544 13932
rect 24952 13880 25004 13932
rect 16580 13812 16632 13864
rect 23664 13855 23716 13864
rect 7840 13676 7892 13728
rect 11796 13676 11848 13728
rect 16672 13719 16724 13728
rect 16672 13685 16681 13719
rect 16681 13685 16715 13719
rect 16715 13685 16724 13719
rect 16672 13676 16724 13685
rect 23664 13821 23673 13855
rect 23673 13821 23707 13855
rect 23707 13821 23716 13855
rect 23664 13812 23716 13821
rect 25228 13923 25280 13932
rect 25228 13889 25237 13923
rect 25237 13889 25271 13923
rect 25271 13889 25280 13923
rect 25228 13880 25280 13889
rect 27068 13923 27120 13932
rect 25320 13812 25372 13864
rect 27068 13889 27077 13923
rect 27077 13889 27111 13923
rect 27111 13889 27120 13923
rect 27068 13880 27120 13889
rect 27988 13923 28040 13932
rect 27988 13889 27997 13923
rect 27997 13889 28031 13923
rect 28031 13889 28040 13923
rect 27988 13880 28040 13889
rect 27896 13812 27948 13864
rect 28264 13880 28316 13932
rect 32128 13880 32180 13932
rect 34520 14016 34572 14068
rect 33140 13948 33192 14000
rect 34244 13948 34296 14000
rect 36452 14016 36504 14068
rect 37740 14059 37792 14068
rect 37740 14025 37749 14059
rect 37749 14025 37783 14059
rect 37783 14025 37792 14059
rect 37740 14016 37792 14025
rect 36728 13948 36780 14000
rect 38292 13948 38344 14000
rect 28632 13812 28684 13864
rect 29184 13812 29236 13864
rect 29644 13812 29696 13864
rect 17500 13676 17552 13728
rect 19432 13719 19484 13728
rect 19432 13685 19441 13719
rect 19441 13685 19475 13719
rect 19475 13685 19484 13719
rect 19432 13676 19484 13685
rect 20260 13676 20312 13728
rect 21272 13719 21324 13728
rect 21272 13685 21281 13719
rect 21281 13685 21315 13719
rect 21315 13685 21324 13719
rect 21272 13676 21324 13685
rect 24768 13719 24820 13728
rect 24768 13685 24777 13719
rect 24777 13685 24811 13719
rect 24811 13685 24820 13719
rect 24768 13676 24820 13685
rect 25504 13744 25556 13796
rect 25780 13744 25832 13796
rect 28080 13676 28132 13728
rect 29000 13676 29052 13728
rect 29828 13676 29880 13728
rect 32404 13719 32456 13728
rect 32404 13685 32413 13719
rect 32413 13685 32447 13719
rect 32447 13685 32456 13719
rect 32404 13676 32456 13685
rect 32864 13744 32916 13796
rect 35900 13880 35952 13932
rect 35992 13880 36044 13932
rect 36636 13923 36688 13932
rect 36636 13889 36645 13923
rect 36645 13889 36679 13923
rect 36679 13889 36688 13923
rect 36636 13880 36688 13889
rect 37372 13923 37424 13932
rect 37372 13889 37381 13923
rect 37381 13889 37415 13923
rect 37415 13889 37424 13923
rect 37372 13880 37424 13889
rect 41236 13880 41288 13932
rect 35532 13812 35584 13864
rect 33048 13676 33100 13728
rect 37832 13676 37884 13728
rect 38016 13676 38068 13728
rect 39120 13676 39172 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 65654 13574 65706 13626
rect 65718 13574 65770 13626
rect 65782 13574 65834 13626
rect 65846 13574 65898 13626
rect 65910 13574 65962 13626
rect 2872 13472 2924 13524
rect 3056 13472 3108 13524
rect 5264 13472 5316 13524
rect 8208 13472 8260 13524
rect 11796 13472 11848 13524
rect 14740 13472 14792 13524
rect 17500 13472 17552 13524
rect 3148 13336 3200 13388
rect 4620 13268 4672 13320
rect 5724 13268 5776 13320
rect 2228 13243 2280 13252
rect 2228 13209 2237 13243
rect 2237 13209 2271 13243
rect 2271 13209 2280 13243
rect 2228 13200 2280 13209
rect 2320 13200 2372 13252
rect 7104 13379 7156 13388
rect 7104 13345 7113 13379
rect 7113 13345 7147 13379
rect 7147 13345 7156 13379
rect 7104 13336 7156 13345
rect 7840 13336 7892 13388
rect 9680 13336 9732 13388
rect 6552 13268 6604 13320
rect 2136 13132 2188 13184
rect 5264 13132 5316 13184
rect 8576 13200 8628 13252
rect 8668 13200 8720 13252
rect 9404 13243 9456 13252
rect 9404 13209 9413 13243
rect 9413 13209 9447 13243
rect 9447 13209 9456 13243
rect 9404 13200 9456 13209
rect 8300 13175 8352 13184
rect 8300 13141 8309 13175
rect 8309 13141 8343 13175
rect 8343 13141 8352 13175
rect 8300 13132 8352 13141
rect 11152 13268 11204 13320
rect 15108 13404 15160 13456
rect 16764 13447 16816 13456
rect 16764 13413 16773 13447
rect 16773 13413 16807 13447
rect 16807 13413 16816 13447
rect 16764 13404 16816 13413
rect 15292 13379 15344 13388
rect 15292 13345 15301 13379
rect 15301 13345 15335 13379
rect 15335 13345 15344 13379
rect 15292 13336 15344 13345
rect 19340 13472 19392 13524
rect 26148 13472 26200 13524
rect 35992 13515 36044 13524
rect 19340 13336 19392 13388
rect 19892 13336 19944 13388
rect 23848 13336 23900 13388
rect 24308 13336 24360 13388
rect 24952 13336 25004 13388
rect 11888 13311 11940 13320
rect 11888 13277 11897 13311
rect 11897 13277 11931 13311
rect 11931 13277 11940 13311
rect 11888 13268 11940 13277
rect 14556 13268 14608 13320
rect 15200 13268 15252 13320
rect 11704 13243 11756 13252
rect 11704 13209 11713 13243
rect 11713 13209 11747 13243
rect 11747 13209 11756 13243
rect 11704 13200 11756 13209
rect 12072 13175 12124 13184
rect 12072 13141 12081 13175
rect 12081 13141 12115 13175
rect 12115 13141 12124 13175
rect 12072 13132 12124 13141
rect 13176 13200 13228 13252
rect 13820 13200 13872 13252
rect 16304 13243 16356 13252
rect 16304 13209 16313 13243
rect 16313 13209 16347 13243
rect 16347 13209 16356 13243
rect 16304 13200 16356 13209
rect 18696 13200 18748 13252
rect 20076 13268 20128 13320
rect 20720 13268 20772 13320
rect 24768 13268 24820 13320
rect 25320 13311 25372 13320
rect 25320 13277 25329 13311
rect 25329 13277 25363 13311
rect 25363 13277 25372 13311
rect 25320 13268 25372 13277
rect 26240 13311 26292 13320
rect 26240 13277 26249 13311
rect 26249 13277 26283 13311
rect 26283 13277 26292 13311
rect 26240 13268 26292 13277
rect 28724 13311 28776 13320
rect 28724 13277 28733 13311
rect 28733 13277 28767 13311
rect 28767 13277 28776 13311
rect 29000 13311 29052 13320
rect 28724 13268 28776 13277
rect 29000 13277 29009 13311
rect 29009 13277 29043 13311
rect 29043 13277 29052 13311
rect 29000 13268 29052 13277
rect 29092 13268 29144 13320
rect 30564 13447 30616 13456
rect 30564 13413 30573 13447
rect 30573 13413 30607 13447
rect 30607 13413 30616 13447
rect 30564 13404 30616 13413
rect 34704 13404 34756 13456
rect 35992 13481 36001 13515
rect 36001 13481 36035 13515
rect 36035 13481 36044 13515
rect 35992 13472 36044 13481
rect 37556 13472 37608 13524
rect 38292 13472 38344 13524
rect 32312 13336 32364 13388
rect 32772 13336 32824 13388
rect 31300 13268 31352 13320
rect 31944 13311 31996 13320
rect 31944 13277 31953 13311
rect 31953 13277 31987 13311
rect 31987 13277 31996 13311
rect 34428 13336 34480 13388
rect 38752 13404 38804 13456
rect 35348 13311 35400 13320
rect 31944 13268 31996 13277
rect 35348 13277 35357 13311
rect 35357 13277 35391 13311
rect 35391 13277 35400 13311
rect 35348 13268 35400 13277
rect 35532 13311 35584 13320
rect 35532 13277 35541 13311
rect 35541 13277 35575 13311
rect 35575 13277 35584 13311
rect 35532 13268 35584 13277
rect 36820 13336 36872 13388
rect 14832 13132 14884 13184
rect 19156 13132 19208 13184
rect 20720 13132 20772 13184
rect 22284 13132 22336 13184
rect 22560 13132 22612 13184
rect 26056 13200 26108 13252
rect 29184 13200 29236 13252
rect 29920 13243 29972 13252
rect 29920 13209 29929 13243
rect 29929 13209 29963 13243
rect 29963 13209 29972 13243
rect 29920 13200 29972 13209
rect 32404 13200 32456 13252
rect 33140 13200 33192 13252
rect 36912 13268 36964 13320
rect 37556 13268 37608 13320
rect 38016 13311 38068 13320
rect 38016 13277 38025 13311
rect 38025 13277 38059 13311
rect 38059 13277 38068 13311
rect 38016 13268 38068 13277
rect 35992 13200 36044 13252
rect 38292 13268 38344 13320
rect 38752 13268 38804 13320
rect 68100 13311 68152 13320
rect 68100 13277 68109 13311
rect 68109 13277 68143 13311
rect 68143 13277 68152 13311
rect 68100 13268 68152 13277
rect 26792 13132 26844 13184
rect 27252 13132 27304 13184
rect 28264 13132 28316 13184
rect 29552 13175 29604 13184
rect 29552 13141 29561 13175
rect 29561 13141 29595 13175
rect 29595 13141 29604 13175
rect 29552 13132 29604 13141
rect 32772 13175 32824 13184
rect 32772 13141 32781 13175
rect 32781 13141 32815 13175
rect 32815 13141 32824 13175
rect 32772 13132 32824 13141
rect 38108 13132 38160 13184
rect 38476 13175 38528 13184
rect 38476 13141 38485 13175
rect 38485 13141 38519 13175
rect 38519 13141 38528 13175
rect 38476 13132 38528 13141
rect 41236 13132 41288 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 2228 12928 2280 12980
rect 5264 12971 5316 12980
rect 3792 12860 3844 12912
rect 5264 12937 5273 12971
rect 5273 12937 5307 12971
rect 5307 12937 5316 12971
rect 5264 12928 5316 12937
rect 5816 12928 5868 12980
rect 6552 12928 6604 12980
rect 8576 12928 8628 12980
rect 9772 12928 9824 12980
rect 3148 12835 3200 12844
rect 3148 12801 3157 12835
rect 3157 12801 3191 12835
rect 3191 12801 3200 12835
rect 3148 12792 3200 12801
rect 3240 12792 3292 12844
rect 6644 12835 6696 12844
rect 6644 12801 6653 12835
rect 6653 12801 6687 12835
rect 6687 12801 6696 12835
rect 6644 12792 6696 12801
rect 8024 12792 8076 12844
rect 8208 12792 8260 12844
rect 2228 12724 2280 12776
rect 7472 12724 7524 12776
rect 7748 12724 7800 12776
rect 8392 12767 8444 12776
rect 8392 12733 8401 12767
rect 8401 12733 8435 12767
rect 8435 12733 8444 12767
rect 8392 12724 8444 12733
rect 10508 12903 10560 12912
rect 10508 12869 10517 12903
rect 10517 12869 10551 12903
rect 10551 12869 10560 12903
rect 11704 12903 11756 12912
rect 10508 12860 10560 12869
rect 11704 12869 11713 12903
rect 11713 12869 11747 12903
rect 11747 12869 11756 12903
rect 11704 12860 11756 12869
rect 10140 12792 10192 12844
rect 10416 12835 10468 12844
rect 10416 12801 10425 12835
rect 10425 12801 10459 12835
rect 10459 12801 10468 12835
rect 10416 12792 10468 12801
rect 10600 12835 10652 12844
rect 10600 12801 10609 12835
rect 10609 12801 10643 12835
rect 10643 12801 10652 12835
rect 10600 12792 10652 12801
rect 11520 12835 11572 12844
rect 11520 12801 11529 12835
rect 11529 12801 11563 12835
rect 11563 12801 11572 12835
rect 11520 12792 11572 12801
rect 11888 12835 11940 12844
rect 11888 12801 11897 12835
rect 11897 12801 11931 12835
rect 11931 12801 11940 12835
rect 16304 12928 16356 12980
rect 17960 12928 18012 12980
rect 18144 12928 18196 12980
rect 15200 12860 15252 12912
rect 11888 12792 11940 12801
rect 13820 12792 13872 12844
rect 14188 12792 14240 12844
rect 15384 12792 15436 12844
rect 15568 12792 15620 12844
rect 19248 12928 19300 12980
rect 20168 12928 20220 12980
rect 22100 12928 22152 12980
rect 23388 12928 23440 12980
rect 25228 12928 25280 12980
rect 26056 12971 26108 12980
rect 26056 12937 26065 12971
rect 26065 12937 26099 12971
rect 26099 12937 26108 12971
rect 26056 12928 26108 12937
rect 27160 12928 27212 12980
rect 27712 12928 27764 12980
rect 28908 12928 28960 12980
rect 38936 12928 38988 12980
rect 19524 12860 19576 12912
rect 9772 12699 9824 12708
rect 9772 12665 9781 12699
rect 9781 12665 9815 12699
rect 9815 12665 9824 12699
rect 9772 12656 9824 12665
rect 11520 12656 11572 12708
rect 12072 12699 12124 12708
rect 12072 12665 12081 12699
rect 12081 12665 12115 12699
rect 12115 12665 12124 12699
rect 12072 12656 12124 12665
rect 12808 12656 12860 12708
rect 16856 12724 16908 12776
rect 17500 12767 17552 12776
rect 17500 12733 17509 12767
rect 17509 12733 17543 12767
rect 17543 12733 17552 12767
rect 17500 12724 17552 12733
rect 18512 12835 18564 12844
rect 18512 12801 18521 12835
rect 18521 12801 18555 12835
rect 18555 12801 18564 12835
rect 18512 12792 18564 12801
rect 18696 12835 18748 12844
rect 18696 12801 18705 12835
rect 18705 12801 18739 12835
rect 18739 12801 18748 12835
rect 19432 12835 19484 12844
rect 18696 12792 18748 12801
rect 19432 12801 19441 12835
rect 19441 12801 19475 12835
rect 19475 12801 19484 12835
rect 19432 12792 19484 12801
rect 19892 12860 19944 12912
rect 19064 12724 19116 12776
rect 19800 12835 19852 12844
rect 19800 12801 19809 12835
rect 19809 12801 19843 12835
rect 19843 12801 19852 12835
rect 20260 12860 20312 12912
rect 22008 12903 22060 12912
rect 19800 12792 19852 12801
rect 21272 12792 21324 12844
rect 22008 12869 22017 12903
rect 22017 12869 22051 12903
rect 22051 12869 22060 12903
rect 22008 12860 22060 12869
rect 22560 12860 22612 12912
rect 25504 12860 25556 12912
rect 27252 12903 27304 12912
rect 14648 12656 14700 12708
rect 15108 12656 15160 12708
rect 15752 12699 15804 12708
rect 15752 12665 15761 12699
rect 15761 12665 15795 12699
rect 15795 12665 15804 12699
rect 15752 12656 15804 12665
rect 22100 12835 22152 12844
rect 22100 12801 22109 12835
rect 22109 12801 22143 12835
rect 22143 12801 22152 12835
rect 22100 12792 22152 12801
rect 22376 12792 22428 12844
rect 23480 12792 23532 12844
rect 23940 12835 23992 12844
rect 23940 12801 23949 12835
rect 23949 12801 23983 12835
rect 23983 12801 23992 12835
rect 23940 12792 23992 12801
rect 24308 12792 24360 12844
rect 25320 12792 25372 12844
rect 25596 12835 25648 12844
rect 25596 12801 25605 12835
rect 25605 12801 25639 12835
rect 25639 12801 25648 12835
rect 25596 12792 25648 12801
rect 27252 12869 27261 12903
rect 27261 12869 27295 12903
rect 27295 12869 27304 12903
rect 27252 12860 27304 12869
rect 27804 12860 27856 12912
rect 29460 12860 29512 12912
rect 32772 12860 32824 12912
rect 35440 12860 35492 12912
rect 35716 12903 35768 12912
rect 35716 12869 35725 12903
rect 35725 12869 35759 12903
rect 35759 12869 35768 12903
rect 35716 12860 35768 12869
rect 38476 12860 38528 12912
rect 26884 12792 26936 12844
rect 26976 12792 27028 12844
rect 23756 12767 23808 12776
rect 23756 12733 23765 12767
rect 23765 12733 23799 12767
rect 23799 12733 23808 12767
rect 23756 12724 23808 12733
rect 26332 12724 26384 12776
rect 27988 12792 28040 12844
rect 29092 12835 29144 12844
rect 29092 12801 29101 12835
rect 29101 12801 29135 12835
rect 29135 12801 29144 12835
rect 29092 12792 29144 12801
rect 31852 12792 31904 12844
rect 32128 12792 32180 12844
rect 35900 12835 35952 12844
rect 35900 12801 35909 12835
rect 35909 12801 35943 12835
rect 35943 12801 35952 12835
rect 37556 12835 37608 12844
rect 35900 12792 35952 12801
rect 35256 12724 35308 12776
rect 35440 12724 35492 12776
rect 37280 12767 37332 12776
rect 37280 12733 37289 12767
rect 37289 12733 37323 12767
rect 37323 12733 37332 12767
rect 37280 12724 37332 12733
rect 37556 12801 37565 12835
rect 37565 12801 37599 12835
rect 37599 12801 37608 12835
rect 37556 12792 37608 12801
rect 38660 12792 38712 12844
rect 38844 12792 38896 12844
rect 41236 12835 41288 12844
rect 41236 12801 41245 12835
rect 41245 12801 41279 12835
rect 41279 12801 41288 12835
rect 41236 12792 41288 12801
rect 10784 12631 10836 12640
rect 10784 12597 10793 12631
rect 10793 12597 10827 12631
rect 10827 12597 10836 12631
rect 10784 12588 10836 12597
rect 11060 12588 11112 12640
rect 11888 12588 11940 12640
rect 14188 12631 14240 12640
rect 14188 12597 14197 12631
rect 14197 12597 14231 12631
rect 14231 12597 14240 12631
rect 14188 12588 14240 12597
rect 17224 12631 17276 12640
rect 17224 12597 17233 12631
rect 17233 12597 17267 12631
rect 17267 12597 17276 12631
rect 17224 12588 17276 12597
rect 17868 12588 17920 12640
rect 25780 12588 25832 12640
rect 27620 12588 27672 12640
rect 30656 12588 30708 12640
rect 32680 12588 32732 12640
rect 34796 12588 34848 12640
rect 36544 12656 36596 12708
rect 35532 12631 35584 12640
rect 35532 12597 35541 12631
rect 35541 12597 35575 12631
rect 35575 12597 35584 12631
rect 35532 12588 35584 12597
rect 37832 12588 37884 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 65654 12486 65706 12538
rect 65718 12486 65770 12538
rect 65782 12486 65834 12538
rect 65846 12486 65898 12538
rect 65910 12486 65962 12538
rect 3240 12384 3292 12436
rect 5908 12384 5960 12436
rect 8208 12427 8260 12436
rect 8208 12393 8217 12427
rect 8217 12393 8251 12427
rect 8251 12393 8260 12427
rect 8208 12384 8260 12393
rect 11704 12384 11756 12436
rect 2320 12316 2372 12368
rect 2044 12248 2096 12300
rect 2136 12223 2188 12232
rect 2136 12189 2145 12223
rect 2145 12189 2179 12223
rect 2179 12189 2188 12223
rect 2136 12180 2188 12189
rect 2228 12223 2280 12232
rect 2228 12189 2237 12223
rect 2237 12189 2271 12223
rect 2271 12189 2280 12223
rect 2228 12180 2280 12189
rect 2504 12180 2556 12232
rect 4620 12180 4672 12232
rect 2780 12112 2832 12164
rect 6368 12180 6420 12232
rect 6644 12223 6696 12232
rect 6644 12189 6653 12223
rect 6653 12189 6687 12223
rect 6687 12189 6696 12223
rect 6644 12180 6696 12189
rect 7196 12180 7248 12232
rect 7748 12316 7800 12368
rect 9864 12316 9916 12368
rect 14280 12316 14332 12368
rect 8300 12248 8352 12300
rect 7932 12223 7984 12232
rect 7932 12189 7941 12223
rect 7941 12189 7975 12223
rect 7975 12189 7984 12223
rect 11060 12248 11112 12300
rect 7932 12180 7984 12189
rect 10600 12180 10652 12232
rect 12624 12223 12676 12232
rect 12624 12189 12626 12223
rect 12626 12189 12660 12223
rect 12660 12189 12676 12223
rect 12624 12180 12676 12189
rect 13084 12223 13136 12232
rect 13084 12189 13093 12223
rect 13093 12189 13127 12223
rect 13127 12189 13136 12223
rect 13084 12180 13136 12189
rect 14372 12223 14424 12232
rect 6184 12087 6236 12096
rect 6184 12053 6193 12087
rect 6193 12053 6227 12087
rect 6227 12053 6236 12087
rect 6184 12044 6236 12053
rect 6460 12044 6512 12096
rect 9036 12087 9088 12096
rect 9036 12053 9045 12087
rect 9045 12053 9079 12087
rect 9079 12053 9088 12087
rect 9036 12044 9088 12053
rect 10416 12112 10468 12164
rect 12900 12112 12952 12164
rect 14372 12189 14381 12223
rect 14381 12189 14415 12223
rect 14415 12189 14424 12223
rect 14372 12180 14424 12189
rect 14556 12180 14608 12232
rect 16212 12384 16264 12436
rect 18512 12384 18564 12436
rect 19800 12384 19852 12436
rect 20260 12384 20312 12436
rect 22192 12384 22244 12436
rect 15292 12316 15344 12368
rect 15476 12316 15528 12368
rect 24952 12384 25004 12436
rect 25596 12384 25648 12436
rect 25872 12384 25924 12436
rect 28264 12427 28316 12436
rect 23940 12316 23992 12368
rect 27620 12316 27672 12368
rect 28264 12393 28273 12427
rect 28273 12393 28307 12427
rect 28307 12393 28316 12427
rect 28264 12384 28316 12393
rect 33140 12427 33192 12436
rect 27896 12248 27948 12300
rect 28080 12291 28132 12300
rect 28080 12257 28089 12291
rect 28089 12257 28123 12291
rect 28123 12257 28132 12291
rect 28080 12248 28132 12257
rect 28172 12248 28224 12300
rect 16212 12223 16264 12232
rect 15384 12112 15436 12164
rect 10048 12087 10100 12096
rect 10048 12053 10057 12087
rect 10057 12053 10091 12087
rect 10091 12053 10100 12087
rect 10048 12044 10100 12053
rect 10968 12044 11020 12096
rect 13176 12044 13228 12096
rect 16212 12189 16221 12223
rect 16221 12189 16255 12223
rect 16255 12189 16264 12223
rect 16212 12180 16264 12189
rect 17868 12180 17920 12232
rect 19340 12180 19392 12232
rect 18144 12155 18196 12164
rect 18144 12121 18153 12155
rect 18153 12121 18187 12155
rect 18187 12121 18196 12155
rect 19800 12180 19852 12232
rect 20260 12180 20312 12232
rect 22376 12180 22428 12232
rect 23020 12180 23072 12232
rect 26976 12180 27028 12232
rect 27988 12223 28040 12232
rect 27988 12189 27997 12223
rect 27997 12189 28031 12223
rect 28031 12189 28040 12223
rect 27988 12180 28040 12189
rect 28264 12223 28316 12232
rect 28264 12189 28273 12223
rect 28273 12189 28307 12223
rect 28307 12189 28316 12223
rect 28264 12180 28316 12189
rect 29092 12180 29144 12232
rect 29920 12223 29972 12232
rect 29920 12189 29929 12223
rect 29929 12189 29963 12223
rect 29963 12189 29972 12223
rect 29920 12180 29972 12189
rect 30104 12223 30156 12232
rect 30104 12189 30113 12223
rect 30113 12189 30147 12223
rect 30147 12189 30156 12223
rect 30104 12180 30156 12189
rect 18144 12112 18196 12121
rect 21272 12112 21324 12164
rect 21548 12112 21600 12164
rect 21916 12155 21968 12164
rect 21916 12121 21925 12155
rect 21925 12121 21959 12155
rect 21959 12121 21968 12155
rect 21916 12112 21968 12121
rect 22284 12112 22336 12164
rect 24308 12112 24360 12164
rect 27620 12112 27672 12164
rect 32312 12180 32364 12232
rect 32680 12316 32732 12368
rect 32772 12316 32824 12368
rect 33140 12393 33149 12427
rect 33149 12393 33183 12427
rect 33183 12393 33192 12427
rect 33140 12384 33192 12393
rect 34520 12384 34572 12436
rect 35348 12384 35400 12436
rect 34796 12248 34848 12300
rect 35532 12223 35584 12232
rect 35532 12189 35541 12223
rect 35541 12189 35575 12223
rect 35575 12189 35584 12223
rect 37280 12248 37332 12300
rect 35532 12180 35584 12189
rect 37464 12180 37516 12232
rect 37556 12180 37608 12232
rect 37832 12223 37884 12232
rect 37832 12189 37841 12223
rect 37841 12189 37875 12223
rect 37875 12189 37884 12223
rect 37832 12180 37884 12189
rect 18972 12044 19024 12096
rect 19340 12044 19392 12096
rect 19524 12044 19576 12096
rect 20076 12087 20128 12096
rect 20076 12053 20085 12087
rect 20085 12053 20119 12087
rect 20119 12053 20128 12087
rect 20076 12044 20128 12053
rect 24768 12044 24820 12096
rect 25872 12044 25924 12096
rect 26240 12044 26292 12096
rect 26516 12044 26568 12096
rect 28448 12087 28500 12096
rect 28448 12053 28457 12087
rect 28457 12053 28491 12087
rect 28491 12053 28500 12087
rect 28448 12044 28500 12053
rect 29184 12044 29236 12096
rect 35992 12112 36044 12164
rect 37188 12112 37240 12164
rect 38016 12223 38068 12232
rect 38016 12189 38025 12223
rect 38025 12189 38059 12223
rect 38059 12189 38068 12223
rect 38016 12180 38068 12189
rect 38200 12180 38252 12232
rect 40500 12180 40552 12232
rect 41236 12223 41288 12232
rect 41236 12189 41245 12223
rect 41245 12189 41279 12223
rect 41279 12189 41288 12223
rect 41236 12180 41288 12189
rect 38108 12112 38160 12164
rect 33416 12044 33468 12096
rect 35072 12087 35124 12096
rect 35072 12053 35081 12087
rect 35081 12053 35115 12087
rect 35115 12053 35124 12087
rect 35072 12044 35124 12053
rect 38660 12044 38712 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 6644 11840 6696 11892
rect 13360 11840 13412 11892
rect 14188 11883 14240 11892
rect 14188 11849 14197 11883
rect 14197 11849 14231 11883
rect 14231 11849 14240 11883
rect 14188 11840 14240 11849
rect 5172 11772 5224 11824
rect 1768 11704 1820 11756
rect 2136 11747 2188 11756
rect 2136 11713 2145 11747
rect 2145 11713 2179 11747
rect 2179 11713 2188 11747
rect 2136 11704 2188 11713
rect 2228 11747 2280 11756
rect 2228 11713 2237 11747
rect 2237 11713 2271 11747
rect 2271 11713 2280 11747
rect 2228 11704 2280 11713
rect 2780 11704 2832 11756
rect 5816 11747 5868 11756
rect 5816 11713 5825 11747
rect 5825 11713 5859 11747
rect 5859 11713 5868 11747
rect 5816 11704 5868 11713
rect 6736 11747 6788 11756
rect 6736 11713 6745 11747
rect 6745 11713 6779 11747
rect 6779 11713 6788 11747
rect 6736 11704 6788 11713
rect 10416 11747 10468 11756
rect 10416 11713 10425 11747
rect 10425 11713 10459 11747
rect 10459 11713 10468 11747
rect 10416 11704 10468 11713
rect 11704 11747 11756 11756
rect 11704 11713 11713 11747
rect 11713 11713 11747 11747
rect 11747 11713 11756 11747
rect 11704 11704 11756 11713
rect 3148 11679 3200 11688
rect 3148 11645 3157 11679
rect 3157 11645 3191 11679
rect 3191 11645 3200 11679
rect 3148 11636 3200 11645
rect 6368 11636 6420 11688
rect 9496 11679 9548 11688
rect 9496 11645 9505 11679
rect 9505 11645 9539 11679
rect 9539 11645 9548 11679
rect 9496 11636 9548 11645
rect 11888 11747 11940 11756
rect 11888 11713 11897 11747
rect 11897 11713 11931 11747
rect 11931 11713 11940 11747
rect 11888 11704 11940 11713
rect 12900 11704 12952 11756
rect 13176 11636 13228 11688
rect 13728 11704 13780 11756
rect 15844 11815 15896 11824
rect 15844 11781 15853 11815
rect 15853 11781 15887 11815
rect 15887 11781 15896 11815
rect 15844 11772 15896 11781
rect 16396 11840 16448 11892
rect 21272 11883 21324 11892
rect 17868 11772 17920 11824
rect 19708 11772 19760 11824
rect 19800 11772 19852 11824
rect 21272 11849 21281 11883
rect 21281 11849 21315 11883
rect 21315 11849 21324 11883
rect 21272 11840 21324 11849
rect 22100 11840 22152 11892
rect 22192 11772 22244 11824
rect 25504 11840 25556 11892
rect 26792 11840 26844 11892
rect 27528 11840 27580 11892
rect 28172 11840 28224 11892
rect 25044 11772 25096 11824
rect 32128 11840 32180 11892
rect 32312 11840 32364 11892
rect 29460 11815 29512 11824
rect 18144 11747 18196 11756
rect 18144 11713 18153 11747
rect 18153 11713 18187 11747
rect 18187 11713 18196 11747
rect 18144 11704 18196 11713
rect 19892 11747 19944 11756
rect 19892 11713 19901 11747
rect 19901 11713 19935 11747
rect 19935 11713 19944 11747
rect 19892 11704 19944 11713
rect 12072 11611 12124 11620
rect 2504 11500 2556 11552
rect 12072 11577 12081 11611
rect 12081 11577 12115 11611
rect 12115 11577 12124 11611
rect 12072 11568 12124 11577
rect 7564 11500 7616 11552
rect 9496 11500 9548 11552
rect 13360 11500 13412 11552
rect 15844 11500 15896 11552
rect 18880 11636 18932 11688
rect 18972 11636 19024 11688
rect 21456 11704 21508 11756
rect 24216 11704 24268 11756
rect 24308 11747 24360 11756
rect 24308 11713 24317 11747
rect 24317 11713 24351 11747
rect 24351 11713 24360 11747
rect 25320 11747 25372 11756
rect 24308 11704 24360 11713
rect 25320 11713 25329 11747
rect 25329 11713 25363 11747
rect 25363 11713 25372 11747
rect 25320 11704 25372 11713
rect 25504 11747 25556 11756
rect 25504 11713 25513 11747
rect 25513 11713 25547 11747
rect 25547 11713 25556 11747
rect 25504 11704 25556 11713
rect 25688 11747 25740 11756
rect 25688 11713 25697 11747
rect 25697 11713 25731 11747
rect 25731 11713 25740 11747
rect 26976 11747 27028 11756
rect 25688 11704 25740 11713
rect 26976 11713 26985 11747
rect 26985 11713 27019 11747
rect 27019 11713 27028 11747
rect 26976 11704 27028 11713
rect 29460 11781 29469 11815
rect 29469 11781 29503 11815
rect 29503 11781 29512 11815
rect 29460 11772 29512 11781
rect 29920 11772 29972 11824
rect 27896 11704 27948 11756
rect 29092 11704 29144 11756
rect 29368 11747 29420 11756
rect 29368 11713 29377 11747
rect 29377 11713 29411 11747
rect 29411 11713 29420 11747
rect 29368 11704 29420 11713
rect 30472 11704 30524 11756
rect 31944 11704 31996 11756
rect 32496 11747 32548 11756
rect 32496 11713 32505 11747
rect 32505 11713 32539 11747
rect 32539 11713 32548 11747
rect 32496 11704 32548 11713
rect 32772 11772 32824 11824
rect 32680 11747 32732 11756
rect 32680 11713 32689 11747
rect 32689 11713 32723 11747
rect 32723 11713 32732 11747
rect 35716 11840 35768 11892
rect 35072 11772 35124 11824
rect 37372 11840 37424 11892
rect 32680 11704 32732 11713
rect 23848 11679 23900 11688
rect 23848 11645 23857 11679
rect 23857 11645 23891 11679
rect 23891 11645 23900 11679
rect 23848 11636 23900 11645
rect 26516 11636 26568 11688
rect 27068 11679 27120 11688
rect 27068 11645 27077 11679
rect 27077 11645 27111 11679
rect 27111 11645 27120 11679
rect 27068 11636 27120 11645
rect 28172 11611 28224 11620
rect 28172 11577 28181 11611
rect 28181 11577 28215 11611
rect 28215 11577 28224 11611
rect 28172 11568 28224 11577
rect 28264 11568 28316 11620
rect 37464 11747 37516 11756
rect 37464 11713 37473 11747
rect 37473 11713 37507 11747
rect 37507 11713 37516 11747
rect 37464 11704 37516 11713
rect 38016 11704 38068 11756
rect 37924 11636 37976 11688
rect 40500 11747 40552 11756
rect 40500 11713 40509 11747
rect 40509 11713 40543 11747
rect 40543 11713 40552 11747
rect 40500 11704 40552 11713
rect 67640 11611 67692 11620
rect 17040 11500 17092 11552
rect 18512 11543 18564 11552
rect 18512 11509 18521 11543
rect 18521 11509 18555 11543
rect 18555 11509 18564 11543
rect 18512 11500 18564 11509
rect 20168 11500 20220 11552
rect 21272 11500 21324 11552
rect 22376 11500 22428 11552
rect 25136 11500 25188 11552
rect 26608 11500 26660 11552
rect 27344 11500 27396 11552
rect 27804 11500 27856 11552
rect 28540 11500 28592 11552
rect 29092 11500 29144 11552
rect 30288 11500 30340 11552
rect 67640 11577 67649 11611
rect 67649 11577 67683 11611
rect 67683 11577 67692 11611
rect 67640 11568 67692 11577
rect 36912 11500 36964 11552
rect 37280 11500 37332 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 65654 11398 65706 11450
rect 65718 11398 65770 11450
rect 65782 11398 65834 11450
rect 65846 11398 65898 11450
rect 65910 11398 65962 11450
rect 2136 11296 2188 11348
rect 2780 11339 2832 11348
rect 2780 11305 2789 11339
rect 2789 11305 2823 11339
rect 2823 11305 2832 11339
rect 2780 11296 2832 11305
rect 5172 11339 5224 11348
rect 5172 11305 5181 11339
rect 5181 11305 5215 11339
rect 5215 11305 5224 11339
rect 5172 11296 5224 11305
rect 7932 11296 7984 11348
rect 13452 11296 13504 11348
rect 12440 11228 12492 11280
rect 16396 11296 16448 11348
rect 17868 11296 17920 11348
rect 18420 11339 18472 11348
rect 18420 11305 18429 11339
rect 18429 11305 18463 11339
rect 18463 11305 18472 11339
rect 18420 11296 18472 11305
rect 19800 11296 19852 11348
rect 22192 11296 22244 11348
rect 23940 11296 23992 11348
rect 24216 11296 24268 11348
rect 24860 11296 24912 11348
rect 25596 11296 25648 11348
rect 25688 11296 25740 11348
rect 26148 11296 26200 11348
rect 8392 11160 8444 11212
rect 19892 11228 19944 11280
rect 2504 11092 2556 11144
rect 3148 11092 3200 11144
rect 7564 11092 7616 11144
rect 2320 11067 2372 11076
rect 2320 11033 2329 11067
rect 2329 11033 2363 11067
rect 2363 11033 2372 11067
rect 2320 11024 2372 11033
rect 6184 11024 6236 11076
rect 7012 11024 7064 11076
rect 7748 11092 7800 11144
rect 7932 11135 7984 11144
rect 7932 11101 7941 11135
rect 7941 11101 7975 11135
rect 7975 11101 7984 11135
rect 7932 11092 7984 11101
rect 8760 11092 8812 11144
rect 13728 11092 13780 11144
rect 19616 11160 19668 11212
rect 19800 11160 19852 11212
rect 9036 10956 9088 11008
rect 10140 10956 10192 11008
rect 13268 11024 13320 11076
rect 15200 11024 15252 11076
rect 18052 11024 18104 11076
rect 19432 11092 19484 11144
rect 20076 11228 20128 11280
rect 20168 11228 20220 11280
rect 20720 11228 20772 11280
rect 21456 11160 21508 11212
rect 29276 11296 29328 11348
rect 32680 11296 32732 11348
rect 33968 11296 34020 11348
rect 34520 11296 34572 11348
rect 38016 11339 38068 11348
rect 38016 11305 38025 11339
rect 38025 11305 38059 11339
rect 38059 11305 38068 11339
rect 38016 11296 38068 11305
rect 29460 11228 29512 11280
rect 30656 11228 30708 11280
rect 21364 11135 21416 11144
rect 21364 11101 21373 11135
rect 21373 11101 21407 11135
rect 21407 11101 21416 11135
rect 21364 11092 21416 11101
rect 24768 11092 24820 11144
rect 25044 11135 25096 11144
rect 25044 11101 25053 11135
rect 25053 11101 25087 11135
rect 25087 11101 25096 11135
rect 25044 11092 25096 11101
rect 25136 11135 25188 11144
rect 25136 11101 25145 11135
rect 25145 11101 25179 11135
rect 25179 11101 25188 11135
rect 25136 11092 25188 11101
rect 25320 11135 25372 11144
rect 25320 11101 25329 11135
rect 25329 11101 25363 11135
rect 25363 11101 25372 11135
rect 26516 11135 26568 11144
rect 25320 11092 25372 11101
rect 26516 11101 26525 11135
rect 26525 11101 26559 11135
rect 26559 11101 26568 11135
rect 26516 11092 26568 11101
rect 26608 11092 26660 11144
rect 28540 11135 28592 11144
rect 19248 11024 19300 11076
rect 22376 11024 22428 11076
rect 28540 11101 28549 11135
rect 28549 11101 28583 11135
rect 28583 11101 28592 11135
rect 28540 11092 28592 11101
rect 28448 11024 28500 11076
rect 29368 11092 29420 11144
rect 30288 11160 30340 11212
rect 29920 11135 29972 11144
rect 29920 11101 29929 11135
rect 29929 11101 29963 11135
rect 29963 11101 29972 11135
rect 29920 11092 29972 11101
rect 30196 11092 30248 11144
rect 31852 11135 31904 11144
rect 31852 11101 31861 11135
rect 31861 11101 31895 11135
rect 31895 11101 31904 11135
rect 31852 11092 31904 11101
rect 32220 11160 32272 11212
rect 32496 11160 32548 11212
rect 34520 11160 34572 11212
rect 32588 11024 32640 11076
rect 34704 11067 34756 11076
rect 34704 11033 34713 11067
rect 34713 11033 34747 11067
rect 34747 11033 34756 11067
rect 34704 11024 34756 11033
rect 34980 11092 35032 11144
rect 35348 11024 35400 11076
rect 35808 11092 35860 11144
rect 37096 11092 37148 11144
rect 37280 11135 37332 11144
rect 37280 11101 37289 11135
rect 37289 11101 37323 11135
rect 37323 11101 37332 11135
rect 37280 11092 37332 11101
rect 38660 11092 38712 11144
rect 13820 10956 13872 11008
rect 14280 10956 14332 11008
rect 18236 10999 18288 11008
rect 18236 10965 18245 10999
rect 18245 10965 18279 10999
rect 18279 10965 18288 10999
rect 18236 10956 18288 10965
rect 20812 10999 20864 11008
rect 20812 10965 20821 10999
rect 20821 10965 20855 10999
rect 20855 10965 20864 10999
rect 20812 10956 20864 10965
rect 21088 10956 21140 11008
rect 33692 10956 33744 11008
rect 35532 10999 35584 11008
rect 35532 10965 35541 10999
rect 35541 10965 35575 10999
rect 35575 10965 35584 10999
rect 35532 10956 35584 10965
rect 37280 10956 37332 11008
rect 38384 10956 38436 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 4528 10795 4580 10804
rect 4528 10761 4537 10795
rect 4537 10761 4571 10795
rect 4571 10761 4580 10795
rect 7748 10795 7800 10804
rect 4528 10752 4580 10761
rect 1768 10659 1820 10668
rect 1768 10625 1777 10659
rect 1777 10625 1811 10659
rect 1811 10625 1820 10659
rect 1768 10616 1820 10625
rect 1860 10616 1912 10668
rect 2228 10684 2280 10736
rect 5816 10684 5868 10736
rect 7748 10761 7757 10795
rect 7757 10761 7791 10795
rect 7791 10761 7800 10795
rect 7748 10752 7800 10761
rect 2136 10659 2188 10668
rect 2136 10625 2145 10659
rect 2145 10625 2179 10659
rect 2179 10625 2188 10659
rect 3148 10659 3200 10668
rect 2136 10616 2188 10625
rect 3148 10625 3157 10659
rect 3157 10625 3191 10659
rect 3191 10625 3200 10659
rect 3148 10616 3200 10625
rect 3240 10616 3292 10668
rect 6828 10659 6880 10668
rect 6828 10625 6837 10659
rect 6837 10625 6871 10659
rect 6871 10625 6880 10659
rect 6828 10616 6880 10625
rect 7012 10659 7064 10668
rect 7012 10625 7021 10659
rect 7021 10625 7055 10659
rect 7055 10625 7064 10659
rect 7012 10616 7064 10625
rect 8760 10616 8812 10668
rect 10140 10659 10192 10668
rect 10140 10625 10149 10659
rect 10149 10625 10183 10659
rect 10183 10625 10192 10659
rect 10140 10616 10192 10625
rect 10416 10752 10468 10804
rect 12164 10752 12216 10804
rect 12532 10684 12584 10736
rect 15200 10752 15252 10804
rect 18420 10752 18472 10804
rect 19248 10752 19300 10804
rect 10600 10616 10652 10668
rect 11428 10616 11480 10668
rect 16396 10684 16448 10736
rect 17132 10684 17184 10736
rect 19800 10684 19852 10736
rect 23940 10752 23992 10804
rect 24768 10795 24820 10804
rect 24768 10761 24777 10795
rect 24777 10761 24811 10795
rect 24811 10761 24820 10795
rect 24768 10752 24820 10761
rect 25504 10752 25556 10804
rect 26240 10795 26292 10804
rect 26240 10761 26249 10795
rect 26249 10761 26283 10795
rect 26283 10761 26292 10795
rect 26240 10752 26292 10761
rect 26608 10752 26660 10804
rect 32680 10795 32732 10804
rect 32680 10761 32689 10795
rect 32689 10761 32723 10795
rect 32723 10761 32732 10795
rect 32680 10752 32732 10761
rect 34520 10795 34572 10804
rect 34520 10761 34529 10795
rect 34529 10761 34563 10795
rect 34563 10761 34572 10795
rect 34520 10752 34572 10761
rect 13912 10659 13964 10668
rect 13912 10625 13921 10659
rect 13921 10625 13955 10659
rect 13955 10625 13964 10659
rect 13912 10616 13964 10625
rect 14280 10659 14332 10668
rect 14280 10625 14289 10659
rect 14289 10625 14323 10659
rect 14323 10625 14332 10659
rect 14280 10616 14332 10625
rect 7932 10548 7984 10600
rect 14004 10591 14056 10600
rect 10692 10523 10744 10532
rect 10692 10489 10701 10523
rect 10701 10489 10735 10523
rect 10735 10489 10744 10523
rect 10692 10480 10744 10489
rect 2044 10412 2096 10464
rect 4528 10412 4580 10464
rect 6368 10455 6420 10464
rect 6368 10421 6377 10455
rect 6377 10421 6411 10455
rect 6411 10421 6420 10455
rect 6368 10412 6420 10421
rect 11520 10455 11572 10464
rect 11520 10421 11529 10455
rect 11529 10421 11563 10455
rect 11563 10421 11572 10455
rect 11520 10412 11572 10421
rect 14004 10557 14013 10591
rect 14013 10557 14047 10591
rect 14047 10557 14056 10591
rect 14004 10548 14056 10557
rect 14096 10591 14148 10600
rect 14096 10557 14105 10591
rect 14105 10557 14139 10591
rect 14139 10557 14148 10591
rect 14096 10548 14148 10557
rect 13268 10480 13320 10532
rect 16304 10616 16356 10668
rect 19984 10616 20036 10668
rect 21548 10616 21600 10668
rect 20812 10548 20864 10600
rect 30748 10684 30800 10736
rect 34980 10684 35032 10736
rect 22192 10659 22244 10668
rect 22192 10625 22201 10659
rect 22201 10625 22235 10659
rect 22235 10625 22244 10659
rect 22192 10616 22244 10625
rect 23020 10659 23072 10668
rect 23020 10625 23029 10659
rect 23029 10625 23063 10659
rect 23063 10625 23072 10659
rect 23020 10616 23072 10625
rect 22836 10591 22888 10600
rect 22836 10557 22845 10591
rect 22845 10557 22879 10591
rect 22879 10557 22888 10591
rect 22836 10548 22888 10557
rect 20536 10480 20588 10532
rect 13452 10412 13504 10464
rect 21088 10412 21140 10464
rect 23572 10412 23624 10464
rect 24124 10616 24176 10668
rect 25412 10616 25464 10668
rect 26148 10616 26200 10668
rect 28816 10659 28868 10668
rect 28816 10625 28825 10659
rect 28825 10625 28859 10659
rect 28859 10625 28868 10659
rect 28816 10616 28868 10625
rect 30656 10616 30708 10668
rect 32680 10616 32732 10668
rect 29460 10591 29512 10600
rect 29460 10557 29469 10591
rect 29469 10557 29503 10591
rect 29503 10557 29512 10591
rect 29460 10548 29512 10557
rect 33692 10659 33744 10668
rect 33692 10625 33701 10659
rect 33701 10625 33735 10659
rect 33735 10625 33744 10659
rect 33692 10616 33744 10625
rect 33876 10659 33928 10668
rect 33876 10625 33885 10659
rect 33885 10625 33919 10659
rect 33919 10625 33928 10659
rect 33876 10616 33928 10625
rect 34520 10616 34572 10668
rect 35440 10727 35492 10736
rect 35440 10693 35449 10727
rect 35449 10693 35483 10727
rect 35483 10693 35492 10727
rect 35440 10684 35492 10693
rect 35808 10616 35860 10668
rect 37464 10616 37516 10668
rect 38016 10659 38068 10668
rect 38016 10625 38025 10659
rect 38025 10625 38059 10659
rect 38059 10625 38068 10659
rect 38016 10616 38068 10625
rect 38200 10659 38252 10668
rect 38200 10625 38209 10659
rect 38209 10625 38243 10659
rect 38243 10625 38252 10659
rect 38200 10616 38252 10625
rect 34796 10548 34848 10600
rect 35532 10548 35584 10600
rect 37924 10548 37976 10600
rect 38384 10659 38436 10668
rect 38384 10625 38393 10659
rect 38393 10625 38427 10659
rect 38427 10625 38436 10659
rect 40500 10659 40552 10668
rect 38384 10616 38436 10625
rect 40500 10625 40509 10659
rect 40509 10625 40543 10659
rect 40543 10625 40552 10659
rect 40500 10616 40552 10625
rect 24860 10480 24912 10532
rect 28724 10480 28776 10532
rect 36820 10480 36872 10532
rect 26148 10412 26200 10464
rect 29552 10455 29604 10464
rect 29552 10421 29561 10455
rect 29561 10421 29595 10455
rect 29595 10421 29604 10455
rect 29552 10412 29604 10421
rect 33232 10455 33284 10464
rect 33232 10421 33241 10455
rect 33241 10421 33275 10455
rect 33275 10421 33284 10455
rect 33232 10412 33284 10421
rect 37372 10412 37424 10464
rect 37924 10412 37976 10464
rect 38108 10412 38160 10464
rect 67640 10455 67692 10464
rect 67640 10421 67649 10455
rect 67649 10421 67683 10455
rect 67683 10421 67692 10455
rect 67640 10412 67692 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 65654 10310 65706 10362
rect 65718 10310 65770 10362
rect 65782 10310 65834 10362
rect 65846 10310 65898 10362
rect 65910 10310 65962 10362
rect 1860 10251 1912 10260
rect 1860 10217 1869 10251
rect 1869 10217 1903 10251
rect 1903 10217 1912 10251
rect 1860 10208 1912 10217
rect 6828 10208 6880 10260
rect 2136 10140 2188 10192
rect 8760 10140 8812 10192
rect 2044 10047 2096 10056
rect 2044 10013 2053 10047
rect 2053 10013 2087 10047
rect 2087 10013 2096 10047
rect 2044 10004 2096 10013
rect 2412 10004 2464 10056
rect 3792 10047 3844 10056
rect 3792 10013 3801 10047
rect 3801 10013 3835 10047
rect 3835 10013 3844 10047
rect 3792 10004 3844 10013
rect 5816 10004 5868 10056
rect 7012 10004 7064 10056
rect 7656 10047 7708 10056
rect 7656 10013 7665 10047
rect 7665 10013 7699 10047
rect 7699 10013 7708 10047
rect 7656 10004 7708 10013
rect 7932 10072 7984 10124
rect 7840 10047 7892 10056
rect 7840 10013 7849 10047
rect 7849 10013 7883 10047
rect 7883 10013 7892 10047
rect 10968 10208 11020 10260
rect 11428 10251 11480 10260
rect 11428 10217 11437 10251
rect 11437 10217 11471 10251
rect 11471 10217 11480 10251
rect 11428 10208 11480 10217
rect 9680 10140 9732 10192
rect 14004 10208 14056 10260
rect 17500 10251 17552 10260
rect 17500 10217 17509 10251
rect 17509 10217 17543 10251
rect 17543 10217 17552 10251
rect 17500 10208 17552 10217
rect 18052 10251 18104 10260
rect 18052 10217 18061 10251
rect 18061 10217 18095 10251
rect 18095 10217 18104 10251
rect 18052 10208 18104 10217
rect 20168 10208 20220 10260
rect 20628 10208 20680 10260
rect 22836 10251 22888 10260
rect 12624 10140 12676 10192
rect 7840 10004 7892 10013
rect 9404 10004 9456 10056
rect 10140 10072 10192 10124
rect 10416 10072 10468 10124
rect 10692 10072 10744 10124
rect 18236 10140 18288 10192
rect 19524 10140 19576 10192
rect 22836 10217 22845 10251
rect 22845 10217 22879 10251
rect 22879 10217 22888 10251
rect 22836 10208 22888 10217
rect 24308 10208 24360 10260
rect 25412 10208 25464 10260
rect 28080 10208 28132 10260
rect 29184 10208 29236 10260
rect 31392 10208 31444 10260
rect 32588 10208 32640 10260
rect 34796 10251 34848 10260
rect 34796 10217 34805 10251
rect 34805 10217 34839 10251
rect 34839 10217 34848 10251
rect 34796 10208 34848 10217
rect 36912 10251 36964 10260
rect 36912 10217 36921 10251
rect 36921 10217 36955 10251
rect 36955 10217 36964 10251
rect 36912 10208 36964 10217
rect 38200 10208 38252 10260
rect 10600 10004 10652 10056
rect 11612 10047 11664 10056
rect 11612 10013 11621 10047
rect 11621 10013 11655 10047
rect 11655 10013 11664 10047
rect 11612 10004 11664 10013
rect 19708 10072 19760 10124
rect 28540 10183 28592 10192
rect 12164 10047 12216 10056
rect 3976 9979 4028 9988
rect 3976 9945 3985 9979
rect 3985 9945 4019 9979
rect 4019 9945 4028 9979
rect 3976 9936 4028 9945
rect 4160 9911 4212 9920
rect 4160 9877 4169 9911
rect 4169 9877 4203 9911
rect 4203 9877 4212 9911
rect 4160 9868 4212 9877
rect 5448 9868 5500 9920
rect 6920 9936 6972 9988
rect 12164 10013 12173 10047
rect 12173 10013 12207 10047
rect 12207 10013 12216 10047
rect 12164 10004 12216 10013
rect 14096 10004 14148 10056
rect 15844 10004 15896 10056
rect 16304 10047 16356 10056
rect 16304 10013 16313 10047
rect 16313 10013 16347 10047
rect 16347 10013 16356 10047
rect 16304 10004 16356 10013
rect 17592 10047 17644 10056
rect 17592 10013 17601 10047
rect 17601 10013 17635 10047
rect 17635 10013 17644 10047
rect 18328 10047 18380 10056
rect 17592 10004 17644 10013
rect 18328 10013 18337 10047
rect 18337 10013 18371 10047
rect 18371 10013 18380 10047
rect 18328 10004 18380 10013
rect 13820 9936 13872 9988
rect 18512 10047 18564 10056
rect 18512 10013 18521 10047
rect 18521 10013 18555 10047
rect 18555 10013 18564 10047
rect 18512 10004 18564 10013
rect 19432 10004 19484 10056
rect 20812 10072 20864 10124
rect 24860 10115 24912 10124
rect 24860 10081 24869 10115
rect 24869 10081 24903 10115
rect 24903 10081 24912 10115
rect 24860 10072 24912 10081
rect 25044 10072 25096 10124
rect 20168 10047 20220 10056
rect 20168 10013 20197 10047
rect 20197 10013 20220 10047
rect 20168 10004 20220 10013
rect 23572 10004 23624 10056
rect 24400 10004 24452 10056
rect 25320 10004 25372 10056
rect 26332 10047 26384 10056
rect 26332 10013 26341 10047
rect 26341 10013 26375 10047
rect 26375 10013 26384 10047
rect 26332 10004 26384 10013
rect 26608 10004 26660 10056
rect 28540 10149 28549 10183
rect 28549 10149 28583 10183
rect 28583 10149 28592 10183
rect 28540 10140 28592 10149
rect 7104 9868 7156 9920
rect 7840 9868 7892 9920
rect 8300 9868 8352 9920
rect 10968 9868 11020 9920
rect 11980 9868 12032 9920
rect 12716 9911 12768 9920
rect 12716 9877 12725 9911
rect 12725 9877 12759 9911
rect 12759 9877 12768 9911
rect 12716 9868 12768 9877
rect 13544 9911 13596 9920
rect 13544 9877 13553 9911
rect 13553 9877 13587 9911
rect 13587 9877 13596 9911
rect 13544 9868 13596 9877
rect 14188 9868 14240 9920
rect 15476 9868 15528 9920
rect 19340 9936 19392 9988
rect 19800 9868 19852 9920
rect 27528 10047 27580 10056
rect 27528 10013 27537 10047
rect 27537 10013 27571 10047
rect 27571 10013 27580 10047
rect 27528 10004 27580 10013
rect 28448 10004 28500 10056
rect 28724 10047 28776 10056
rect 28724 10013 28733 10047
rect 28733 10013 28767 10047
rect 28767 10013 28776 10047
rect 28724 10004 28776 10013
rect 28816 10047 28868 10056
rect 28816 10013 28825 10047
rect 28825 10013 28859 10047
rect 28859 10013 28868 10047
rect 28816 10004 28868 10013
rect 29000 10047 29052 10056
rect 29000 10013 29009 10047
rect 29009 10013 29043 10047
rect 29043 10013 29052 10047
rect 29000 10004 29052 10013
rect 27804 9936 27856 9988
rect 39028 10072 39080 10124
rect 33232 10004 33284 10056
rect 34520 10004 34572 10056
rect 35348 10004 35400 10056
rect 35716 10004 35768 10056
rect 35808 10004 35860 10056
rect 37096 10047 37148 10056
rect 34244 9936 34296 9988
rect 20076 9868 20128 9920
rect 20720 9868 20772 9920
rect 21088 9868 21140 9920
rect 26792 9911 26844 9920
rect 26792 9877 26801 9911
rect 26801 9877 26835 9911
rect 26835 9877 26844 9911
rect 26792 9868 26844 9877
rect 31392 9868 31444 9920
rect 34060 9868 34112 9920
rect 37096 10013 37105 10047
rect 37105 10013 37139 10047
rect 37139 10013 37148 10047
rect 37096 10004 37148 10013
rect 37004 9936 37056 9988
rect 37280 9979 37332 9988
rect 37280 9945 37289 9979
rect 37289 9945 37323 9979
rect 37323 9945 37332 9979
rect 37280 9936 37332 9945
rect 37740 10004 37792 10056
rect 38108 10047 38160 10056
rect 38108 10013 38117 10047
rect 38117 10013 38151 10047
rect 38151 10013 38160 10047
rect 38108 10004 38160 10013
rect 37924 9979 37976 9988
rect 37924 9945 37933 9979
rect 37933 9945 37967 9979
rect 37967 9945 37976 9979
rect 37924 9936 37976 9945
rect 37372 9868 37424 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 4160 9664 4212 9716
rect 1768 9528 1820 9580
rect 4620 9596 4672 9648
rect 5172 9673 5181 9686
rect 5181 9673 5215 9686
rect 5215 9673 5224 9686
rect 5172 9634 5224 9673
rect 7656 9664 7708 9716
rect 10968 9664 11020 9716
rect 14280 9664 14332 9716
rect 18788 9664 18840 9716
rect 19340 9664 19392 9716
rect 19524 9664 19576 9716
rect 20076 9664 20128 9716
rect 32680 9707 32732 9716
rect 32680 9673 32689 9707
rect 32689 9673 32723 9707
rect 32723 9673 32732 9707
rect 32680 9664 32732 9673
rect 5264 9596 5316 9648
rect 8300 9639 8352 9648
rect 2320 9392 2372 9444
rect 2412 9324 2464 9376
rect 2688 9367 2740 9376
rect 2688 9333 2697 9367
rect 2697 9333 2731 9367
rect 2731 9333 2740 9367
rect 2688 9324 2740 9333
rect 4068 9571 4120 9580
rect 4068 9537 4102 9571
rect 4102 9537 4120 9571
rect 4068 9528 4120 9537
rect 5816 9528 5868 9580
rect 7104 9324 7156 9376
rect 7564 9528 7616 9580
rect 8300 9605 8334 9639
rect 8334 9605 8352 9639
rect 8300 9596 8352 9605
rect 10416 9596 10468 9648
rect 8760 9528 8812 9580
rect 9956 9571 10008 9580
rect 9956 9537 9965 9571
rect 9965 9537 9999 9571
rect 9999 9537 10008 9571
rect 9956 9528 10008 9537
rect 10140 9571 10192 9580
rect 10140 9537 10149 9571
rect 10149 9537 10183 9571
rect 10183 9537 10192 9571
rect 10140 9528 10192 9537
rect 10600 9528 10652 9580
rect 12164 9571 12216 9580
rect 12164 9537 12173 9571
rect 12173 9537 12207 9571
rect 12207 9537 12216 9571
rect 12164 9528 12216 9537
rect 12624 9528 12676 9580
rect 15568 9571 15620 9580
rect 9864 9460 9916 9512
rect 12532 9503 12584 9512
rect 12532 9469 12541 9503
rect 12541 9469 12575 9503
rect 12575 9469 12584 9503
rect 12532 9460 12584 9469
rect 13360 9460 13412 9512
rect 14740 9503 14792 9512
rect 14740 9469 14749 9503
rect 14749 9469 14783 9503
rect 14783 9469 14792 9503
rect 14740 9460 14792 9469
rect 9404 9367 9456 9376
rect 9404 9333 9413 9367
rect 9413 9333 9447 9367
rect 9447 9333 9456 9367
rect 9404 9324 9456 9333
rect 10508 9367 10560 9376
rect 10508 9333 10517 9367
rect 10517 9333 10551 9367
rect 10551 9333 10560 9367
rect 10508 9324 10560 9333
rect 11520 9367 11572 9376
rect 11520 9333 11529 9367
rect 11529 9333 11563 9367
rect 11563 9333 11572 9367
rect 11520 9324 11572 9333
rect 13360 9367 13412 9376
rect 13360 9333 13369 9367
rect 13369 9333 13403 9367
rect 13403 9333 13412 9367
rect 13360 9324 13412 9333
rect 15568 9537 15577 9571
rect 15577 9537 15611 9571
rect 15611 9537 15620 9571
rect 15568 9528 15620 9537
rect 17224 9596 17276 9648
rect 18052 9596 18104 9648
rect 16396 9528 16448 9580
rect 17868 9571 17920 9580
rect 17868 9537 17877 9571
rect 17877 9537 17911 9571
rect 17911 9537 17920 9571
rect 17868 9528 17920 9537
rect 18420 9571 18472 9580
rect 15292 9460 15344 9512
rect 16948 9460 17000 9512
rect 18420 9537 18429 9571
rect 18429 9537 18463 9571
rect 18463 9537 18472 9571
rect 18420 9528 18472 9537
rect 20628 9596 20680 9648
rect 19524 9528 19576 9580
rect 22192 9596 22244 9648
rect 20076 9503 20128 9512
rect 20076 9469 20085 9503
rect 20085 9469 20119 9503
rect 20119 9469 20128 9503
rect 20076 9460 20128 9469
rect 20444 9460 20496 9512
rect 21548 9460 21600 9512
rect 22928 9528 22980 9580
rect 24308 9528 24360 9580
rect 24860 9596 24912 9648
rect 25412 9596 25464 9648
rect 26332 9596 26384 9648
rect 26516 9596 26568 9648
rect 24584 9571 24636 9580
rect 24584 9537 24593 9571
rect 24593 9537 24627 9571
rect 24627 9537 24636 9571
rect 24584 9528 24636 9537
rect 25320 9528 25372 9580
rect 27436 9528 27488 9580
rect 27988 9571 28040 9580
rect 27988 9537 27997 9571
rect 27997 9537 28031 9571
rect 28031 9537 28040 9571
rect 27988 9528 28040 9537
rect 28908 9571 28960 9580
rect 25596 9460 25648 9512
rect 28080 9503 28132 9512
rect 28080 9469 28089 9503
rect 28089 9469 28123 9503
rect 28123 9469 28132 9503
rect 28080 9460 28132 9469
rect 28908 9537 28917 9571
rect 28917 9537 28951 9571
rect 28951 9537 28960 9571
rect 28908 9528 28960 9537
rect 29000 9528 29052 9580
rect 29736 9528 29788 9580
rect 34244 9664 34296 9716
rect 34520 9596 34572 9648
rect 29552 9460 29604 9512
rect 18328 9392 18380 9444
rect 28172 9392 28224 9444
rect 28448 9435 28500 9444
rect 28448 9401 28457 9435
rect 28457 9401 28491 9435
rect 28491 9401 28500 9435
rect 28448 9392 28500 9401
rect 15384 9367 15436 9376
rect 15384 9333 15393 9367
rect 15393 9333 15427 9367
rect 15427 9333 15436 9367
rect 15384 9324 15436 9333
rect 17132 9367 17184 9376
rect 17132 9333 17141 9367
rect 17141 9333 17175 9367
rect 17175 9333 17184 9367
rect 17132 9324 17184 9333
rect 17316 9324 17368 9376
rect 17776 9367 17828 9376
rect 17776 9333 17785 9367
rect 17785 9333 17819 9367
rect 17819 9333 17828 9367
rect 17776 9324 17828 9333
rect 20076 9324 20128 9376
rect 24124 9367 24176 9376
rect 24124 9333 24133 9367
rect 24133 9333 24167 9367
rect 24167 9333 24176 9367
rect 24124 9324 24176 9333
rect 29276 9392 29328 9444
rect 33600 9571 33652 9580
rect 33600 9537 33609 9571
rect 33609 9537 33643 9571
rect 33643 9537 33652 9571
rect 33600 9528 33652 9537
rect 34428 9528 34480 9580
rect 34612 9528 34664 9580
rect 34704 9528 34756 9580
rect 35716 9571 35768 9580
rect 35716 9537 35725 9571
rect 35725 9537 35759 9571
rect 35759 9537 35768 9571
rect 35716 9528 35768 9537
rect 37556 9528 37608 9580
rect 38016 9571 38068 9580
rect 38016 9537 38025 9571
rect 38025 9537 38059 9571
rect 38059 9537 38068 9571
rect 38016 9528 38068 9537
rect 38384 9596 38436 9648
rect 39028 9571 39080 9580
rect 34520 9460 34572 9512
rect 35624 9460 35676 9512
rect 37188 9460 37240 9512
rect 39028 9537 39037 9571
rect 39037 9537 39071 9571
rect 39071 9537 39080 9571
rect 39028 9528 39080 9537
rect 35532 9392 35584 9444
rect 29092 9367 29144 9376
rect 29092 9333 29101 9367
rect 29101 9333 29135 9367
rect 29135 9333 29144 9367
rect 29092 9324 29144 9333
rect 29368 9367 29420 9376
rect 29368 9333 29377 9367
rect 29377 9333 29411 9367
rect 29411 9333 29420 9367
rect 29368 9324 29420 9333
rect 31116 9324 31168 9376
rect 35900 9324 35952 9376
rect 37188 9324 37240 9376
rect 37832 9324 37884 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 65654 9222 65706 9274
rect 65718 9222 65770 9274
rect 65782 9222 65834 9274
rect 65846 9222 65898 9274
rect 65910 9222 65962 9274
rect 1768 8916 1820 8968
rect 2320 8984 2372 9036
rect 3240 9120 3292 9172
rect 6920 9120 6972 9172
rect 9956 9120 10008 9172
rect 12532 9120 12584 9172
rect 15292 9120 15344 9172
rect 15568 9163 15620 9172
rect 15568 9129 15577 9163
rect 15577 9129 15611 9163
rect 15611 9129 15620 9163
rect 15568 9120 15620 9129
rect 17684 9163 17736 9172
rect 8116 9052 8168 9104
rect 9864 9052 9916 9104
rect 12072 9052 12124 9104
rect 11980 8984 12032 9036
rect 12440 9027 12492 9036
rect 12440 8993 12449 9027
rect 12449 8993 12483 9027
rect 12483 8993 12492 9027
rect 12440 8984 12492 8993
rect 4620 8916 4672 8968
rect 6368 8916 6420 8968
rect 10876 8916 10928 8968
rect 13636 9052 13688 9104
rect 15016 8984 15068 9036
rect 17684 9129 17693 9163
rect 17693 9129 17727 9163
rect 17727 9129 17736 9163
rect 17684 9120 17736 9129
rect 19524 9095 19576 9104
rect 19524 9061 19533 9095
rect 19533 9061 19567 9095
rect 19567 9061 19576 9095
rect 19524 9052 19576 9061
rect 20352 9052 20404 9104
rect 3792 8891 3844 8900
rect 3792 8857 3801 8891
rect 3801 8857 3835 8891
rect 3835 8857 3844 8891
rect 3792 8848 3844 8857
rect 5172 8848 5224 8900
rect 5448 8848 5500 8900
rect 10324 8848 10376 8900
rect 4068 8780 4120 8832
rect 5080 8780 5132 8832
rect 7288 8780 7340 8832
rect 8484 8780 8536 8832
rect 14280 8916 14332 8968
rect 14740 8916 14792 8968
rect 19984 8984 20036 9036
rect 15384 8916 15436 8968
rect 17776 8959 17828 8968
rect 17776 8925 17785 8959
rect 17785 8925 17819 8959
rect 17819 8925 17828 8959
rect 17776 8916 17828 8925
rect 16764 8848 16816 8900
rect 17224 8780 17276 8832
rect 17500 8823 17552 8832
rect 17500 8789 17509 8823
rect 17509 8789 17543 8823
rect 17543 8789 17552 8823
rect 17500 8780 17552 8789
rect 18144 8916 18196 8968
rect 18420 8959 18472 8968
rect 18420 8925 18429 8959
rect 18429 8925 18463 8959
rect 18463 8925 18472 8959
rect 18420 8916 18472 8925
rect 17960 8848 18012 8900
rect 19892 8916 19944 8968
rect 20536 8984 20588 9036
rect 24584 9120 24636 9172
rect 25320 9163 25372 9172
rect 25320 9129 25329 9163
rect 25329 9129 25363 9163
rect 25363 9129 25372 9163
rect 27436 9163 27488 9172
rect 25320 9120 25372 9129
rect 27436 9129 27445 9163
rect 27445 9129 27479 9163
rect 27479 9129 27488 9163
rect 27436 9120 27488 9129
rect 28908 9120 28960 9172
rect 30840 9163 30892 9172
rect 30840 9129 30849 9163
rect 30849 9129 30883 9163
rect 30883 9129 30892 9163
rect 30840 9120 30892 9129
rect 33600 9120 33652 9172
rect 34612 9120 34664 9172
rect 35256 9120 35308 9172
rect 38016 9163 38068 9172
rect 38016 9129 38025 9163
rect 38025 9129 38059 9163
rect 38059 9129 38068 9163
rect 38016 9120 38068 9129
rect 29736 9052 29788 9104
rect 21916 8916 21968 8968
rect 23388 8916 23440 8968
rect 20720 8848 20772 8900
rect 24124 8848 24176 8900
rect 24400 8891 24452 8900
rect 24400 8857 24409 8891
rect 24409 8857 24443 8891
rect 24443 8857 24452 8891
rect 24400 8848 24452 8857
rect 19892 8780 19944 8832
rect 20444 8780 20496 8832
rect 23204 8780 23256 8832
rect 25596 8848 25648 8900
rect 33324 8984 33376 9036
rect 34796 8984 34848 9036
rect 35716 8984 35768 9036
rect 26792 8916 26844 8968
rect 31024 8959 31076 8968
rect 31024 8925 31033 8959
rect 31033 8925 31067 8959
rect 31067 8925 31076 8959
rect 31024 8916 31076 8925
rect 31116 8959 31168 8968
rect 31116 8925 31125 8959
rect 31125 8925 31159 8959
rect 31159 8925 31168 8959
rect 31116 8916 31168 8925
rect 31208 8891 31260 8900
rect 31208 8857 31217 8891
rect 31217 8857 31251 8891
rect 31251 8857 31260 8891
rect 31208 8848 31260 8857
rect 31392 8959 31444 8968
rect 31392 8925 31401 8959
rect 31401 8925 31435 8959
rect 31435 8925 31444 8959
rect 31392 8916 31444 8925
rect 34612 8916 34664 8968
rect 35440 8916 35492 8968
rect 35624 8959 35676 8968
rect 35624 8925 35633 8959
rect 35633 8925 35667 8959
rect 35667 8925 35676 8959
rect 35624 8916 35676 8925
rect 37096 8984 37148 9036
rect 37004 8959 37056 8968
rect 37004 8925 37013 8959
rect 37013 8925 37047 8959
rect 37047 8925 37056 8959
rect 37004 8916 37056 8925
rect 37280 8916 37332 8968
rect 37832 8959 37884 8968
rect 37832 8925 37841 8959
rect 37841 8925 37875 8959
rect 37875 8925 37884 8959
rect 37832 8916 37884 8925
rect 32496 8780 32548 8832
rect 34520 8780 34572 8832
rect 38568 8848 38620 8900
rect 68100 8959 68152 8968
rect 68100 8925 68109 8959
rect 68109 8925 68143 8959
rect 68143 8925 68152 8959
rect 68100 8916 68152 8925
rect 41236 8848 41288 8900
rect 37464 8780 37516 8832
rect 38844 8823 38896 8832
rect 38844 8789 38853 8823
rect 38853 8789 38887 8823
rect 38887 8789 38896 8823
rect 38844 8780 38896 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 3148 8576 3200 8628
rect 3976 8619 4028 8628
rect 3976 8585 3985 8619
rect 3985 8585 4019 8619
rect 4019 8585 4028 8619
rect 3976 8576 4028 8585
rect 6736 8576 6788 8628
rect 2688 8508 2740 8560
rect 5724 8551 5776 8560
rect 5724 8517 5733 8551
rect 5733 8517 5767 8551
rect 5767 8517 5776 8551
rect 7380 8576 7432 8628
rect 12440 8576 12492 8628
rect 14280 8576 14332 8628
rect 19524 8576 19576 8628
rect 20076 8576 20128 8628
rect 5724 8508 5776 8517
rect 2044 8440 2096 8492
rect 3884 8440 3936 8492
rect 4804 8483 4856 8492
rect 4804 8449 4813 8483
rect 4813 8449 4847 8483
rect 4847 8449 4856 8483
rect 4804 8440 4856 8449
rect 3976 8372 4028 8424
rect 10416 8508 10468 8560
rect 7656 8440 7708 8492
rect 8208 8483 8260 8492
rect 7840 8372 7892 8424
rect 8208 8449 8217 8483
rect 8217 8449 8251 8483
rect 8251 8449 8260 8483
rect 8208 8440 8260 8449
rect 11152 8508 11204 8560
rect 12072 8483 12124 8492
rect 8668 8372 8720 8424
rect 7748 8304 7800 8356
rect 9680 8304 9732 8356
rect 11244 8372 11296 8424
rect 12072 8449 12081 8483
rect 12081 8449 12115 8483
rect 12115 8449 12124 8483
rect 12072 8440 12124 8449
rect 12164 8440 12216 8492
rect 19432 8508 19484 8560
rect 12532 8440 12584 8492
rect 16396 8440 16448 8492
rect 18052 8440 18104 8492
rect 19616 8440 19668 8492
rect 20260 8576 20312 8628
rect 23664 8576 23716 8628
rect 24308 8576 24360 8628
rect 28632 8576 28684 8628
rect 28816 8619 28868 8628
rect 28816 8585 28825 8619
rect 28825 8585 28859 8619
rect 28859 8585 28868 8619
rect 28816 8576 28868 8585
rect 32128 8619 32180 8628
rect 32128 8585 32137 8619
rect 32137 8585 32171 8619
rect 32171 8585 32180 8619
rect 32128 8576 32180 8585
rect 20812 8508 20864 8560
rect 23204 8551 23256 8560
rect 23204 8517 23213 8551
rect 23213 8517 23247 8551
rect 23247 8517 23256 8551
rect 23204 8508 23256 8517
rect 24860 8508 24912 8560
rect 27804 8508 27856 8560
rect 11980 8372 12032 8424
rect 13636 8415 13688 8424
rect 13636 8381 13645 8415
rect 13645 8381 13679 8415
rect 13679 8381 13688 8415
rect 13636 8372 13688 8381
rect 15292 8372 15344 8424
rect 15844 8372 15896 8424
rect 21916 8440 21968 8492
rect 23112 8483 23164 8492
rect 23112 8449 23121 8483
rect 23121 8449 23155 8483
rect 23155 8449 23164 8483
rect 23112 8440 23164 8449
rect 23572 8440 23624 8492
rect 31024 8508 31076 8560
rect 32496 8551 32548 8560
rect 26148 8483 26200 8492
rect 26148 8449 26157 8483
rect 26157 8449 26191 8483
rect 26191 8449 26200 8483
rect 26148 8440 26200 8449
rect 27160 8440 27212 8492
rect 28632 8483 28684 8492
rect 20444 8372 20496 8424
rect 25044 8372 25096 8424
rect 10784 8347 10836 8356
rect 10784 8313 10793 8347
rect 10793 8313 10827 8347
rect 10827 8313 10836 8347
rect 10784 8304 10836 8313
rect 11428 8304 11480 8356
rect 11888 8304 11940 8356
rect 12256 8304 12308 8356
rect 2964 8236 3016 8288
rect 5080 8236 5132 8288
rect 17040 8304 17092 8356
rect 17224 8304 17276 8356
rect 12808 8279 12860 8288
rect 12808 8245 12817 8279
rect 12817 8245 12851 8279
rect 12851 8245 12860 8279
rect 12808 8236 12860 8245
rect 13360 8236 13412 8288
rect 16212 8236 16264 8288
rect 17408 8236 17460 8288
rect 19340 8279 19392 8288
rect 19340 8245 19349 8279
rect 19349 8245 19383 8279
rect 19383 8245 19392 8279
rect 19984 8304 20036 8356
rect 20536 8304 20588 8356
rect 23572 8304 23624 8356
rect 26700 8372 26752 8424
rect 27712 8372 27764 8424
rect 28632 8449 28641 8483
rect 28641 8449 28675 8483
rect 28675 8449 28684 8483
rect 28632 8440 28684 8449
rect 29276 8483 29328 8492
rect 29276 8449 29285 8483
rect 29285 8449 29319 8483
rect 29319 8449 29328 8483
rect 29276 8440 29328 8449
rect 29460 8483 29512 8492
rect 29460 8449 29469 8483
rect 29469 8449 29503 8483
rect 29503 8449 29512 8483
rect 29460 8440 29512 8449
rect 32496 8517 32505 8551
rect 32505 8517 32539 8551
rect 32539 8517 32548 8551
rect 32496 8508 32548 8517
rect 32404 8483 32456 8492
rect 32404 8449 32413 8483
rect 32413 8449 32447 8483
rect 32447 8449 32456 8483
rect 32404 8440 32456 8449
rect 32588 8440 32640 8492
rect 39028 8576 39080 8628
rect 39856 8576 39908 8628
rect 34796 8508 34848 8560
rect 38752 8551 38804 8560
rect 38752 8517 38761 8551
rect 38761 8517 38795 8551
rect 38795 8517 38804 8551
rect 38752 8508 38804 8517
rect 34060 8483 34112 8492
rect 34060 8449 34069 8483
rect 34069 8449 34103 8483
rect 34103 8449 34112 8483
rect 34060 8440 34112 8449
rect 34428 8483 34480 8492
rect 28724 8372 28776 8424
rect 34428 8449 34437 8483
rect 34437 8449 34471 8483
rect 34471 8449 34480 8483
rect 34428 8440 34480 8449
rect 34704 8440 34756 8492
rect 35716 8483 35768 8492
rect 35716 8449 35725 8483
rect 35725 8449 35759 8483
rect 35759 8449 35768 8483
rect 35716 8440 35768 8449
rect 37096 8440 37148 8492
rect 34520 8372 34572 8424
rect 35992 8415 36044 8424
rect 35992 8381 36001 8415
rect 36001 8381 36035 8415
rect 36035 8381 36044 8415
rect 35992 8372 36044 8381
rect 37280 8415 37332 8424
rect 37280 8381 37289 8415
rect 37289 8381 37323 8415
rect 37323 8381 37332 8415
rect 37280 8372 37332 8381
rect 28172 8304 28224 8356
rect 31208 8304 31260 8356
rect 32680 8304 32732 8356
rect 33876 8347 33928 8356
rect 33876 8313 33885 8347
rect 33885 8313 33919 8347
rect 33919 8313 33928 8347
rect 33876 8304 33928 8313
rect 35900 8304 35952 8356
rect 38568 8304 38620 8356
rect 19340 8236 19392 8245
rect 20904 8236 20956 8288
rect 29736 8236 29788 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 65654 8134 65706 8186
rect 65718 8134 65770 8186
rect 65782 8134 65834 8186
rect 65846 8134 65898 8186
rect 65910 8134 65962 8186
rect 2596 8032 2648 8084
rect 2872 8032 2924 8084
rect 7748 8075 7800 8084
rect 7748 8041 7757 8075
rect 7757 8041 7791 8075
rect 7791 8041 7800 8075
rect 7748 8032 7800 8041
rect 2688 7964 2740 8016
rect 3332 7964 3384 8016
rect 6828 7964 6880 8016
rect 2320 7939 2372 7948
rect 2320 7905 2329 7939
rect 2329 7905 2363 7939
rect 2363 7905 2372 7939
rect 2320 7896 2372 7905
rect 2596 7828 2648 7880
rect 4620 7828 4672 7880
rect 5080 7871 5132 7880
rect 5080 7837 5114 7871
rect 5114 7837 5132 7871
rect 5080 7828 5132 7837
rect 4436 7760 4488 7812
rect 8208 7828 8260 7880
rect 12164 8032 12216 8084
rect 12532 7964 12584 8016
rect 12164 7896 12216 7948
rect 7656 7760 7708 7812
rect 9496 7828 9548 7880
rect 11796 7828 11848 7880
rect 12808 7828 12860 7880
rect 13452 7828 13504 7880
rect 16304 7828 16356 7880
rect 16396 7828 16448 7880
rect 17500 8032 17552 8084
rect 18052 8032 18104 8084
rect 21916 8075 21968 8084
rect 21916 8041 21925 8075
rect 21925 8041 21959 8075
rect 21959 8041 21968 8075
rect 21916 8032 21968 8041
rect 23756 8075 23808 8084
rect 23756 8041 23765 8075
rect 23765 8041 23799 8075
rect 23799 8041 23808 8075
rect 23756 8032 23808 8041
rect 27068 8032 27120 8084
rect 17868 7964 17920 8016
rect 25596 7964 25648 8016
rect 26056 7964 26108 8016
rect 17408 7871 17460 7880
rect 9680 7760 9732 7812
rect 1860 7692 1912 7744
rect 2872 7692 2924 7744
rect 3332 7692 3384 7744
rect 4896 7692 4948 7744
rect 7196 7692 7248 7744
rect 8392 7692 8444 7744
rect 11060 7735 11112 7744
rect 11060 7701 11069 7735
rect 11069 7701 11103 7735
rect 11103 7701 11112 7735
rect 11060 7692 11112 7701
rect 12440 7692 12492 7744
rect 14740 7692 14792 7744
rect 14924 7760 14976 7812
rect 16948 7760 17000 7812
rect 17408 7837 17417 7871
rect 17417 7837 17451 7871
rect 17451 7837 17460 7871
rect 17408 7828 17460 7837
rect 18328 7828 18380 7880
rect 20536 7871 20588 7880
rect 20536 7837 20545 7871
rect 20545 7837 20579 7871
rect 20579 7837 20588 7871
rect 20536 7828 20588 7837
rect 20812 7871 20864 7880
rect 20812 7837 20846 7871
rect 20846 7837 20864 7871
rect 20812 7828 20864 7837
rect 23480 7896 23532 7948
rect 24952 7896 25004 7948
rect 23572 7871 23624 7880
rect 23572 7837 23581 7871
rect 23581 7837 23615 7871
rect 23615 7837 23624 7871
rect 23572 7828 23624 7837
rect 24400 7871 24452 7880
rect 24400 7837 24409 7871
rect 24409 7837 24443 7871
rect 24443 7837 24452 7871
rect 24400 7828 24452 7837
rect 25780 7828 25832 7880
rect 25964 7828 26016 7880
rect 22652 7760 22704 7812
rect 23112 7760 23164 7812
rect 18512 7692 18564 7744
rect 20444 7692 20496 7744
rect 23664 7760 23716 7812
rect 27528 7896 27580 7948
rect 27804 7896 27856 7948
rect 28540 7896 28592 7948
rect 26700 7871 26752 7880
rect 26700 7837 26709 7871
rect 26709 7837 26743 7871
rect 26743 7837 26752 7871
rect 26700 7828 26752 7837
rect 29092 7828 29144 7880
rect 29736 7964 29788 8016
rect 29828 7964 29880 8016
rect 33784 7964 33836 8016
rect 33692 7896 33744 7948
rect 31208 7871 31260 7880
rect 31208 7837 31217 7871
rect 31217 7837 31251 7871
rect 31251 7837 31260 7871
rect 31208 7828 31260 7837
rect 32956 7828 33008 7880
rect 24860 7692 24912 7744
rect 25596 7692 25648 7744
rect 26240 7692 26292 7744
rect 30196 7735 30248 7744
rect 30196 7701 30205 7735
rect 30205 7701 30239 7735
rect 30239 7701 30248 7735
rect 30196 7692 30248 7701
rect 32588 7735 32640 7744
rect 32588 7701 32597 7735
rect 32597 7701 32631 7735
rect 32631 7701 32640 7735
rect 32588 7692 32640 7701
rect 33968 7865 34020 7874
rect 33968 7831 33977 7865
rect 33977 7831 34011 7865
rect 34011 7831 34020 7865
rect 33968 7822 34020 7831
rect 34244 7828 34296 7880
rect 34520 8032 34572 8084
rect 37280 8032 37332 8084
rect 41236 8075 41288 8084
rect 41236 8041 41245 8075
rect 41245 8041 41279 8075
rect 41279 8041 41288 8075
rect 41236 8032 41288 8041
rect 36176 7896 36228 7948
rect 37004 7896 37056 7948
rect 37372 7828 37424 7880
rect 37556 7828 37608 7880
rect 37924 7871 37976 7880
rect 37924 7837 37933 7871
rect 37933 7837 37967 7871
rect 37967 7837 37976 7871
rect 37924 7828 37976 7837
rect 38844 7896 38896 7948
rect 39856 7939 39908 7948
rect 39856 7905 39865 7939
rect 39865 7905 39899 7939
rect 39899 7905 39908 7939
rect 39856 7896 39908 7905
rect 35992 7760 36044 7812
rect 38292 7871 38344 7880
rect 38292 7837 38301 7871
rect 38301 7837 38335 7871
rect 38335 7837 38344 7871
rect 38292 7828 38344 7837
rect 68100 7871 68152 7880
rect 68100 7837 68109 7871
rect 68109 7837 68143 7871
rect 68143 7837 68152 7871
rect 68100 7828 68152 7837
rect 38384 7692 38436 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 4436 7488 4488 7540
rect 4804 7488 4856 7540
rect 2136 7395 2188 7404
rect 2136 7361 2145 7395
rect 2145 7361 2179 7395
rect 2179 7361 2188 7395
rect 2136 7352 2188 7361
rect 6368 7352 6420 7404
rect 10692 7488 10744 7540
rect 14924 7531 14976 7540
rect 2688 7284 2740 7336
rect 2964 7327 3016 7336
rect 2964 7293 2973 7327
rect 2973 7293 3007 7327
rect 3007 7293 3016 7327
rect 2964 7284 3016 7293
rect 6920 7284 6972 7336
rect 5816 7216 5868 7268
rect 6092 7148 6144 7200
rect 6460 7191 6512 7200
rect 6460 7157 6469 7191
rect 6469 7157 6503 7191
rect 6503 7157 6512 7191
rect 6460 7148 6512 7157
rect 8300 7420 8352 7472
rect 9220 7420 9272 7472
rect 12072 7420 12124 7472
rect 8392 7395 8444 7404
rect 7656 7284 7708 7336
rect 8392 7361 8401 7395
rect 8401 7361 8435 7395
rect 8435 7361 8444 7395
rect 8392 7352 8444 7361
rect 9680 7352 9732 7404
rect 10140 7352 10192 7404
rect 7196 7259 7248 7268
rect 7196 7225 7205 7259
rect 7205 7225 7239 7259
rect 7239 7225 7248 7259
rect 11060 7352 11112 7404
rect 11612 7284 11664 7336
rect 11980 7352 12032 7404
rect 13820 7420 13872 7472
rect 14004 7352 14056 7404
rect 14280 7395 14332 7404
rect 14280 7361 14289 7395
rect 14289 7361 14323 7395
rect 14323 7361 14332 7395
rect 14280 7352 14332 7361
rect 14924 7497 14933 7531
rect 14933 7497 14967 7531
rect 14967 7497 14976 7531
rect 14924 7488 14976 7497
rect 23572 7488 23624 7540
rect 24952 7488 25004 7540
rect 28080 7488 28132 7540
rect 29000 7488 29052 7540
rect 29460 7488 29512 7540
rect 33968 7488 34020 7540
rect 37372 7531 37424 7540
rect 37372 7497 37381 7531
rect 37381 7497 37415 7531
rect 37415 7497 37424 7531
rect 37372 7488 37424 7497
rect 38476 7488 38528 7540
rect 38752 7488 38804 7540
rect 15108 7420 15160 7472
rect 13544 7284 13596 7336
rect 14832 7352 14884 7404
rect 16672 7395 16724 7404
rect 16672 7361 16681 7395
rect 16681 7361 16715 7395
rect 16715 7361 16724 7395
rect 16672 7352 16724 7361
rect 19984 7420 20036 7472
rect 23664 7420 23716 7472
rect 27528 7463 27580 7472
rect 27528 7429 27537 7463
rect 27537 7429 27571 7463
rect 27571 7429 27580 7463
rect 27528 7420 27580 7429
rect 28448 7420 28500 7472
rect 29644 7420 29696 7472
rect 30196 7420 30248 7472
rect 32588 7420 32640 7472
rect 18512 7395 18564 7404
rect 18512 7361 18521 7395
rect 18521 7361 18555 7395
rect 18555 7361 18564 7395
rect 18512 7352 18564 7361
rect 21548 7352 21600 7404
rect 22652 7395 22704 7404
rect 22652 7361 22661 7395
rect 22661 7361 22695 7395
rect 22695 7361 22704 7395
rect 22652 7352 22704 7361
rect 24860 7352 24912 7404
rect 25320 7352 25372 7404
rect 18420 7284 18472 7336
rect 22376 7327 22428 7336
rect 22376 7293 22385 7327
rect 22385 7293 22419 7327
rect 22419 7293 22428 7327
rect 22376 7284 22428 7293
rect 25044 7284 25096 7336
rect 7196 7216 7248 7225
rect 19708 7216 19760 7268
rect 25780 7395 25832 7404
rect 25780 7361 25789 7395
rect 25789 7361 25823 7395
rect 25823 7361 25832 7395
rect 27344 7395 27396 7404
rect 25780 7352 25832 7361
rect 27344 7361 27353 7395
rect 27353 7361 27387 7395
rect 27387 7361 27396 7395
rect 27344 7352 27396 7361
rect 27712 7395 27764 7404
rect 27712 7361 27721 7395
rect 27721 7361 27755 7395
rect 27755 7361 27764 7395
rect 27712 7352 27764 7361
rect 27804 7352 27856 7404
rect 28540 7395 28592 7404
rect 28540 7361 28549 7395
rect 28549 7361 28583 7395
rect 28583 7361 28592 7395
rect 28540 7352 28592 7361
rect 29552 7352 29604 7404
rect 35900 7420 35952 7472
rect 36176 7463 36228 7472
rect 36176 7429 36185 7463
rect 36185 7429 36219 7463
rect 36219 7429 36228 7463
rect 36176 7420 36228 7429
rect 31208 7284 31260 7336
rect 31576 7284 31628 7336
rect 34428 7352 34480 7404
rect 36084 7395 36136 7404
rect 36084 7361 36093 7395
rect 36093 7361 36127 7395
rect 36127 7361 36136 7395
rect 36360 7395 36412 7404
rect 36084 7352 36136 7361
rect 36360 7361 36369 7395
rect 36369 7361 36403 7395
rect 36403 7361 36412 7395
rect 36360 7352 36412 7361
rect 37924 7395 37976 7404
rect 37924 7361 37933 7395
rect 37933 7361 37967 7395
rect 37967 7361 37976 7395
rect 37924 7352 37976 7361
rect 37096 7284 37148 7336
rect 38476 7352 38528 7404
rect 38384 7284 38436 7336
rect 38200 7216 38252 7268
rect 13912 7148 13964 7200
rect 14004 7148 14056 7200
rect 14740 7148 14792 7200
rect 16120 7191 16172 7200
rect 16120 7157 16129 7191
rect 16129 7157 16163 7191
rect 16163 7157 16172 7191
rect 16120 7148 16172 7157
rect 17500 7148 17552 7200
rect 20260 7148 20312 7200
rect 23848 7148 23900 7200
rect 25320 7148 25372 7200
rect 26332 7191 26384 7200
rect 26332 7157 26341 7191
rect 26341 7157 26375 7191
rect 26375 7157 26384 7191
rect 26332 7148 26384 7157
rect 26424 7148 26476 7200
rect 29092 7148 29144 7200
rect 34060 7148 34112 7200
rect 39948 7148 40000 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 65654 7046 65706 7098
rect 65718 7046 65770 7098
rect 65782 7046 65834 7098
rect 65846 7046 65898 7098
rect 65910 7046 65962 7098
rect 2136 6944 2188 6996
rect 6368 6987 6420 6996
rect 6368 6953 6377 6987
rect 6377 6953 6411 6987
rect 6411 6953 6420 6987
rect 6368 6944 6420 6953
rect 12808 6944 12860 6996
rect 13176 6944 13228 6996
rect 16672 6944 16724 6996
rect 34428 6944 34480 6996
rect 36360 6944 36412 6996
rect 38200 6987 38252 6996
rect 38200 6953 38209 6987
rect 38209 6953 38243 6987
rect 38243 6953 38252 6987
rect 38200 6944 38252 6953
rect 9864 6919 9916 6928
rect 9864 6885 9873 6919
rect 9873 6885 9907 6919
rect 9907 6885 9916 6919
rect 9864 6876 9916 6885
rect 1768 6808 1820 6860
rect 5908 6808 5960 6860
rect 6828 6851 6880 6860
rect 6828 6817 6837 6851
rect 6837 6817 6871 6851
rect 6871 6817 6880 6851
rect 6828 6808 6880 6817
rect 8116 6851 8168 6860
rect 1860 6783 1912 6792
rect 1860 6749 1869 6783
rect 1869 6749 1903 6783
rect 1903 6749 1912 6783
rect 1860 6740 1912 6749
rect 5080 6740 5132 6792
rect 6644 6740 6696 6792
rect 8116 6817 8125 6851
rect 8125 6817 8159 6851
rect 8159 6817 8168 6851
rect 8116 6808 8168 6817
rect 7656 6783 7708 6792
rect 7656 6749 7665 6783
rect 7665 6749 7699 6783
rect 7699 6749 7708 6783
rect 7656 6740 7708 6749
rect 7932 6783 7984 6792
rect 7932 6749 7941 6783
rect 7941 6749 7975 6783
rect 7975 6749 7984 6783
rect 7932 6740 7984 6749
rect 9772 6808 9824 6860
rect 10600 6851 10652 6860
rect 5540 6672 5592 6724
rect 6920 6672 6972 6724
rect 4620 6604 4672 6656
rect 6460 6604 6512 6656
rect 6828 6604 6880 6656
rect 7012 6604 7064 6656
rect 9220 6672 9272 6724
rect 9496 6783 9548 6792
rect 9496 6749 9505 6783
rect 9505 6749 9539 6783
rect 9539 6749 9548 6783
rect 9680 6783 9732 6792
rect 9496 6740 9548 6749
rect 9680 6749 9689 6783
rect 9689 6749 9723 6783
rect 9723 6749 9732 6783
rect 9680 6740 9732 6749
rect 10600 6817 10609 6851
rect 10609 6817 10643 6851
rect 10643 6817 10652 6851
rect 10600 6808 10652 6817
rect 25044 6876 25096 6928
rect 10692 6783 10744 6792
rect 10048 6672 10100 6724
rect 10692 6749 10701 6783
rect 10701 6749 10735 6783
rect 10735 6749 10744 6783
rect 10692 6740 10744 6749
rect 11704 6740 11756 6792
rect 11612 6672 11664 6724
rect 12624 6808 12676 6860
rect 15476 6808 15528 6860
rect 16304 6851 16356 6860
rect 16304 6817 16313 6851
rect 16313 6817 16347 6851
rect 16347 6817 16356 6851
rect 16304 6808 16356 6817
rect 20536 6851 20588 6860
rect 13360 6740 13412 6792
rect 13728 6740 13780 6792
rect 15752 6740 15804 6792
rect 16396 6740 16448 6792
rect 18512 6783 18564 6792
rect 18512 6749 18521 6783
rect 18521 6749 18555 6783
rect 18555 6749 18564 6783
rect 18512 6740 18564 6749
rect 19432 6783 19484 6792
rect 15936 6672 15988 6724
rect 16672 6672 16724 6724
rect 17224 6672 17276 6724
rect 19432 6749 19441 6783
rect 19441 6749 19475 6783
rect 19475 6749 19484 6783
rect 19432 6740 19484 6749
rect 11060 6647 11112 6656
rect 11060 6613 11069 6647
rect 11069 6613 11103 6647
rect 11103 6613 11112 6647
rect 11060 6604 11112 6613
rect 11152 6604 11204 6656
rect 12348 6604 12400 6656
rect 16856 6604 16908 6656
rect 19432 6604 19484 6656
rect 19800 6783 19852 6792
rect 19800 6749 19809 6783
rect 19809 6749 19843 6783
rect 19843 6749 19852 6783
rect 19800 6740 19852 6749
rect 20168 6740 20220 6792
rect 20536 6817 20545 6851
rect 20545 6817 20579 6851
rect 20579 6817 20588 6851
rect 20536 6808 20588 6817
rect 21548 6808 21600 6860
rect 22376 6783 22428 6792
rect 22376 6749 22385 6783
rect 22385 6749 22419 6783
rect 22419 6749 22428 6783
rect 22376 6740 22428 6749
rect 26240 6740 26292 6792
rect 26424 6783 26476 6792
rect 26424 6749 26433 6783
rect 26433 6749 26467 6783
rect 26467 6749 26476 6783
rect 26424 6740 26476 6749
rect 29828 6876 29880 6928
rect 30196 6876 30248 6928
rect 25596 6715 25648 6724
rect 25596 6681 25605 6715
rect 25605 6681 25639 6715
rect 25639 6681 25648 6715
rect 25596 6672 25648 6681
rect 26792 6783 26844 6792
rect 26792 6749 26801 6783
rect 26801 6749 26835 6783
rect 26835 6749 26844 6783
rect 26792 6740 26844 6749
rect 29276 6740 29328 6792
rect 29644 6740 29696 6792
rect 31576 6808 31628 6860
rect 37004 6808 37056 6860
rect 39856 6851 39908 6860
rect 32864 6740 32916 6792
rect 34612 6740 34664 6792
rect 37096 6740 37148 6792
rect 39856 6817 39865 6851
rect 39865 6817 39899 6851
rect 39899 6817 39908 6851
rect 39856 6808 39908 6817
rect 38568 6783 38620 6792
rect 19984 6604 20036 6656
rect 23756 6647 23808 6656
rect 23756 6613 23765 6647
rect 23765 6613 23799 6647
rect 23799 6613 23808 6647
rect 23756 6604 23808 6613
rect 25044 6647 25096 6656
rect 25044 6613 25053 6647
rect 25053 6613 25087 6647
rect 25087 6613 25096 6647
rect 27068 6647 27120 6656
rect 25044 6604 25096 6613
rect 27068 6613 27077 6647
rect 27077 6613 27111 6647
rect 27111 6613 27120 6647
rect 27068 6604 27120 6613
rect 28908 6647 28960 6656
rect 28908 6613 28917 6647
rect 28917 6613 28951 6647
rect 28951 6613 28960 6647
rect 28908 6604 28960 6613
rect 29552 6604 29604 6656
rect 32128 6672 32180 6724
rect 33600 6672 33652 6724
rect 35164 6672 35216 6724
rect 35808 6672 35860 6724
rect 38568 6749 38577 6783
rect 38577 6749 38611 6783
rect 38611 6749 38620 6783
rect 38568 6740 38620 6749
rect 39948 6740 40000 6792
rect 29920 6647 29972 6656
rect 29920 6613 29929 6647
rect 29929 6613 29963 6647
rect 29963 6613 29972 6647
rect 29920 6604 29972 6613
rect 34612 6604 34664 6656
rect 34704 6604 34756 6656
rect 36820 6604 36872 6656
rect 37648 6604 37700 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 2320 6332 2372 6384
rect 4068 6400 4120 6452
rect 5816 6400 5868 6452
rect 5908 6400 5960 6452
rect 7196 6400 7248 6452
rect 9220 6400 9272 6452
rect 9496 6400 9548 6452
rect 10692 6400 10744 6452
rect 16304 6400 16356 6452
rect 18052 6400 18104 6452
rect 19432 6400 19484 6452
rect 23664 6443 23716 6452
rect 23664 6409 23673 6443
rect 23673 6409 23707 6443
rect 23707 6409 23716 6443
rect 23664 6400 23716 6409
rect 25044 6400 25096 6452
rect 26792 6400 26844 6452
rect 2964 6332 3016 6384
rect 4620 6332 4672 6384
rect 5448 6332 5500 6384
rect 5724 6332 5776 6384
rect 6460 6332 6512 6384
rect 1768 6307 1820 6316
rect 1768 6273 1777 6307
rect 1777 6273 1811 6307
rect 1811 6273 1820 6307
rect 1768 6264 1820 6273
rect 1952 6060 2004 6112
rect 3056 6307 3108 6316
rect 3056 6273 3090 6307
rect 3090 6273 3108 6307
rect 3056 6264 3108 6273
rect 6920 6264 6972 6316
rect 8300 6332 8352 6384
rect 9128 6332 9180 6384
rect 11060 6332 11112 6384
rect 4068 6196 4120 6248
rect 6644 6196 6696 6248
rect 6828 6196 6880 6248
rect 7656 6196 7708 6248
rect 8024 6307 8076 6316
rect 8024 6273 8033 6307
rect 8033 6273 8067 6307
rect 8067 6273 8076 6307
rect 8024 6264 8076 6273
rect 9312 6264 9364 6316
rect 10140 6264 10192 6316
rect 12440 6332 12492 6384
rect 12624 6332 12676 6384
rect 17040 6375 17092 6384
rect 13452 6264 13504 6316
rect 15936 6307 15988 6316
rect 9588 6239 9640 6248
rect 9588 6205 9597 6239
rect 9597 6205 9631 6239
rect 9631 6205 9640 6239
rect 9588 6196 9640 6205
rect 9956 6196 10008 6248
rect 10876 6196 10928 6248
rect 15936 6273 15945 6307
rect 15945 6273 15979 6307
rect 15979 6273 15988 6307
rect 15936 6264 15988 6273
rect 17040 6341 17049 6375
rect 17049 6341 17083 6375
rect 17083 6341 17092 6375
rect 17040 6332 17092 6341
rect 19156 6264 19208 6316
rect 19984 6264 20036 6316
rect 20720 6307 20772 6316
rect 20720 6273 20729 6307
rect 20729 6273 20763 6307
rect 20763 6273 20772 6307
rect 20720 6264 20772 6273
rect 22100 6264 22152 6316
rect 23388 6332 23440 6384
rect 26332 6332 26384 6384
rect 27068 6332 27120 6384
rect 29644 6400 29696 6452
rect 33600 6443 33652 6452
rect 33600 6409 33609 6443
rect 33609 6409 33643 6443
rect 33643 6409 33652 6443
rect 33600 6400 33652 6409
rect 33692 6400 33744 6452
rect 35164 6443 35216 6452
rect 29736 6332 29788 6384
rect 35164 6409 35173 6443
rect 35173 6409 35207 6443
rect 35207 6409 35216 6443
rect 35164 6400 35216 6409
rect 35992 6400 36044 6452
rect 23848 6264 23900 6316
rect 27620 6264 27672 6316
rect 29092 6307 29144 6316
rect 29092 6273 29101 6307
rect 29101 6273 29135 6307
rect 29135 6273 29144 6307
rect 29092 6264 29144 6273
rect 10508 6128 10560 6180
rect 15660 6239 15712 6248
rect 15660 6205 15669 6239
rect 15669 6205 15703 6239
rect 15703 6205 15712 6239
rect 15660 6196 15712 6205
rect 17684 6196 17736 6248
rect 29000 6196 29052 6248
rect 15200 6128 15252 6180
rect 26240 6128 26292 6180
rect 29552 6264 29604 6316
rect 30472 6264 30524 6316
rect 33876 6307 33928 6316
rect 33876 6273 33885 6307
rect 33885 6273 33919 6307
rect 33919 6273 33928 6307
rect 33876 6264 33928 6273
rect 34060 6307 34112 6316
rect 34060 6273 34069 6307
rect 34069 6273 34103 6307
rect 34103 6273 34112 6307
rect 34060 6264 34112 6273
rect 34244 6307 34296 6316
rect 34244 6273 34253 6307
rect 34253 6273 34287 6307
rect 34287 6273 34296 6307
rect 34244 6264 34296 6273
rect 34612 6264 34664 6316
rect 35440 6307 35492 6316
rect 35440 6273 35449 6307
rect 35449 6273 35483 6307
rect 35483 6273 35492 6307
rect 35440 6264 35492 6273
rect 36360 6332 36412 6384
rect 38568 6400 38620 6452
rect 37648 6332 37700 6384
rect 38660 6332 38712 6384
rect 30196 6196 30248 6248
rect 31576 6239 31628 6248
rect 31576 6205 31585 6239
rect 31585 6205 31619 6239
rect 31619 6205 31628 6239
rect 31576 6196 31628 6205
rect 29276 6128 29328 6180
rect 30564 6128 30616 6180
rect 37372 6264 37424 6316
rect 38108 6307 38160 6316
rect 38108 6273 38117 6307
rect 38117 6273 38151 6307
rect 38151 6273 38160 6307
rect 38108 6264 38160 6273
rect 37188 6128 37240 6180
rect 38476 6307 38528 6316
rect 38476 6273 38485 6307
rect 38485 6273 38519 6307
rect 38519 6273 38528 6307
rect 38476 6264 38528 6273
rect 67640 6171 67692 6180
rect 67640 6137 67649 6171
rect 67649 6137 67683 6171
rect 67683 6137 67692 6171
rect 67640 6128 67692 6137
rect 8116 6060 8168 6112
rect 10600 6060 10652 6112
rect 11336 6060 11388 6112
rect 11704 6060 11756 6112
rect 14556 6060 14608 6112
rect 20076 6103 20128 6112
rect 20076 6069 20085 6103
rect 20085 6069 20119 6103
rect 20119 6069 20128 6103
rect 20076 6060 20128 6069
rect 23020 6060 23072 6112
rect 28264 6060 28316 6112
rect 30288 6060 30340 6112
rect 30932 6060 30984 6112
rect 38752 6103 38804 6112
rect 38752 6069 38761 6103
rect 38761 6069 38795 6103
rect 38795 6069 38804 6103
rect 38752 6060 38804 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 65654 5958 65706 6010
rect 65718 5958 65770 6010
rect 65782 5958 65834 6010
rect 65846 5958 65898 6010
rect 65910 5958 65962 6010
rect 3056 5856 3108 5908
rect 3240 5899 3292 5908
rect 3240 5865 3249 5899
rect 3249 5865 3283 5899
rect 3283 5865 3292 5899
rect 3240 5856 3292 5865
rect 5540 5856 5592 5908
rect 6736 5856 6788 5908
rect 9588 5856 9640 5908
rect 15660 5899 15712 5908
rect 5264 5788 5316 5840
rect 9220 5788 9272 5840
rect 13636 5788 13688 5840
rect 13820 5788 13872 5840
rect 8208 5720 8260 5772
rect 9864 5720 9916 5772
rect 15660 5865 15669 5899
rect 15669 5865 15703 5899
rect 15703 5865 15712 5899
rect 15660 5856 15712 5865
rect 16672 5899 16724 5908
rect 16672 5865 16681 5899
rect 16681 5865 16715 5899
rect 16715 5865 16724 5899
rect 16672 5856 16724 5865
rect 17868 5899 17920 5908
rect 17868 5865 17877 5899
rect 17877 5865 17911 5899
rect 17911 5865 17920 5899
rect 17868 5856 17920 5865
rect 18880 5856 18932 5908
rect 23480 5899 23532 5908
rect 17776 5788 17828 5840
rect 23480 5865 23489 5899
rect 23489 5865 23523 5899
rect 23523 5865 23532 5899
rect 23480 5856 23532 5865
rect 26332 5856 26384 5908
rect 28908 5856 28960 5908
rect 29276 5856 29328 5908
rect 30472 5899 30524 5908
rect 30472 5865 30481 5899
rect 30481 5865 30515 5899
rect 30515 5865 30524 5899
rect 30472 5856 30524 5865
rect 35440 5856 35492 5908
rect 35992 5899 36044 5908
rect 35992 5865 36001 5899
rect 36001 5865 36035 5899
rect 36035 5865 36044 5899
rect 35992 5856 36044 5865
rect 38476 5856 38528 5908
rect 26424 5788 26476 5840
rect 30932 5831 30984 5840
rect 30932 5797 30941 5831
rect 30941 5797 30975 5831
rect 30975 5797 30984 5831
rect 30932 5788 30984 5797
rect 1952 5695 2004 5704
rect 1952 5661 1961 5695
rect 1961 5661 1995 5695
rect 1995 5661 2004 5695
rect 1952 5652 2004 5661
rect 5816 5652 5868 5704
rect 7748 5652 7800 5704
rect 7840 5695 7892 5704
rect 7840 5661 7849 5695
rect 7849 5661 7883 5695
rect 7883 5661 7892 5695
rect 7840 5652 7892 5661
rect 3792 5559 3844 5568
rect 3792 5525 3801 5559
rect 3801 5525 3835 5559
rect 3835 5525 3844 5559
rect 3792 5516 3844 5525
rect 6368 5516 6420 5568
rect 6460 5516 6512 5568
rect 7196 5584 7248 5636
rect 9312 5652 9364 5704
rect 13176 5652 13228 5704
rect 14188 5652 14240 5704
rect 15384 5652 15436 5704
rect 9956 5627 10008 5636
rect 9956 5593 9965 5627
rect 9965 5593 9999 5627
rect 9999 5593 10008 5627
rect 9956 5584 10008 5593
rect 11888 5584 11940 5636
rect 16672 5652 16724 5704
rect 16856 5695 16908 5704
rect 16856 5661 16865 5695
rect 16865 5661 16899 5695
rect 16899 5661 16908 5695
rect 16856 5652 16908 5661
rect 17592 5720 17644 5772
rect 6736 5559 6788 5568
rect 6736 5525 6745 5559
rect 6745 5525 6779 5559
rect 6779 5525 6788 5559
rect 6736 5516 6788 5525
rect 7564 5516 7616 5568
rect 7932 5516 7984 5568
rect 16948 5584 17000 5636
rect 17040 5584 17092 5636
rect 17316 5652 17368 5704
rect 17684 5652 17736 5704
rect 19432 5720 19484 5772
rect 19616 5695 19668 5704
rect 19616 5661 19625 5695
rect 19625 5661 19659 5695
rect 19659 5661 19668 5695
rect 20260 5720 20312 5772
rect 19616 5652 19668 5661
rect 20168 5652 20220 5704
rect 22100 5763 22152 5772
rect 22100 5729 22109 5763
rect 22109 5729 22143 5763
rect 22143 5729 22152 5763
rect 22100 5720 22152 5729
rect 37188 5720 37240 5772
rect 23388 5652 23440 5704
rect 24676 5652 24728 5704
rect 28448 5652 28500 5704
rect 29092 5652 29144 5704
rect 29920 5652 29972 5704
rect 30104 5695 30156 5704
rect 30104 5661 30113 5695
rect 30113 5661 30147 5695
rect 30147 5661 30156 5695
rect 30104 5652 30156 5661
rect 30288 5652 30340 5704
rect 12348 5516 12400 5568
rect 12624 5516 12676 5568
rect 13544 5559 13596 5568
rect 13544 5525 13553 5559
rect 13553 5525 13587 5559
rect 13587 5525 13596 5559
rect 13544 5516 13596 5525
rect 14372 5516 14424 5568
rect 15936 5516 15988 5568
rect 17132 5516 17184 5568
rect 17316 5516 17368 5568
rect 19156 5516 19208 5568
rect 23296 5584 23348 5636
rect 25044 5627 25096 5636
rect 20260 5516 20312 5568
rect 23020 5516 23072 5568
rect 25044 5593 25053 5627
rect 25053 5593 25087 5627
rect 25087 5593 25096 5627
rect 25044 5584 25096 5593
rect 25596 5627 25648 5636
rect 25596 5593 25605 5627
rect 25605 5593 25639 5627
rect 25639 5593 25648 5627
rect 25596 5584 25648 5593
rect 26424 5627 26476 5636
rect 26424 5593 26433 5627
rect 26433 5593 26467 5627
rect 26467 5593 26476 5627
rect 26424 5584 26476 5593
rect 27160 5584 27212 5636
rect 29184 5584 29236 5636
rect 24768 5516 24820 5568
rect 27620 5516 27672 5568
rect 35532 5695 35584 5704
rect 35532 5661 35541 5695
rect 35541 5661 35575 5695
rect 35575 5661 35584 5695
rect 35532 5652 35584 5661
rect 36452 5652 36504 5704
rect 37280 5695 37332 5704
rect 31576 5584 31628 5636
rect 37280 5661 37289 5695
rect 37289 5661 37323 5695
rect 37323 5661 37332 5695
rect 37280 5652 37332 5661
rect 38292 5720 38344 5772
rect 38108 5584 38160 5636
rect 34704 5516 34756 5568
rect 37372 5516 37424 5568
rect 37740 5559 37792 5568
rect 37740 5525 37749 5559
rect 37749 5525 37783 5559
rect 37783 5525 37792 5559
rect 37740 5516 37792 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 8116 5355 8168 5364
rect 6828 5287 6880 5296
rect 6828 5253 6837 5287
rect 6837 5253 6871 5287
rect 6871 5253 6880 5287
rect 6828 5244 6880 5253
rect 2228 5219 2280 5228
rect 2228 5185 2237 5219
rect 2237 5185 2271 5219
rect 2271 5185 2280 5219
rect 2228 5176 2280 5185
rect 5540 5108 5592 5160
rect 8116 5321 8125 5355
rect 8125 5321 8159 5355
rect 8159 5321 8168 5355
rect 8116 5312 8168 5321
rect 9496 5355 9548 5364
rect 9496 5321 9505 5355
rect 9505 5321 9539 5355
rect 9539 5321 9548 5355
rect 9496 5312 9548 5321
rect 11244 5312 11296 5364
rect 13084 5312 13136 5364
rect 8852 5244 8904 5296
rect 7656 5219 7708 5228
rect 7656 5185 7665 5219
rect 7665 5185 7699 5219
rect 7699 5185 7708 5219
rect 7656 5176 7708 5185
rect 7932 5219 7984 5228
rect 7932 5185 7941 5219
rect 7941 5185 7975 5219
rect 7975 5185 7984 5219
rect 7932 5176 7984 5185
rect 9496 5219 9548 5228
rect 9496 5185 9505 5219
rect 9505 5185 9539 5219
rect 9539 5185 9548 5219
rect 9496 5176 9548 5185
rect 9772 5219 9824 5228
rect 9772 5185 9781 5219
rect 9781 5185 9815 5219
rect 9815 5185 9824 5219
rect 9772 5176 9824 5185
rect 10048 5219 10100 5228
rect 10048 5185 10057 5219
rect 10057 5185 10091 5219
rect 10091 5185 10100 5219
rect 10048 5176 10100 5185
rect 6920 5151 6972 5160
rect 2964 4972 3016 5024
rect 4712 4972 4764 5024
rect 6920 5117 6929 5151
rect 6929 5117 6963 5151
rect 6963 5117 6972 5151
rect 6920 5108 6972 5117
rect 7472 5108 7524 5160
rect 11060 5244 11112 5296
rect 10968 5219 11020 5228
rect 10968 5185 10977 5219
rect 10977 5185 11011 5219
rect 11011 5185 11020 5219
rect 10968 5176 11020 5185
rect 13268 5244 13320 5296
rect 14648 5312 14700 5364
rect 17132 5355 17184 5364
rect 17132 5321 17141 5355
rect 17141 5321 17175 5355
rect 17175 5321 17184 5355
rect 17132 5312 17184 5321
rect 18236 5312 18288 5364
rect 23296 5355 23348 5364
rect 23296 5321 23305 5355
rect 23305 5321 23339 5355
rect 23339 5321 23348 5355
rect 23296 5312 23348 5321
rect 28448 5312 28500 5364
rect 32864 5312 32916 5364
rect 34612 5312 34664 5364
rect 37280 5312 37332 5364
rect 38660 5312 38712 5364
rect 13912 5244 13964 5296
rect 16672 5244 16724 5296
rect 7196 5040 7248 5092
rect 10876 5108 10928 5160
rect 12348 5176 12400 5228
rect 14096 5176 14148 5228
rect 15200 5219 15252 5228
rect 15200 5185 15209 5219
rect 15209 5185 15243 5219
rect 15243 5185 15252 5219
rect 15200 5176 15252 5185
rect 16948 5176 17000 5228
rect 17316 5219 17368 5228
rect 17316 5185 17325 5219
rect 17325 5185 17359 5219
rect 17359 5185 17368 5219
rect 17316 5176 17368 5185
rect 17592 5219 17644 5228
rect 17592 5185 17619 5219
rect 17619 5185 17644 5219
rect 17592 5176 17644 5185
rect 11980 5108 12032 5160
rect 13912 5108 13964 5160
rect 8944 5040 8996 5092
rect 7840 4972 7892 5024
rect 10968 4972 11020 5024
rect 12900 5040 12952 5092
rect 12532 4972 12584 5024
rect 13636 5040 13688 5092
rect 13820 5040 13872 5092
rect 14372 5108 14424 5160
rect 14740 5040 14792 5092
rect 21272 5244 21324 5296
rect 24676 5244 24728 5296
rect 18788 5176 18840 5228
rect 19156 5219 19208 5228
rect 19156 5185 19165 5219
rect 19165 5185 19199 5219
rect 19199 5185 19208 5219
rect 19156 5176 19208 5185
rect 22008 5219 22060 5228
rect 22008 5185 22017 5219
rect 22017 5185 22051 5219
rect 22051 5185 22060 5219
rect 22008 5176 22060 5185
rect 22744 5176 22796 5228
rect 18512 5108 18564 5160
rect 19984 5108 20036 5160
rect 20444 5151 20496 5160
rect 20444 5117 20453 5151
rect 20453 5117 20487 5151
rect 20487 5117 20496 5151
rect 20444 5108 20496 5117
rect 18144 5040 18196 5092
rect 19432 5040 19484 5092
rect 23388 5108 23440 5160
rect 23756 5219 23808 5226
rect 23756 5185 23770 5219
rect 23770 5185 23804 5219
rect 23804 5185 23808 5219
rect 23756 5174 23808 5185
rect 24584 5219 24636 5228
rect 23204 5040 23256 5092
rect 24584 5185 24593 5219
rect 24593 5185 24627 5219
rect 24627 5185 24636 5219
rect 24584 5176 24636 5185
rect 24768 5219 24820 5228
rect 24768 5185 24777 5219
rect 24777 5185 24811 5219
rect 24811 5185 24820 5219
rect 24768 5176 24820 5185
rect 25044 5244 25096 5296
rect 29000 5244 29052 5296
rect 30840 5244 30892 5296
rect 24952 5219 25004 5228
rect 24952 5185 24961 5219
rect 24961 5185 24995 5219
rect 24995 5185 25004 5219
rect 24952 5176 25004 5185
rect 27252 5176 27304 5228
rect 27804 5176 27856 5228
rect 30564 5176 30616 5228
rect 31576 5244 31628 5296
rect 33324 5219 33376 5228
rect 33324 5185 33333 5219
rect 33333 5185 33367 5219
rect 33367 5185 33376 5219
rect 33324 5176 33376 5185
rect 26792 5108 26844 5160
rect 33876 5176 33928 5228
rect 34428 5219 34480 5228
rect 34428 5185 34437 5219
rect 34437 5185 34471 5219
rect 34471 5185 34480 5219
rect 34428 5176 34480 5185
rect 35348 5176 35400 5228
rect 35992 5176 36044 5228
rect 37188 5244 37240 5296
rect 37464 5287 37516 5296
rect 37464 5253 37473 5287
rect 37473 5253 37507 5287
rect 37507 5253 37516 5287
rect 37464 5244 37516 5253
rect 38752 5244 38804 5296
rect 36268 5219 36320 5228
rect 36268 5185 36277 5219
rect 36277 5185 36311 5219
rect 36311 5185 36320 5219
rect 36268 5176 36320 5185
rect 36452 5219 36504 5228
rect 36452 5185 36461 5219
rect 36461 5185 36495 5219
rect 36495 5185 36504 5219
rect 36452 5176 36504 5185
rect 37372 5176 37424 5228
rect 38752 5108 38804 5160
rect 58808 5108 58860 5160
rect 14004 4972 14056 5024
rect 17868 4972 17920 5024
rect 19340 4972 19392 5024
rect 19984 5015 20036 5024
rect 19984 4981 19993 5015
rect 19993 4981 20027 5015
rect 20027 4981 20036 5015
rect 19984 4972 20036 4981
rect 20076 4972 20128 5024
rect 22744 5015 22796 5024
rect 22744 4981 22753 5015
rect 22753 4981 22787 5015
rect 22787 4981 22796 5015
rect 22744 4972 22796 4981
rect 59268 5040 59320 5092
rect 25228 5015 25280 5024
rect 25228 4981 25237 5015
rect 25237 4981 25271 5015
rect 25271 4981 25280 5015
rect 25228 4972 25280 4981
rect 26700 4972 26752 5024
rect 27620 4972 27672 5024
rect 32864 5015 32916 5024
rect 32864 4981 32873 5015
rect 32873 4981 32907 5015
rect 32907 4981 32916 5015
rect 32864 4972 32916 4981
rect 33784 4972 33836 5024
rect 35624 4972 35676 5024
rect 58716 4972 58768 5024
rect 67640 5015 67692 5024
rect 67640 4981 67649 5015
rect 67649 4981 67683 5015
rect 67683 4981 67692 5015
rect 67640 4972 67692 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 65654 4870 65706 4922
rect 65718 4870 65770 4922
rect 65782 4870 65834 4922
rect 65846 4870 65898 4922
rect 65910 4870 65962 4922
rect 6920 4768 6972 4820
rect 9772 4768 9824 4820
rect 10600 4811 10652 4820
rect 10600 4777 10609 4811
rect 10609 4777 10643 4811
rect 10643 4777 10652 4811
rect 10600 4768 10652 4777
rect 11980 4811 12032 4820
rect 11980 4777 11989 4811
rect 11989 4777 12023 4811
rect 12023 4777 12032 4811
rect 11980 4768 12032 4777
rect 13728 4768 13780 4820
rect 17960 4768 18012 4820
rect 18236 4768 18288 4820
rect 22100 4768 22152 4820
rect 2780 4700 2832 4752
rect 6644 4700 6696 4752
rect 2320 4632 2372 4684
rect 7472 4675 7524 4684
rect 7472 4641 7481 4675
rect 7481 4641 7515 4675
rect 7515 4641 7524 4675
rect 7472 4632 7524 4641
rect 1400 4607 1452 4616
rect 1400 4573 1409 4607
rect 1409 4573 1443 4607
rect 1443 4573 1452 4607
rect 1400 4564 1452 4573
rect 3884 4564 3936 4616
rect 4712 4607 4764 4616
rect 4712 4573 4746 4607
rect 4746 4573 4764 4607
rect 4252 4496 4304 4548
rect 4712 4564 4764 4573
rect 8208 4607 8260 4616
rect 8208 4573 8217 4607
rect 8217 4573 8251 4607
rect 8251 4573 8260 4607
rect 8208 4564 8260 4573
rect 8944 4607 8996 4616
rect 8944 4573 8953 4607
rect 8953 4573 8987 4607
rect 8987 4573 8996 4607
rect 8944 4564 8996 4573
rect 10048 4700 10100 4752
rect 11704 4743 11756 4752
rect 11704 4709 11728 4743
rect 11728 4709 11756 4743
rect 11704 4700 11756 4709
rect 11796 4743 11848 4752
rect 11796 4709 11805 4743
rect 11805 4709 11839 4743
rect 11839 4709 11848 4743
rect 11796 4700 11848 4709
rect 12072 4700 12124 4752
rect 12532 4700 12584 4752
rect 13452 4700 13504 4752
rect 13820 4700 13872 4752
rect 14096 4743 14148 4752
rect 14096 4709 14105 4743
rect 14105 4709 14139 4743
rect 14139 4709 14148 4743
rect 14096 4700 14148 4709
rect 9496 4607 9548 4616
rect 9496 4573 9505 4607
rect 9505 4573 9539 4607
rect 9539 4573 9548 4607
rect 9496 4564 9548 4573
rect 10048 4564 10100 4616
rect 12440 4564 12492 4616
rect 13636 4632 13688 4684
rect 4620 4496 4672 4548
rect 7840 4496 7892 4548
rect 9036 4496 9088 4548
rect 11152 4496 11204 4548
rect 11980 4496 12032 4548
rect 13912 4564 13964 4616
rect 14464 4564 14516 4616
rect 14740 4632 14792 4684
rect 15936 4675 15988 4684
rect 15936 4641 15945 4675
rect 15945 4641 15979 4675
rect 15979 4641 15988 4675
rect 15936 4632 15988 4641
rect 16028 4675 16080 4684
rect 16028 4641 16037 4675
rect 16037 4641 16071 4675
rect 16071 4641 16080 4675
rect 16028 4632 16080 4641
rect 17960 4632 18012 4684
rect 18144 4700 18196 4752
rect 18696 4743 18748 4752
rect 18696 4709 18705 4743
rect 18705 4709 18739 4743
rect 18739 4709 18748 4743
rect 18696 4700 18748 4709
rect 20260 4700 20312 4752
rect 23756 4768 23808 4820
rect 27160 4811 27212 4820
rect 27160 4777 27169 4811
rect 27169 4777 27203 4811
rect 27203 4777 27212 4811
rect 27160 4768 27212 4777
rect 27344 4768 27396 4820
rect 33324 4768 33376 4820
rect 33876 4811 33928 4820
rect 33876 4777 33885 4811
rect 33885 4777 33919 4811
rect 33919 4777 33928 4811
rect 33876 4768 33928 4777
rect 34428 4768 34480 4820
rect 36268 4768 36320 4820
rect 37464 4768 37516 4820
rect 22744 4700 22796 4752
rect 25596 4700 25648 4752
rect 57244 4700 57296 4752
rect 58256 4700 58308 4752
rect 24308 4632 24360 4684
rect 29000 4675 29052 4684
rect 29000 4641 29009 4675
rect 29009 4641 29043 4675
rect 29043 4641 29052 4675
rect 29000 4632 29052 4641
rect 38752 4675 38804 4684
rect 38752 4641 38761 4675
rect 38761 4641 38795 4675
rect 38795 4641 38804 4675
rect 38752 4632 38804 4641
rect 58900 4632 58952 4684
rect 19156 4564 19208 4616
rect 1952 4428 2004 4480
rect 2412 4471 2464 4480
rect 2412 4437 2421 4471
rect 2421 4437 2455 4471
rect 2455 4437 2464 4471
rect 2412 4428 2464 4437
rect 2688 4428 2740 4480
rect 4712 4428 4764 4480
rect 8392 4471 8444 4480
rect 8392 4437 8401 4471
rect 8401 4437 8435 4471
rect 8435 4437 8444 4471
rect 8392 4428 8444 4437
rect 9312 4428 9364 4480
rect 10140 4428 10192 4480
rect 10324 4428 10376 4480
rect 12532 4428 12584 4480
rect 13636 4496 13688 4548
rect 15568 4428 15620 4480
rect 15844 4471 15896 4480
rect 15844 4437 15853 4471
rect 15853 4437 15887 4471
rect 15887 4437 15896 4471
rect 15844 4428 15896 4437
rect 18052 4496 18104 4548
rect 19984 4564 20036 4616
rect 23020 4564 23072 4616
rect 23480 4564 23532 4616
rect 25228 4564 25280 4616
rect 32404 4564 32456 4616
rect 34796 4564 34848 4616
rect 36084 4564 36136 4616
rect 37740 4564 37792 4616
rect 57152 4564 57204 4616
rect 57612 4564 57664 4616
rect 18236 4428 18288 4480
rect 18880 4428 18932 4480
rect 19432 4428 19484 4480
rect 21272 4496 21324 4548
rect 24952 4496 25004 4548
rect 27712 4496 27764 4548
rect 34704 4496 34756 4548
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 2228 4224 2280 4276
rect 2964 4156 3016 4208
rect 8668 4224 8720 4276
rect 9404 4224 9456 4276
rect 9496 4224 9548 4276
rect 10600 4267 10652 4276
rect 10600 4233 10609 4267
rect 10609 4233 10643 4267
rect 10643 4233 10652 4267
rect 10600 4224 10652 4233
rect 1952 4131 2004 4140
rect 1952 4097 1961 4131
rect 1961 4097 1995 4131
rect 1995 4097 2004 4131
rect 1952 4088 2004 4097
rect 1768 4063 1820 4072
rect 1768 4029 1777 4063
rect 1777 4029 1811 4063
rect 1811 4029 1820 4063
rect 1768 4020 1820 4029
rect 1952 3884 2004 3936
rect 3700 4088 3752 4140
rect 5080 4088 5132 4140
rect 5632 4131 5684 4140
rect 5632 4097 5641 4131
rect 5641 4097 5675 4131
rect 5675 4097 5684 4131
rect 5632 4088 5684 4097
rect 8208 4156 8260 4208
rect 10324 4156 10376 4208
rect 2872 4063 2924 4072
rect 2872 4029 2881 4063
rect 2881 4029 2915 4063
rect 2915 4029 2924 4063
rect 2872 4020 2924 4029
rect 3056 3884 3108 3936
rect 6736 4063 6788 4072
rect 6736 4029 6745 4063
rect 6745 4029 6779 4063
rect 6779 4029 6788 4063
rect 6736 4020 6788 4029
rect 8024 4088 8076 4140
rect 8300 4088 8352 4140
rect 9128 4131 9180 4140
rect 9128 4097 9137 4131
rect 9137 4097 9171 4131
rect 9171 4097 9180 4131
rect 9128 4088 9180 4097
rect 9772 4131 9824 4140
rect 9772 4097 9781 4131
rect 9781 4097 9815 4131
rect 9815 4097 9824 4131
rect 9772 4088 9824 4097
rect 10692 4088 10744 4140
rect 12072 4224 12124 4276
rect 13268 4224 13320 4276
rect 14372 4224 14424 4276
rect 16212 4224 16264 4276
rect 18144 4224 18196 4276
rect 18236 4224 18288 4276
rect 18604 4224 18656 4276
rect 19432 4224 19484 4276
rect 20444 4224 20496 4276
rect 23388 4224 23440 4276
rect 11704 4156 11756 4208
rect 11888 4156 11940 4208
rect 12348 4156 12400 4208
rect 15108 4156 15160 4208
rect 17960 4156 18012 4208
rect 19064 4156 19116 4208
rect 7840 4063 7892 4072
rect 7840 4029 7849 4063
rect 7849 4029 7883 4063
rect 7883 4029 7892 4063
rect 7840 4020 7892 4029
rect 9312 4020 9364 4072
rect 13728 4088 13780 4140
rect 34796 4224 34848 4276
rect 36084 4224 36136 4276
rect 26792 4156 26844 4208
rect 15384 4131 15436 4140
rect 15384 4097 15393 4131
rect 15393 4097 15427 4131
rect 15427 4097 15436 4131
rect 15384 4088 15436 4097
rect 15568 4131 15620 4140
rect 15568 4097 15577 4131
rect 15577 4097 15611 4131
rect 15611 4097 15620 4131
rect 15568 4088 15620 4097
rect 17776 4131 17828 4140
rect 17776 4097 17794 4131
rect 17794 4097 17828 4131
rect 18052 4131 18104 4140
rect 17776 4088 17828 4097
rect 18052 4097 18061 4131
rect 18061 4097 18095 4131
rect 18095 4097 18104 4131
rect 18052 4088 18104 4097
rect 18696 4131 18748 4140
rect 18696 4097 18705 4131
rect 18705 4097 18739 4131
rect 18739 4097 18748 4131
rect 18696 4088 18748 4097
rect 23204 4131 23256 4140
rect 23204 4097 23213 4131
rect 23213 4097 23247 4131
rect 23247 4097 23256 4131
rect 23204 4088 23256 4097
rect 12072 4020 12124 4072
rect 12348 4063 12400 4072
rect 12348 4029 12357 4063
rect 12357 4029 12391 4063
rect 12391 4029 12400 4063
rect 12348 4020 12400 4029
rect 12808 4020 12860 4072
rect 13452 4063 13504 4072
rect 13452 4029 13461 4063
rect 13461 4029 13495 4063
rect 13495 4029 13504 4063
rect 13452 4020 13504 4029
rect 8208 3952 8260 4004
rect 4252 3927 4304 3936
rect 4252 3893 4261 3927
rect 4261 3893 4295 3927
rect 4295 3893 4304 3927
rect 4252 3884 4304 3893
rect 10692 3952 10744 4004
rect 9128 3884 9180 3936
rect 11244 3952 11296 4004
rect 11796 3995 11848 4004
rect 11796 3961 11805 3995
rect 11805 3961 11839 3995
rect 11839 3961 11848 3995
rect 11796 3952 11848 3961
rect 11888 3952 11940 4004
rect 10968 3884 11020 3936
rect 12072 3884 12124 3936
rect 12164 3927 12216 3936
rect 12164 3893 12173 3927
rect 12173 3893 12207 3927
rect 12207 3893 12216 3927
rect 14096 4020 14148 4072
rect 15108 4020 15160 4072
rect 18512 4063 18564 4072
rect 13912 3995 13964 4004
rect 13912 3961 13921 3995
rect 13921 3961 13955 3995
rect 13955 3961 13964 3995
rect 13912 3952 13964 3961
rect 13820 3927 13872 3936
rect 12164 3884 12216 3893
rect 13820 3893 13829 3927
rect 13829 3893 13863 3927
rect 13863 3893 13872 3927
rect 13820 3884 13872 3893
rect 15200 3884 15252 3936
rect 18512 4029 18521 4063
rect 18521 4029 18555 4063
rect 18555 4029 18564 4063
rect 18512 4020 18564 4029
rect 18604 4020 18656 4072
rect 20168 4020 20220 4072
rect 23112 4020 23164 4072
rect 23664 4088 23716 4140
rect 24308 4131 24360 4140
rect 24308 4097 24317 4131
rect 24317 4097 24351 4131
rect 24351 4097 24360 4131
rect 24308 4088 24360 4097
rect 15936 3952 15988 4004
rect 18696 3952 18748 4004
rect 18972 3952 19024 4004
rect 20260 3952 20312 4004
rect 27344 4131 27396 4140
rect 27344 4097 27353 4131
rect 27353 4097 27387 4131
rect 27387 4097 27396 4131
rect 27344 4088 27396 4097
rect 27528 4131 27580 4140
rect 27528 4097 27537 4131
rect 27537 4097 27571 4131
rect 27571 4097 27580 4131
rect 27528 4088 27580 4097
rect 27896 4088 27948 4140
rect 30840 4088 30892 4140
rect 33140 4088 33192 4140
rect 33784 4131 33836 4140
rect 33784 4097 33818 4131
rect 33818 4097 33836 4131
rect 33784 4088 33836 4097
rect 35900 4156 35952 4208
rect 38752 4156 38804 4208
rect 35624 4131 35676 4140
rect 35624 4097 35658 4131
rect 35658 4097 35676 4131
rect 35624 4088 35676 4097
rect 57980 4088 58032 4140
rect 20444 3884 20496 3936
rect 21180 3927 21232 3936
rect 21180 3893 21189 3927
rect 21189 3893 21223 3927
rect 21223 3893 21232 3927
rect 25964 3952 26016 4004
rect 59176 4020 59228 4072
rect 27804 3952 27856 4004
rect 57520 3952 57572 4004
rect 58624 3952 58676 4004
rect 21180 3884 21232 3893
rect 22376 3884 22428 3936
rect 26332 3927 26384 3936
rect 26332 3893 26341 3927
rect 26341 3893 26375 3927
rect 26375 3893 26384 3927
rect 26332 3884 26384 3893
rect 32588 3884 32640 3936
rect 56140 3884 56192 3936
rect 56324 3884 56376 3936
rect 56968 3884 57020 3936
rect 58072 3884 58124 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 65654 3782 65706 3834
rect 65718 3782 65770 3834
rect 65782 3782 65834 3834
rect 65846 3782 65898 3834
rect 65910 3782 65962 3834
rect 3884 3680 3936 3732
rect 2320 3544 2372 3596
rect 3792 3587 3844 3596
rect 3792 3553 3801 3587
rect 3801 3553 3835 3587
rect 3835 3553 3844 3587
rect 3792 3544 3844 3553
rect 3056 3519 3108 3528
rect 3056 3485 3065 3519
rect 3065 3485 3099 3519
rect 3099 3485 3108 3519
rect 3056 3476 3108 3485
rect 3884 3476 3936 3528
rect 7472 3680 7524 3732
rect 7748 3723 7800 3732
rect 7748 3689 7757 3723
rect 7757 3689 7791 3723
rect 7791 3689 7800 3723
rect 7748 3680 7800 3689
rect 9036 3680 9088 3732
rect 9312 3723 9364 3732
rect 9312 3689 9321 3723
rect 9321 3689 9355 3723
rect 9355 3689 9364 3723
rect 9312 3680 9364 3689
rect 9864 3680 9916 3732
rect 10784 3723 10836 3732
rect 10784 3689 10793 3723
rect 10793 3689 10827 3723
rect 10827 3689 10836 3723
rect 10784 3680 10836 3689
rect 10876 3680 10928 3732
rect 11796 3723 11848 3732
rect 11796 3689 11805 3723
rect 11805 3689 11839 3723
rect 11839 3689 11848 3723
rect 11796 3680 11848 3689
rect 11888 3723 11940 3732
rect 11888 3689 11897 3723
rect 11897 3689 11931 3723
rect 11931 3689 11940 3723
rect 11888 3680 11940 3689
rect 12900 3680 12952 3732
rect 14096 3680 14148 3732
rect 14372 3680 14424 3732
rect 15844 3680 15896 3732
rect 21180 3680 21232 3732
rect 23112 3680 23164 3732
rect 27712 3680 27764 3732
rect 32404 3680 32456 3732
rect 57796 3680 57848 3732
rect 58072 3680 58124 3732
rect 7932 3612 7984 3664
rect 8392 3612 8444 3664
rect 8208 3544 8260 3596
rect 6368 3476 6420 3528
rect 6552 3476 6604 3528
rect 7288 3476 7340 3528
rect 7932 3519 7984 3528
rect 7932 3485 7941 3519
rect 7941 3485 7975 3519
rect 7975 3485 7984 3519
rect 7932 3476 7984 3485
rect 9128 3519 9180 3528
rect 1768 3340 1820 3392
rect 2228 3383 2280 3392
rect 2228 3349 2237 3383
rect 2237 3349 2271 3383
rect 2271 3349 2280 3383
rect 2228 3340 2280 3349
rect 7564 3408 7616 3460
rect 5264 3383 5316 3392
rect 5264 3349 5273 3383
rect 5273 3349 5307 3383
rect 5307 3349 5316 3383
rect 5264 3340 5316 3349
rect 5356 3383 5408 3392
rect 5356 3349 5365 3383
rect 5365 3349 5399 3383
rect 5399 3349 5408 3383
rect 5356 3340 5408 3349
rect 6460 3340 6512 3392
rect 7104 3340 7156 3392
rect 7196 3340 7248 3392
rect 9128 3485 9137 3519
rect 9137 3485 9171 3519
rect 9171 3485 9180 3519
rect 9128 3476 9180 3485
rect 11244 3544 11296 3596
rect 10416 3408 10468 3460
rect 10600 3451 10652 3460
rect 10600 3417 10609 3451
rect 10609 3417 10643 3451
rect 10643 3417 10652 3451
rect 10600 3408 10652 3417
rect 9680 3340 9732 3392
rect 10140 3383 10192 3392
rect 10140 3349 10149 3383
rect 10149 3349 10183 3383
rect 10183 3349 10192 3383
rect 10140 3340 10192 3349
rect 14740 3612 14792 3664
rect 15200 3612 15252 3664
rect 17960 3612 18012 3664
rect 18972 3612 19024 3664
rect 19340 3655 19392 3664
rect 19340 3621 19349 3655
rect 19349 3621 19383 3655
rect 19383 3621 19392 3655
rect 19340 3612 19392 3621
rect 22652 3612 22704 3664
rect 41144 3612 41196 3664
rect 56508 3612 56560 3664
rect 58348 3612 58400 3664
rect 12348 3544 12400 3596
rect 18880 3544 18932 3596
rect 20076 3544 20128 3596
rect 24584 3544 24636 3596
rect 11796 3408 11848 3460
rect 12900 3476 12952 3528
rect 14280 3408 14332 3460
rect 14464 3519 14516 3528
rect 14464 3485 14473 3519
rect 14473 3485 14507 3519
rect 14507 3485 14516 3519
rect 14464 3476 14516 3485
rect 14832 3408 14884 3460
rect 12440 3340 12492 3392
rect 13360 3340 13412 3392
rect 14372 3340 14424 3392
rect 15660 3476 15712 3528
rect 17408 3476 17460 3528
rect 17868 3519 17920 3528
rect 17868 3485 17877 3519
rect 17877 3485 17911 3519
rect 17911 3485 17920 3519
rect 17868 3476 17920 3485
rect 19984 3476 20036 3528
rect 20996 3476 21048 3528
rect 23204 3476 23256 3528
rect 24860 3476 24912 3528
rect 25688 3476 25740 3528
rect 26240 3476 26292 3528
rect 27344 3544 27396 3596
rect 33140 3587 33192 3596
rect 33140 3553 33149 3587
rect 33149 3553 33183 3587
rect 33183 3553 33192 3587
rect 33140 3544 33192 3553
rect 55772 3544 55824 3596
rect 56784 3544 56836 3596
rect 58992 3544 59044 3596
rect 26700 3519 26752 3528
rect 26700 3485 26709 3519
rect 26709 3485 26743 3519
rect 26743 3485 26752 3519
rect 26700 3476 26752 3485
rect 26792 3519 26844 3528
rect 26792 3485 26801 3519
rect 26801 3485 26835 3519
rect 26835 3485 26844 3519
rect 26792 3476 26844 3485
rect 26976 3476 27028 3528
rect 27896 3476 27948 3528
rect 28724 3476 28776 3528
rect 29552 3476 29604 3528
rect 30656 3519 30708 3528
rect 30656 3485 30665 3519
rect 30665 3485 30699 3519
rect 30699 3485 30708 3519
rect 30656 3476 30708 3485
rect 31208 3476 31260 3528
rect 32864 3519 32916 3528
rect 32864 3485 32882 3519
rect 32882 3485 32916 3519
rect 32864 3476 32916 3485
rect 39212 3476 39264 3528
rect 40040 3476 40092 3528
rect 40868 3476 40920 3528
rect 42524 3476 42576 3528
rect 43076 3476 43128 3528
rect 45008 3476 45060 3528
rect 45284 3476 45336 3528
rect 46112 3476 46164 3528
rect 46940 3476 46992 3528
rect 47768 3476 47820 3528
rect 48872 3476 48924 3528
rect 50160 3476 50212 3528
rect 50804 3476 50856 3528
rect 51356 3476 51408 3528
rect 52736 3476 52788 3528
rect 53012 3476 53064 3528
rect 54668 3476 54720 3528
rect 55496 3476 55548 3528
rect 56232 3476 56284 3528
rect 57336 3476 57388 3528
rect 60464 3519 60516 3528
rect 60464 3485 60473 3519
rect 60473 3485 60507 3519
rect 60507 3485 60516 3519
rect 60464 3476 60516 3485
rect 68100 3519 68152 3528
rect 68100 3485 68109 3519
rect 68109 3485 68143 3519
rect 68143 3485 68152 3519
rect 68100 3476 68152 3485
rect 15108 3408 15160 3460
rect 18420 3408 18472 3460
rect 16488 3383 16540 3392
rect 16488 3349 16497 3383
rect 16497 3349 16531 3383
rect 16531 3349 16540 3383
rect 16488 3340 16540 3349
rect 19432 3408 19484 3460
rect 20076 3451 20128 3460
rect 20076 3417 20085 3451
rect 20085 3417 20119 3451
rect 20119 3417 20128 3451
rect 20076 3408 20128 3417
rect 23020 3408 23072 3460
rect 25964 3408 26016 3460
rect 20168 3340 20220 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 1400 3136 1452 3188
rect 3976 3179 4028 3188
rect 3976 3145 3985 3179
rect 3985 3145 4019 3179
rect 4019 3145 4028 3179
rect 3976 3136 4028 3145
rect 1768 3043 1820 3052
rect 1768 3009 1777 3043
rect 1777 3009 1811 3043
rect 1811 3009 1820 3043
rect 1768 3000 1820 3009
rect 1952 3043 2004 3052
rect 1952 3009 1961 3043
rect 1961 3009 1995 3043
rect 1995 3009 2004 3043
rect 1952 3000 2004 3009
rect 2964 3068 3016 3120
rect 2872 3043 2924 3052
rect 2872 3009 2906 3043
rect 2906 3009 2924 3043
rect 4620 3136 4672 3188
rect 5356 3136 5408 3188
rect 7012 3136 7064 3188
rect 8024 3136 8076 3188
rect 8116 3136 8168 3188
rect 8944 3136 8996 3188
rect 10140 3136 10192 3188
rect 11612 3136 11664 3188
rect 11888 3136 11940 3188
rect 11980 3136 12032 3188
rect 12256 3136 12308 3188
rect 12992 3136 13044 3188
rect 13360 3136 13412 3188
rect 16488 3136 16540 3188
rect 19340 3136 19392 3188
rect 19432 3136 19484 3188
rect 20260 3136 20312 3188
rect 22008 3136 22060 3188
rect 26424 3136 26476 3188
rect 26976 3179 27028 3188
rect 26976 3145 26985 3179
rect 26985 3145 27019 3179
rect 27019 3145 27028 3179
rect 26976 3136 27028 3145
rect 55956 3136 56008 3188
rect 58072 3136 58124 3188
rect 4712 3111 4764 3120
rect 4712 3077 4746 3111
rect 4746 3077 4764 3111
rect 4712 3068 4764 3077
rect 2872 3000 2924 3009
rect 6460 3000 6512 3052
rect 7104 3000 7156 3052
rect 6368 2796 6420 2848
rect 9220 3000 9272 3052
rect 9956 3068 10008 3120
rect 10048 3068 10100 3120
rect 12900 3068 12952 3120
rect 13084 3111 13136 3120
rect 13084 3077 13093 3111
rect 13093 3077 13127 3111
rect 13127 3077 13136 3111
rect 13084 3068 13136 3077
rect 13820 3068 13872 3120
rect 15108 3068 15160 3120
rect 17868 3068 17920 3120
rect 20628 3068 20680 3120
rect 57704 3068 57756 3120
rect 60464 3068 60516 3120
rect 11612 3000 11664 3052
rect 11796 3000 11848 3052
rect 11244 2932 11296 2984
rect 12164 3000 12216 3052
rect 12348 3043 12400 3052
rect 12348 3009 12357 3043
rect 12357 3009 12391 3043
rect 12391 3009 12400 3043
rect 12348 3000 12400 3009
rect 12440 2932 12492 2984
rect 13544 3043 13596 3052
rect 13544 3009 13553 3043
rect 13553 3009 13587 3043
rect 13587 3009 13596 3043
rect 13544 3000 13596 3009
rect 13912 3000 13964 3052
rect 14556 3000 14608 3052
rect 16856 3000 16908 3052
rect 17592 3043 17644 3052
rect 17592 3009 17601 3043
rect 17601 3009 17635 3043
rect 17635 3009 17644 3043
rect 17592 3000 17644 3009
rect 20076 3000 20128 3052
rect 58164 3000 58216 3052
rect 14280 2932 14332 2984
rect 18696 2932 18748 2984
rect 20720 2932 20772 2984
rect 21824 2932 21876 2984
rect 25136 2932 25188 2984
rect 29000 2932 29052 2984
rect 30932 2932 30984 2984
rect 37280 2932 37332 2984
rect 44732 2932 44784 2984
rect 48596 2932 48648 2984
rect 52460 2932 52512 2984
rect 53564 2932 53616 2984
rect 55220 2932 55272 2984
rect 56692 2932 56744 2984
rect 11796 2864 11848 2916
rect 11888 2864 11940 2916
rect 11704 2796 11756 2848
rect 13268 2864 13320 2916
rect 13636 2864 13688 2916
rect 20260 2864 20312 2916
rect 14188 2796 14240 2848
rect 17776 2796 17828 2848
rect 20168 2796 20220 2848
rect 22008 2864 22060 2916
rect 23480 2864 23532 2916
rect 21272 2796 21324 2848
rect 23756 2796 23808 2848
rect 24308 2796 24360 2848
rect 25964 2864 26016 2916
rect 27068 2864 27120 2916
rect 38384 2864 38436 2916
rect 39764 2864 39816 2916
rect 42248 2864 42300 2916
rect 43628 2864 43680 2916
rect 47492 2864 47544 2916
rect 49424 2864 49476 2916
rect 50620 2864 50672 2916
rect 53288 2864 53340 2916
rect 54392 2864 54444 2916
rect 55680 2864 55732 2916
rect 57060 2864 57112 2916
rect 58440 2932 58492 2984
rect 26792 2796 26844 2848
rect 28172 2796 28224 2848
rect 29276 2796 29328 2848
rect 30104 2796 30156 2848
rect 31484 2796 31536 2848
rect 32036 2796 32088 2848
rect 33140 2796 33192 2848
rect 33692 2796 33744 2848
rect 34244 2796 34296 2848
rect 34520 2796 34572 2848
rect 35348 2796 35400 2848
rect 36176 2796 36228 2848
rect 36728 2796 36780 2848
rect 37832 2796 37884 2848
rect 38936 2796 38988 2848
rect 40316 2796 40368 2848
rect 41696 2796 41748 2848
rect 42800 2796 42852 2848
rect 44180 2796 44232 2848
rect 45560 2796 45612 2848
rect 46664 2796 46716 2848
rect 48044 2796 48096 2848
rect 49976 2796 50028 2848
rect 51908 2796 51960 2848
rect 53840 2796 53892 2848
rect 55404 2796 55456 2848
rect 56048 2796 56100 2848
rect 59360 2864 59412 2916
rect 59452 2796 59504 2848
rect 60464 2839 60516 2848
rect 60464 2805 60473 2839
rect 60473 2805 60507 2839
rect 60507 2805 60516 2839
rect 60464 2796 60516 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 65654 2694 65706 2746
rect 65718 2694 65770 2746
rect 65782 2694 65834 2746
rect 65846 2694 65898 2746
rect 65910 2694 65962 2746
rect 8300 2592 8352 2644
rect 10416 2592 10468 2644
rect 10508 2592 10560 2644
rect 12808 2592 12860 2644
rect 14832 2635 14884 2644
rect 14832 2601 14841 2635
rect 14841 2601 14875 2635
rect 14875 2601 14884 2635
rect 14832 2592 14884 2601
rect 17960 2592 18012 2644
rect 10784 2524 10836 2576
rect 11060 2524 11112 2576
rect 12440 2524 12492 2576
rect 14464 2524 14516 2576
rect 17592 2524 17644 2576
rect 55220 2592 55272 2644
rect 57428 2592 57480 2644
rect 1768 2431 1820 2440
rect 1768 2397 1777 2431
rect 1777 2397 1811 2431
rect 1811 2397 1820 2431
rect 1768 2388 1820 2397
rect 2504 2388 2556 2440
rect 2964 2388 3016 2440
rect 5172 2456 5224 2508
rect 4896 2431 4948 2440
rect 4896 2397 4905 2431
rect 4905 2397 4939 2431
rect 4939 2397 4948 2431
rect 4896 2388 4948 2397
rect 6368 2388 6420 2440
rect 8484 2456 8536 2508
rect 10048 2456 10100 2508
rect 7656 2431 7708 2440
rect 7656 2397 7665 2431
rect 7665 2397 7699 2431
rect 7699 2397 7708 2431
rect 7656 2388 7708 2397
rect 4344 2320 4396 2372
rect 3240 2295 3292 2304
rect 3240 2261 3249 2295
rect 3249 2261 3283 2295
rect 3283 2261 3292 2295
rect 3240 2252 3292 2261
rect 7196 2320 7248 2372
rect 8760 2388 8812 2440
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 5080 2295 5132 2304
rect 5080 2261 5089 2295
rect 5089 2261 5123 2295
rect 5123 2261 5132 2295
rect 5080 2252 5132 2261
rect 6736 2295 6788 2304
rect 6736 2261 6745 2295
rect 6745 2261 6779 2295
rect 6779 2261 6788 2295
rect 6736 2252 6788 2261
rect 8208 2295 8260 2304
rect 8208 2261 8217 2295
rect 8217 2261 8251 2295
rect 8251 2261 8260 2295
rect 8484 2320 8536 2372
rect 10508 2388 10560 2440
rect 11152 2388 11204 2440
rect 11704 2456 11756 2508
rect 12164 2456 12216 2508
rect 13544 2456 13596 2508
rect 21548 2524 21600 2576
rect 24032 2524 24084 2576
rect 27344 2524 27396 2576
rect 32864 2524 32916 2576
rect 40592 2524 40644 2576
rect 44456 2524 44508 2576
rect 48320 2524 48372 2576
rect 52184 2524 52236 2576
rect 55864 2524 55916 2576
rect 58072 2524 58124 2576
rect 13176 2388 13228 2440
rect 14924 2388 14976 2440
rect 9956 2363 10008 2372
rect 9956 2329 9965 2363
rect 9965 2329 9999 2363
rect 9999 2329 10008 2363
rect 9956 2320 10008 2329
rect 11888 2320 11940 2372
rect 12716 2320 12768 2372
rect 13544 2320 13596 2372
rect 13728 2320 13780 2372
rect 8208 2252 8260 2261
rect 11060 2252 11112 2304
rect 12992 2295 13044 2304
rect 12992 2261 13001 2295
rect 13001 2261 13035 2295
rect 13035 2261 13044 2295
rect 12992 2252 13044 2261
rect 14096 2252 14148 2304
rect 18144 2431 18196 2440
rect 16764 2295 16816 2304
rect 16764 2261 16773 2295
rect 16773 2261 16807 2295
rect 16807 2261 16816 2295
rect 18144 2397 18153 2431
rect 18153 2397 18187 2431
rect 18187 2397 18196 2431
rect 18144 2388 18196 2397
rect 17592 2363 17644 2372
rect 17592 2329 17601 2363
rect 17601 2329 17635 2363
rect 17635 2329 17644 2363
rect 22100 2456 22152 2508
rect 24584 2456 24636 2508
rect 26516 2456 26568 2508
rect 28448 2456 28500 2508
rect 30380 2456 30432 2508
rect 37004 2456 37056 2508
rect 38108 2456 38160 2508
rect 41420 2456 41472 2508
rect 43352 2456 43404 2508
rect 46388 2456 46440 2508
rect 49148 2456 49200 2508
rect 51080 2456 51132 2508
rect 54944 2456 54996 2508
rect 63684 2499 63736 2508
rect 17592 2320 17644 2329
rect 20536 2320 20588 2372
rect 22928 2388 22980 2440
rect 25412 2388 25464 2440
rect 27620 2388 27672 2440
rect 29828 2388 29880 2440
rect 32312 2388 32364 2440
rect 33416 2388 33468 2440
rect 33968 2388 34020 2440
rect 34796 2388 34848 2440
rect 35072 2388 35124 2440
rect 35624 2388 35676 2440
rect 35900 2388 35952 2440
rect 36452 2388 36504 2440
rect 37556 2388 37608 2440
rect 38660 2388 38712 2440
rect 31760 2320 31812 2372
rect 39488 2320 39540 2372
rect 41972 2388 42024 2440
rect 43904 2320 43956 2372
rect 45836 2388 45888 2440
rect 47216 2320 47268 2372
rect 49700 2388 49752 2440
rect 51632 2388 51684 2440
rect 54116 2320 54168 2372
rect 56416 2388 56468 2440
rect 16764 2252 16816 2261
rect 18788 2252 18840 2304
rect 19248 2252 19300 2304
rect 20628 2252 20680 2304
rect 56876 2252 56928 2304
rect 63684 2465 63693 2499
rect 63693 2465 63727 2499
rect 63727 2465 63736 2499
rect 63684 2456 63736 2465
rect 61752 2431 61804 2440
rect 61752 2397 61761 2431
rect 61761 2397 61795 2431
rect 61795 2397 61804 2431
rect 61752 2388 61804 2397
rect 63040 2431 63092 2440
rect 63040 2397 63049 2431
rect 63049 2397 63083 2431
rect 63083 2397 63092 2431
rect 63040 2388 63092 2397
rect 66996 2431 67048 2440
rect 66996 2397 67005 2431
rect 67005 2397 67039 2431
rect 67039 2397 67048 2431
rect 66996 2388 67048 2397
rect 67548 2388 67600 2440
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 6736 2048 6788 2100
rect 11704 2048 11756 2100
rect 13176 2048 13228 2100
rect 20352 2048 20404 2100
rect 58072 2048 58124 2100
rect 61752 2048 61804 2100
rect 5080 1980 5132 2032
rect 12164 1980 12216 2032
rect 12348 1980 12400 2032
rect 13728 1980 13780 2032
rect 16764 1980 16816 2032
rect 22744 1980 22796 2032
rect 59084 1980 59136 2032
rect 63684 1980 63736 2032
rect 8852 1912 8904 1964
rect 9956 1912 10008 1964
rect 11244 1912 11296 1964
rect 58532 1912 58584 1964
rect 63040 1912 63092 1964
rect 9128 1844 9180 1896
rect 16672 1844 16724 1896
rect 4344 1776 4396 1828
rect 9864 1776 9916 1828
rect 3240 1708 3292 1760
rect 10600 1708 10652 1760
rect 19800 1708 19852 1760
rect 20628 1708 20680 1760
rect 2964 1640 3016 1692
rect 11060 1640 11112 1692
rect 12624 1368 12676 1420
rect 13176 1368 13228 1420
rect 1768 1300 1820 1352
rect 10324 1300 10376 1352
rect 10692 1300 10744 1352
rect 13084 1300 13136 1352
rect 13544 1368 13596 1420
rect 17592 1368 17644 1420
rect 19524 1300 19576 1352
rect 20168 1300 20220 1352
rect 5172 1232 5224 1284
rect 11888 1232 11940 1284
rect 13544 1232 13596 1284
rect 56784 1164 56836 1216
rect 57060 1164 57112 1216
rect 57060 1028 57112 1080
rect 59452 1028 59504 1080
rect 4896 960 4948 1012
rect 9680 892 9732 944
rect 10876 892 10928 944
rect 12900 892 12952 944
rect 2504 144 2556 196
rect 9680 144 9732 196
<< metal2 >>
rect 5170 59200 5226 60000
rect 15106 59200 15162 60000
rect 25042 59200 25098 60000
rect 34978 59200 35034 60000
rect 44914 59200 44970 60000
rect 54850 59200 54906 60000
rect 64786 59200 64842 60000
rect 67546 59256 67602 59265
rect 5184 57458 5212 59200
rect 15120 57882 15148 59200
rect 15120 57854 15240 57882
rect 15212 57458 15240 57854
rect 19574 57692 19882 57701
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57627 19882 57636
rect 25056 57458 25084 59200
rect 34992 57458 35020 59200
rect 44928 57458 44956 59200
rect 50294 57692 50602 57701
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57627 50602 57636
rect 54864 57458 54892 59200
rect 64800 57458 64828 59200
rect 67546 59191 67602 59200
rect 66994 57896 67050 57905
rect 66994 57831 67050 57840
rect 67008 57458 67036 57831
rect 67560 57458 67588 59191
rect 5172 57452 5224 57458
rect 5172 57394 5224 57400
rect 15200 57452 15252 57458
rect 15200 57394 15252 57400
rect 25044 57452 25096 57458
rect 25044 57394 25096 57400
rect 34980 57452 35032 57458
rect 34980 57394 35032 57400
rect 44916 57452 44968 57458
rect 44916 57394 44968 57400
rect 54852 57452 54904 57458
rect 54852 57394 54904 57400
rect 64788 57452 64840 57458
rect 64788 57394 64840 57400
rect 66996 57452 67048 57458
rect 66996 57394 67048 57400
rect 67548 57452 67600 57458
rect 67548 57394 67600 57400
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 65654 57148 65962 57157
rect 65654 57146 65660 57148
rect 65716 57146 65740 57148
rect 65796 57146 65820 57148
rect 65876 57146 65900 57148
rect 65956 57146 65962 57148
rect 65716 57094 65718 57146
rect 65898 57094 65900 57146
rect 65654 57092 65660 57094
rect 65716 57092 65740 57094
rect 65796 57092 65820 57094
rect 65876 57092 65900 57094
rect 65956 57092 65962 57094
rect 65654 57083 65962 57092
rect 68100 56840 68152 56846
rect 68100 56782 68152 56788
rect 19574 56604 19882 56613
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56539 19882 56548
rect 50294 56604 50602 56613
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56539 50602 56548
rect 68112 56545 68140 56782
rect 68098 56536 68154 56545
rect 68098 56471 68154 56480
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 65654 56060 65962 56069
rect 65654 56058 65660 56060
rect 65716 56058 65740 56060
rect 65796 56058 65820 56060
rect 65876 56058 65900 56060
rect 65956 56058 65962 56060
rect 65716 56006 65718 56058
rect 65898 56006 65900 56058
rect 65654 56004 65660 56006
rect 65716 56004 65740 56006
rect 65796 56004 65820 56006
rect 65876 56004 65900 56006
rect 65956 56004 65962 56006
rect 65654 55995 65962 56004
rect 19574 55516 19882 55525
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55451 19882 55460
rect 50294 55516 50602 55525
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55451 50602 55460
rect 67638 55176 67694 55185
rect 67638 55111 67640 55120
rect 67692 55111 67694 55120
rect 67640 55082 67692 55088
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 65654 54972 65962 54981
rect 65654 54970 65660 54972
rect 65716 54970 65740 54972
rect 65796 54970 65820 54972
rect 65876 54970 65900 54972
rect 65956 54970 65962 54972
rect 65716 54918 65718 54970
rect 65898 54918 65900 54970
rect 65654 54916 65660 54918
rect 65716 54916 65740 54918
rect 65796 54916 65820 54918
rect 65876 54916 65900 54918
rect 65956 54916 65962 54918
rect 65654 54907 65962 54916
rect 19574 54428 19882 54437
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54363 19882 54372
rect 50294 54428 50602 54437
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54363 50602 54372
rect 67548 53984 67600 53990
rect 67548 53926 67600 53932
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 65654 53884 65962 53893
rect 65654 53882 65660 53884
rect 65716 53882 65740 53884
rect 65796 53882 65820 53884
rect 65876 53882 65900 53884
rect 65956 53882 65962 53884
rect 65716 53830 65718 53882
rect 65898 53830 65900 53882
rect 65654 53828 65660 53830
rect 65716 53828 65740 53830
rect 65796 53828 65820 53830
rect 65876 53828 65900 53830
rect 65956 53828 65962 53830
rect 65654 53819 65962 53828
rect 67560 53825 67588 53926
rect 67546 53816 67602 53825
rect 67546 53751 67602 53760
rect 19574 53340 19882 53349
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53275 19882 53284
rect 50294 53340 50602 53349
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53275 50602 53284
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 65654 52796 65962 52805
rect 65654 52794 65660 52796
rect 65716 52794 65740 52796
rect 65796 52794 65820 52796
rect 65876 52794 65900 52796
rect 65956 52794 65962 52796
rect 65716 52742 65718 52794
rect 65898 52742 65900 52794
rect 65654 52740 65660 52742
rect 65716 52740 65740 52742
rect 65796 52740 65820 52742
rect 65876 52740 65900 52742
rect 65956 52740 65962 52742
rect 65654 52731 65962 52740
rect 68100 52488 68152 52494
rect 68098 52456 68100 52465
rect 68152 52456 68154 52465
rect 68098 52391 68154 52400
rect 19574 52252 19882 52261
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52187 19882 52196
rect 50294 52252 50602 52261
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52187 50602 52196
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 65654 51708 65962 51717
rect 65654 51706 65660 51708
rect 65716 51706 65740 51708
rect 65796 51706 65820 51708
rect 65876 51706 65900 51708
rect 65956 51706 65962 51708
rect 65716 51654 65718 51706
rect 65898 51654 65900 51706
rect 65654 51652 65660 51654
rect 65716 51652 65740 51654
rect 65796 51652 65820 51654
rect 65876 51652 65900 51654
rect 65956 51652 65962 51654
rect 65654 51643 65962 51652
rect 68100 51400 68152 51406
rect 68100 51342 68152 51348
rect 19574 51164 19882 51173
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51099 19882 51108
rect 50294 51164 50602 51173
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51099 50602 51108
rect 68112 51105 68140 51342
rect 68098 51096 68154 51105
rect 68098 51031 68154 51040
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 65654 50620 65962 50629
rect 65654 50618 65660 50620
rect 65716 50618 65740 50620
rect 65796 50618 65820 50620
rect 65876 50618 65900 50620
rect 65956 50618 65962 50620
rect 65716 50566 65718 50618
rect 65898 50566 65900 50618
rect 65654 50564 65660 50566
rect 65716 50564 65740 50566
rect 65796 50564 65820 50566
rect 65876 50564 65900 50566
rect 65956 50564 65962 50566
rect 65654 50555 65962 50564
rect 19574 50076 19882 50085
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50011 19882 50020
rect 50294 50076 50602 50085
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50011 50602 50020
rect 67640 49768 67692 49774
rect 67638 49736 67640 49745
rect 67692 49736 67694 49745
rect 67638 49671 67694 49680
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 65654 49532 65962 49541
rect 65654 49530 65660 49532
rect 65716 49530 65740 49532
rect 65796 49530 65820 49532
rect 65876 49530 65900 49532
rect 65956 49530 65962 49532
rect 65716 49478 65718 49530
rect 65898 49478 65900 49530
rect 65654 49476 65660 49478
rect 65716 49476 65740 49478
rect 65796 49476 65820 49478
rect 65876 49476 65900 49478
rect 65956 49476 65962 49478
rect 65654 49467 65962 49476
rect 19574 48988 19882 48997
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48923 19882 48932
rect 50294 48988 50602 48997
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48923 50602 48932
rect 67640 48544 67692 48550
rect 67640 48486 67692 48492
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 65654 48444 65962 48453
rect 65654 48442 65660 48444
rect 65716 48442 65740 48444
rect 65796 48442 65820 48444
rect 65876 48442 65900 48444
rect 65956 48442 65962 48444
rect 65716 48390 65718 48442
rect 65898 48390 65900 48442
rect 65654 48388 65660 48390
rect 65716 48388 65740 48390
rect 65796 48388 65820 48390
rect 65876 48388 65900 48390
rect 65956 48388 65962 48390
rect 65654 48379 65962 48388
rect 67652 48385 67680 48486
rect 67638 48376 67694 48385
rect 67638 48311 67694 48320
rect 19574 47900 19882 47909
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47835 19882 47844
rect 50294 47900 50602 47909
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47835 50602 47844
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 65654 47356 65962 47365
rect 65654 47354 65660 47356
rect 65716 47354 65740 47356
rect 65796 47354 65820 47356
rect 65876 47354 65900 47356
rect 65956 47354 65962 47356
rect 65716 47302 65718 47354
rect 65898 47302 65900 47354
rect 65654 47300 65660 47302
rect 65716 47300 65740 47302
rect 65796 47300 65820 47302
rect 65876 47300 65900 47302
rect 65956 47300 65962 47302
rect 65654 47291 65962 47300
rect 68100 47048 68152 47054
rect 68098 47016 68100 47025
rect 68152 47016 68154 47025
rect 68098 46951 68154 46960
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 50294 46812 50602 46821
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46747 50602 46756
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 65654 46268 65962 46277
rect 65654 46266 65660 46268
rect 65716 46266 65740 46268
rect 65796 46266 65820 46268
rect 65876 46266 65900 46268
rect 65956 46266 65962 46268
rect 65716 46214 65718 46266
rect 65898 46214 65900 46266
rect 65654 46212 65660 46214
rect 65716 46212 65740 46214
rect 65796 46212 65820 46214
rect 65876 46212 65900 46214
rect 65956 46212 65962 46214
rect 65654 46203 65962 46212
rect 68100 45960 68152 45966
rect 68100 45902 68152 45908
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 50294 45724 50602 45733
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45659 50602 45668
rect 68112 45665 68140 45902
rect 68098 45656 68154 45665
rect 68098 45591 68154 45600
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 65654 45180 65962 45189
rect 65654 45178 65660 45180
rect 65716 45178 65740 45180
rect 65796 45178 65820 45180
rect 65876 45178 65900 45180
rect 65956 45178 65962 45180
rect 65716 45126 65718 45178
rect 65898 45126 65900 45178
rect 65654 45124 65660 45126
rect 65716 45124 65740 45126
rect 65796 45124 65820 45126
rect 65876 45124 65900 45126
rect 65956 45124 65962 45126
rect 65654 45115 65962 45124
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 50294 44636 50602 44645
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44571 50602 44580
rect 67638 44296 67694 44305
rect 67638 44231 67640 44240
rect 67692 44231 67694 44240
rect 67640 44202 67692 44208
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 65654 44092 65962 44101
rect 65654 44090 65660 44092
rect 65716 44090 65740 44092
rect 65796 44090 65820 44092
rect 65876 44090 65900 44092
rect 65956 44090 65962 44092
rect 65716 44038 65718 44090
rect 65898 44038 65900 44090
rect 65654 44036 65660 44038
rect 65716 44036 65740 44038
rect 65796 44036 65820 44038
rect 65876 44036 65900 44038
rect 65956 44036 65962 44038
rect 65654 44027 65962 44036
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 50294 43548 50602 43557
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43483 50602 43492
rect 67640 43104 67692 43110
rect 67640 43046 67692 43052
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 65654 43004 65962 43013
rect 65654 43002 65660 43004
rect 65716 43002 65740 43004
rect 65796 43002 65820 43004
rect 65876 43002 65900 43004
rect 65956 43002 65962 43004
rect 65716 42950 65718 43002
rect 65898 42950 65900 43002
rect 65654 42948 65660 42950
rect 65716 42948 65740 42950
rect 65796 42948 65820 42950
rect 65876 42948 65900 42950
rect 65956 42948 65962 42950
rect 65654 42939 65962 42948
rect 67652 42945 67680 43046
rect 67638 42936 67694 42945
rect 67638 42871 67694 42880
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 50294 42460 50602 42469
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42395 50602 42404
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 65654 41916 65962 41925
rect 65654 41914 65660 41916
rect 65716 41914 65740 41916
rect 65796 41914 65820 41916
rect 65876 41914 65900 41916
rect 65956 41914 65962 41916
rect 65716 41862 65718 41914
rect 65898 41862 65900 41914
rect 65654 41860 65660 41862
rect 65716 41860 65740 41862
rect 65796 41860 65820 41862
rect 65876 41860 65900 41862
rect 65956 41860 65962 41862
rect 65654 41851 65962 41860
rect 68100 41608 68152 41614
rect 68098 41576 68100 41585
rect 68152 41576 68154 41585
rect 68098 41511 68154 41520
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 50294 41372 50602 41381
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41307 50602 41316
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 65654 40828 65962 40837
rect 65654 40826 65660 40828
rect 65716 40826 65740 40828
rect 65796 40826 65820 40828
rect 65876 40826 65900 40828
rect 65956 40826 65962 40828
rect 65716 40774 65718 40826
rect 65898 40774 65900 40826
rect 65654 40772 65660 40774
rect 65716 40772 65740 40774
rect 65796 40772 65820 40774
rect 65876 40772 65900 40774
rect 65956 40772 65962 40774
rect 65654 40763 65962 40772
rect 68100 40520 68152 40526
rect 68100 40462 68152 40468
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 50294 40284 50602 40293
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40219 50602 40228
rect 68112 40225 68140 40462
rect 68098 40216 68154 40225
rect 68098 40151 68154 40160
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 65654 39740 65962 39749
rect 65654 39738 65660 39740
rect 65716 39738 65740 39740
rect 65796 39738 65820 39740
rect 65876 39738 65900 39740
rect 65956 39738 65962 39740
rect 65716 39686 65718 39738
rect 65898 39686 65900 39738
rect 65654 39684 65660 39686
rect 65716 39684 65740 39686
rect 65796 39684 65820 39686
rect 65876 39684 65900 39686
rect 65956 39684 65962 39686
rect 65654 39675 65962 39684
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 67638 38856 67694 38865
rect 67638 38791 67640 38800
rect 67692 38791 67694 38800
rect 67640 38762 67692 38768
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 65654 38652 65962 38661
rect 65654 38650 65660 38652
rect 65716 38650 65740 38652
rect 65796 38650 65820 38652
rect 65876 38650 65900 38652
rect 65956 38650 65962 38652
rect 65716 38598 65718 38650
rect 65898 38598 65900 38650
rect 65654 38596 65660 38598
rect 65716 38596 65740 38598
rect 65796 38596 65820 38598
rect 65876 38596 65900 38598
rect 65956 38596 65962 38598
rect 65654 38587 65962 38596
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 67640 37664 67692 37670
rect 67640 37606 67692 37612
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 65654 37564 65962 37573
rect 65654 37562 65660 37564
rect 65716 37562 65740 37564
rect 65796 37562 65820 37564
rect 65876 37562 65900 37564
rect 65956 37562 65962 37564
rect 65716 37510 65718 37562
rect 65898 37510 65900 37562
rect 65654 37508 65660 37510
rect 65716 37508 65740 37510
rect 65796 37508 65820 37510
rect 65876 37508 65900 37510
rect 65956 37508 65962 37510
rect 65654 37499 65962 37508
rect 67652 37505 67680 37606
rect 67638 37496 67694 37505
rect 67638 37431 67694 37440
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 65654 36476 65962 36485
rect 65654 36474 65660 36476
rect 65716 36474 65740 36476
rect 65796 36474 65820 36476
rect 65876 36474 65900 36476
rect 65956 36474 65962 36476
rect 65716 36422 65718 36474
rect 65898 36422 65900 36474
rect 65654 36420 65660 36422
rect 65716 36420 65740 36422
rect 65796 36420 65820 36422
rect 65876 36420 65900 36422
rect 65956 36420 65962 36422
rect 65654 36411 65962 36420
rect 68100 36168 68152 36174
rect 68098 36136 68100 36145
rect 68152 36136 68154 36145
rect 68098 36071 68154 36080
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 65654 35388 65962 35397
rect 65654 35386 65660 35388
rect 65716 35386 65740 35388
rect 65796 35386 65820 35388
rect 65876 35386 65900 35388
rect 65956 35386 65962 35388
rect 65716 35334 65718 35386
rect 65898 35334 65900 35386
rect 65654 35332 65660 35334
rect 65716 35332 65740 35334
rect 65796 35332 65820 35334
rect 65876 35332 65900 35334
rect 65956 35332 65962 35334
rect 65654 35323 65962 35332
rect 68100 35080 68152 35086
rect 68100 35022 68152 35028
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 68112 34785 68140 35022
rect 68098 34776 68154 34785
rect 68098 34711 68154 34720
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 65654 34300 65962 34309
rect 65654 34298 65660 34300
rect 65716 34298 65740 34300
rect 65796 34298 65820 34300
rect 65876 34298 65900 34300
rect 65956 34298 65962 34300
rect 65716 34246 65718 34298
rect 65898 34246 65900 34298
rect 65654 34244 65660 34246
rect 65716 34244 65740 34246
rect 65796 34244 65820 34246
rect 65876 34244 65900 34246
rect 65956 34244 65962 34246
rect 65654 34235 65962 34244
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 67638 33416 67694 33425
rect 67638 33351 67640 33360
rect 67692 33351 67694 33360
rect 67640 33322 67692 33328
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 65654 33212 65962 33221
rect 65654 33210 65660 33212
rect 65716 33210 65740 33212
rect 65796 33210 65820 33212
rect 65876 33210 65900 33212
rect 65956 33210 65962 33212
rect 65716 33158 65718 33210
rect 65898 33158 65900 33210
rect 65654 33156 65660 33158
rect 65716 33156 65740 33158
rect 65796 33156 65820 33158
rect 65876 33156 65900 33158
rect 65956 33156 65962 33158
rect 65654 33147 65962 33156
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 21364 32224 21416 32230
rect 21364 32166 21416 32172
rect 22468 32224 22520 32230
rect 22468 32166 22520 32172
rect 67640 32224 67692 32230
rect 67640 32166 67692 32172
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 21376 31890 21404 32166
rect 21824 32020 21876 32026
rect 21824 31962 21876 31968
rect 21364 31884 21416 31890
rect 21364 31826 21416 31832
rect 15108 31748 15160 31754
rect 15108 31690 15160 31696
rect 15292 31748 15344 31754
rect 15292 31690 15344 31696
rect 21364 31748 21416 31754
rect 21364 31690 21416 31696
rect 12624 31408 12676 31414
rect 12624 31350 12676 31356
rect 3424 31340 3476 31346
rect 3424 31282 3476 31288
rect 12440 31340 12492 31346
rect 12440 31282 12492 31288
rect 2872 31136 2924 31142
rect 2872 31078 2924 31084
rect 1676 30320 1728 30326
rect 1676 30262 1728 30268
rect 1688 28558 1716 30262
rect 2688 30252 2740 30258
rect 2688 30194 2740 30200
rect 2136 30048 2188 30054
rect 2136 29990 2188 29996
rect 2504 30048 2556 30054
rect 2504 29990 2556 29996
rect 2148 29646 2176 29990
rect 1952 29640 2004 29646
rect 1952 29582 2004 29588
rect 2136 29640 2188 29646
rect 2136 29582 2188 29588
rect 1964 29170 1992 29582
rect 2412 29572 2464 29578
rect 2412 29514 2464 29520
rect 2424 29306 2452 29514
rect 2412 29300 2464 29306
rect 2412 29242 2464 29248
rect 1952 29164 2004 29170
rect 1952 29106 2004 29112
rect 1676 28552 1728 28558
rect 1676 28494 1728 28500
rect 1688 27470 1716 28494
rect 1860 28484 1912 28490
rect 1860 28426 1912 28432
rect 1872 28218 1900 28426
rect 2044 28416 2096 28422
rect 2044 28358 2096 28364
rect 1860 28212 1912 28218
rect 1860 28154 1912 28160
rect 2056 28082 2084 28358
rect 2424 28150 2452 29242
rect 2516 29170 2544 29990
rect 2700 29578 2728 30194
rect 2884 30190 2912 31078
rect 2872 30184 2924 30190
rect 2872 30126 2924 30132
rect 3436 29850 3464 31282
rect 4804 31272 4856 31278
rect 4804 31214 4856 31220
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4816 30326 4844 31214
rect 6736 30728 6788 30734
rect 6736 30670 6788 30676
rect 11060 30728 11112 30734
rect 11060 30670 11112 30676
rect 6748 30326 6776 30670
rect 7104 30660 7156 30666
rect 7104 30602 7156 30608
rect 9220 30660 9272 30666
rect 9220 30602 9272 30608
rect 10968 30660 11020 30666
rect 10968 30602 11020 30608
rect 4804 30320 4856 30326
rect 4804 30262 4856 30268
rect 6736 30320 6788 30326
rect 6736 30262 6788 30268
rect 4712 30252 4764 30258
rect 4712 30194 4764 30200
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 3424 29844 3476 29850
rect 3424 29786 3476 29792
rect 2780 29776 2832 29782
rect 2780 29718 2832 29724
rect 2688 29572 2740 29578
rect 2688 29514 2740 29520
rect 2504 29164 2556 29170
rect 2504 29106 2556 29112
rect 2792 29034 2820 29718
rect 4160 29504 4212 29510
rect 4160 29446 4212 29452
rect 2596 29028 2648 29034
rect 2596 28970 2648 28976
rect 2688 29028 2740 29034
rect 2688 28970 2740 28976
rect 2780 29028 2832 29034
rect 4172 29016 4200 29446
rect 4724 29306 4752 30194
rect 4712 29300 4764 29306
rect 4712 29242 4764 29248
rect 4816 29238 4844 30262
rect 5814 30152 5870 30161
rect 6748 30122 6776 30262
rect 5814 30087 5816 30096
rect 5868 30087 5870 30096
rect 6736 30116 6788 30122
rect 5816 30058 5868 30064
rect 6736 30058 6788 30064
rect 5448 29572 5500 29578
rect 5448 29514 5500 29520
rect 4804 29232 4856 29238
rect 4804 29174 4856 29180
rect 4620 29164 4672 29170
rect 4620 29106 4672 29112
rect 2780 28970 2832 28976
rect 4080 28988 4200 29016
rect 2608 28558 2636 28970
rect 2596 28552 2648 28558
rect 2596 28494 2648 28500
rect 2412 28144 2464 28150
rect 2412 28086 2464 28092
rect 2044 28076 2096 28082
rect 2044 28018 2096 28024
rect 2608 28014 2636 28494
rect 2596 28008 2648 28014
rect 2596 27950 2648 27956
rect 2608 27470 2636 27950
rect 1676 27464 1728 27470
rect 1676 27406 1728 27412
rect 2320 27464 2372 27470
rect 2320 27406 2372 27412
rect 2596 27464 2648 27470
rect 2596 27406 2648 27412
rect 2136 27396 2188 27402
rect 2136 27338 2188 27344
rect 1676 27328 1728 27334
rect 1676 27270 1728 27276
rect 1688 25906 1716 27270
rect 2148 27130 2176 27338
rect 2332 27130 2360 27406
rect 2136 27124 2188 27130
rect 2136 27066 2188 27072
rect 2320 27124 2372 27130
rect 2320 27066 2372 27072
rect 2332 26994 2360 27066
rect 2320 26988 2372 26994
rect 2320 26930 2372 26936
rect 2608 26450 2636 27406
rect 2596 26444 2648 26450
rect 2596 26386 2648 26392
rect 1676 25900 1728 25906
rect 1676 25842 1728 25848
rect 1688 25158 1716 25842
rect 2412 25696 2464 25702
rect 2412 25638 2464 25644
rect 2320 25288 2372 25294
rect 2320 25230 2372 25236
rect 1676 25152 1728 25158
rect 1676 25094 1728 25100
rect 1688 24886 1716 25094
rect 1676 24880 1728 24886
rect 1676 24822 1728 24828
rect 1688 24138 1716 24822
rect 2332 24750 2360 25230
rect 2424 24818 2452 25638
rect 2700 25242 2728 28970
rect 4080 28694 4108 28988
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4632 28762 4660 29106
rect 5460 29073 5488 29514
rect 6644 29504 6696 29510
rect 6644 29446 6696 29452
rect 6656 29170 6684 29446
rect 7116 29306 7144 30602
rect 8116 30592 8168 30598
rect 8116 30534 8168 30540
rect 7748 30116 7800 30122
rect 7748 30058 7800 30064
rect 7288 29640 7340 29646
rect 7286 29608 7288 29617
rect 7340 29608 7342 29617
rect 7196 29572 7248 29578
rect 7286 29543 7342 29552
rect 7196 29514 7248 29520
rect 7104 29300 7156 29306
rect 7104 29242 7156 29248
rect 7208 29238 7236 29514
rect 7656 29504 7708 29510
rect 7656 29446 7708 29452
rect 7196 29232 7248 29238
rect 7196 29174 7248 29180
rect 6644 29164 6696 29170
rect 6644 29106 6696 29112
rect 6828 29164 6880 29170
rect 6828 29106 6880 29112
rect 5446 29064 5502 29073
rect 5446 28999 5448 29008
rect 5500 28999 5502 29008
rect 5448 28970 5500 28976
rect 4620 28756 4672 28762
rect 4620 28698 4672 28704
rect 4068 28688 4120 28694
rect 4068 28630 4120 28636
rect 5632 28620 5684 28626
rect 5632 28562 5684 28568
rect 3332 28484 3384 28490
rect 3332 28426 3384 28432
rect 3344 28150 3372 28426
rect 3332 28144 3384 28150
rect 3332 28086 3384 28092
rect 5080 28144 5132 28150
rect 5080 28086 5132 28092
rect 3148 28076 3200 28082
rect 3148 28018 3200 28024
rect 2872 27872 2924 27878
rect 2872 27814 2924 27820
rect 2884 27674 2912 27814
rect 2872 27668 2924 27674
rect 2872 27610 2924 27616
rect 3056 27396 3108 27402
rect 3056 27338 3108 27344
rect 3068 27130 3096 27338
rect 3056 27124 3108 27130
rect 3056 27066 3108 27072
rect 3056 26308 3108 26314
rect 3056 26250 3108 26256
rect 2964 25900 3016 25906
rect 2964 25842 3016 25848
rect 2872 25696 2924 25702
rect 2872 25638 2924 25644
rect 2884 25430 2912 25638
rect 2976 25498 3004 25842
rect 2964 25492 3016 25498
rect 2964 25434 3016 25440
rect 2872 25424 2924 25430
rect 2872 25366 2924 25372
rect 2608 25214 2728 25242
rect 2504 25152 2556 25158
rect 2504 25094 2556 25100
rect 2516 24818 2544 25094
rect 2412 24812 2464 24818
rect 2412 24754 2464 24760
rect 2504 24812 2556 24818
rect 2504 24754 2556 24760
rect 2320 24744 2372 24750
rect 2320 24686 2372 24692
rect 1676 24132 1728 24138
rect 1676 24074 1728 24080
rect 1688 22030 1716 24074
rect 1952 24064 2004 24070
rect 1952 24006 2004 24012
rect 1964 23186 1992 24006
rect 2332 23662 2360 24686
rect 2516 24342 2544 24754
rect 2504 24336 2556 24342
rect 2504 24278 2556 24284
rect 2320 23656 2372 23662
rect 2320 23598 2372 23604
rect 1952 23180 2004 23186
rect 1952 23122 2004 23128
rect 2332 23118 2360 23598
rect 2608 23322 2636 25214
rect 3068 24750 3096 26250
rect 3056 24744 3108 24750
rect 3056 24686 3108 24692
rect 2780 24064 2832 24070
rect 2780 24006 2832 24012
rect 2792 23662 2820 24006
rect 2780 23656 2832 23662
rect 2780 23598 2832 23604
rect 2412 23316 2464 23322
rect 2412 23258 2464 23264
rect 2596 23316 2648 23322
rect 2596 23258 2648 23264
rect 1860 23112 1912 23118
rect 1860 23054 1912 23060
rect 2320 23112 2372 23118
rect 2320 23054 2372 23060
rect 1676 22024 1728 22030
rect 1676 21966 1728 21972
rect 1872 21350 1900 23054
rect 2044 23044 2096 23050
rect 2044 22986 2096 22992
rect 2056 22642 2084 22986
rect 2332 22710 2360 23054
rect 2320 22704 2372 22710
rect 2320 22646 2372 22652
rect 1952 22636 2004 22642
rect 1952 22578 2004 22584
rect 2044 22636 2096 22642
rect 2044 22578 2096 22584
rect 1964 22234 1992 22578
rect 1952 22228 2004 22234
rect 1952 22170 2004 22176
rect 1860 21344 1912 21350
rect 1860 21286 1912 21292
rect 2320 20936 2372 20942
rect 2320 20878 2372 20884
rect 1952 20460 2004 20466
rect 1952 20402 2004 20408
rect 2136 20460 2188 20466
rect 2136 20402 2188 20408
rect 1964 20369 1992 20402
rect 1950 20360 2006 20369
rect 1950 20295 2006 20304
rect 2044 20256 2096 20262
rect 2044 20198 2096 20204
rect 2056 19854 2084 20198
rect 1860 19848 1912 19854
rect 1860 19790 1912 19796
rect 2044 19848 2096 19854
rect 2044 19790 2096 19796
rect 1872 19378 1900 19790
rect 2148 19417 2176 20402
rect 2332 19990 2360 20878
rect 2320 19984 2372 19990
rect 2320 19926 2372 19932
rect 2424 19854 2452 23258
rect 2504 22772 2556 22778
rect 2504 22714 2556 22720
rect 2516 22642 2544 22714
rect 2504 22636 2556 22642
rect 2504 22578 2556 22584
rect 2516 21894 2544 22578
rect 2504 21888 2556 21894
rect 2504 21830 2556 21836
rect 2412 19848 2464 19854
rect 2412 19790 2464 19796
rect 2228 19712 2280 19718
rect 2228 19654 2280 19660
rect 2240 19446 2268 19654
rect 2424 19514 2452 19790
rect 2412 19508 2464 19514
rect 2412 19450 2464 19456
rect 2228 19440 2280 19446
rect 2134 19408 2190 19417
rect 1860 19372 1912 19378
rect 2228 19382 2280 19388
rect 2134 19343 2190 19352
rect 1860 19314 1912 19320
rect 1872 18290 1900 19314
rect 2148 18766 2176 19343
rect 2136 18760 2188 18766
rect 2136 18702 2188 18708
rect 1860 18284 1912 18290
rect 1860 18226 1912 18232
rect 2044 18284 2096 18290
rect 2044 18226 2096 18232
rect 2136 18284 2188 18290
rect 2240 18272 2268 19382
rect 2320 19372 2372 19378
rect 2320 19314 2372 19320
rect 2332 18970 2360 19314
rect 2320 18964 2372 18970
rect 2320 18906 2372 18912
rect 2188 18244 2268 18272
rect 2136 18226 2188 18232
rect 2056 17746 2084 18226
rect 2044 17740 2096 17746
rect 2044 17682 2096 17688
rect 1858 17232 1914 17241
rect 1858 17167 1860 17176
rect 1912 17167 1914 17176
rect 1860 17138 1912 17144
rect 1872 15502 1900 17138
rect 2044 16584 2096 16590
rect 2044 16526 2096 16532
rect 2056 16114 2084 16526
rect 2044 16108 2096 16114
rect 2044 16050 2096 16056
rect 1860 15496 1912 15502
rect 1860 15438 1912 15444
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 1964 14414 1992 14758
rect 1768 14408 1820 14414
rect 1768 14350 1820 14356
rect 1952 14408 2004 14414
rect 1952 14350 2004 14356
rect 1780 13870 1808 14350
rect 1768 13864 1820 13870
rect 1768 13806 1820 13812
rect 1780 11762 1808 13806
rect 2056 12306 2084 16050
rect 2148 14550 2176 18226
rect 2424 17338 2452 19450
rect 2412 17332 2464 17338
rect 2412 17274 2464 17280
rect 2320 17264 2372 17270
rect 2320 17206 2372 17212
rect 2228 16992 2280 16998
rect 2228 16934 2280 16940
rect 2240 16590 2268 16934
rect 2228 16584 2280 16590
rect 2228 16526 2280 16532
rect 2332 16454 2360 17206
rect 2320 16448 2372 16454
rect 2320 16390 2372 16396
rect 2332 16114 2360 16390
rect 2228 16108 2280 16114
rect 2228 16050 2280 16056
rect 2320 16108 2372 16114
rect 2320 16050 2372 16056
rect 2240 15706 2268 16050
rect 2228 15700 2280 15706
rect 2228 15642 2280 15648
rect 2136 14544 2188 14550
rect 2136 14486 2188 14492
rect 2228 14544 2280 14550
rect 2228 14486 2280 14492
rect 2240 14414 2268 14486
rect 2228 14408 2280 14414
rect 2228 14350 2280 14356
rect 2516 13433 2544 21830
rect 2596 21344 2648 21350
rect 2596 21286 2648 21292
rect 2502 13424 2558 13433
rect 2502 13359 2558 13368
rect 2228 13252 2280 13258
rect 2228 13194 2280 13200
rect 2320 13252 2372 13258
rect 2320 13194 2372 13200
rect 2136 13184 2188 13190
rect 2136 13126 2188 13132
rect 2044 12300 2096 12306
rect 2044 12242 2096 12248
rect 2148 12238 2176 13126
rect 2240 12986 2268 13194
rect 2228 12980 2280 12986
rect 2228 12922 2280 12928
rect 2228 12776 2280 12782
rect 2228 12718 2280 12724
rect 2240 12238 2268 12718
rect 2332 12374 2360 13194
rect 2320 12368 2372 12374
rect 2320 12310 2372 12316
rect 2136 12232 2188 12238
rect 2136 12174 2188 12180
rect 2228 12232 2280 12238
rect 2228 12174 2280 12180
rect 2240 11762 2268 12174
rect 1768 11756 1820 11762
rect 1768 11698 1820 11704
rect 2136 11756 2188 11762
rect 2136 11698 2188 11704
rect 2228 11756 2280 11762
rect 2228 11698 2280 11704
rect 1780 10674 1808 11698
rect 2148 11354 2176 11698
rect 2136 11348 2188 11354
rect 2136 11290 2188 11296
rect 2240 10742 2268 11698
rect 2332 11082 2360 12310
rect 2516 12238 2544 13359
rect 2504 12232 2556 12238
rect 2504 12174 2556 12180
rect 2504 11552 2556 11558
rect 2504 11494 2556 11500
rect 2516 11150 2544 11494
rect 2504 11144 2556 11150
rect 2504 11086 2556 11092
rect 2320 11076 2372 11082
rect 2372 11036 2452 11064
rect 2320 11018 2372 11024
rect 2228 10736 2280 10742
rect 2280 10696 2360 10724
rect 2228 10678 2280 10684
rect 1768 10668 1820 10674
rect 1768 10610 1820 10616
rect 1860 10668 1912 10674
rect 1860 10610 1912 10616
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 1780 9586 1808 10610
rect 1872 10266 1900 10610
rect 2044 10464 2096 10470
rect 2044 10406 2096 10412
rect 1860 10260 1912 10266
rect 1860 10202 1912 10208
rect 2056 10062 2084 10406
rect 2148 10198 2176 10610
rect 2136 10192 2188 10198
rect 2136 10134 2188 10140
rect 2044 10056 2096 10062
rect 2044 9998 2096 10004
rect 1768 9580 1820 9586
rect 1768 9522 1820 9528
rect 1780 8974 1808 9522
rect 2332 9450 2360 10696
rect 2424 10062 2452 11036
rect 2412 10056 2464 10062
rect 2412 9998 2464 10004
rect 2320 9444 2372 9450
rect 2320 9386 2372 9392
rect 2332 9042 2360 9386
rect 2412 9376 2464 9382
rect 2412 9318 2464 9324
rect 2320 9036 2372 9042
rect 2320 8978 2372 8984
rect 1768 8968 1820 8974
rect 1768 8910 1820 8916
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 1860 7744 1912 7750
rect 1860 7686 1912 7692
rect 1768 6860 1820 6866
rect 1768 6802 1820 6808
rect 1780 6322 1808 6802
rect 1872 6798 1900 7686
rect 1860 6792 1912 6798
rect 1860 6734 1912 6740
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 1400 4616 1452 4622
rect 1400 4558 1452 4564
rect 1412 3194 1440 4558
rect 1780 4078 1808 6258
rect 1952 6112 2004 6118
rect 1952 6054 2004 6060
rect 1964 5710 1992 6054
rect 1952 5704 2004 5710
rect 1952 5646 2004 5652
rect 1952 4480 2004 4486
rect 1952 4422 2004 4428
rect 1964 4146 1992 4422
rect 2056 4162 2084 8434
rect 2320 7948 2372 7954
rect 2320 7890 2372 7896
rect 2136 7404 2188 7410
rect 2136 7346 2188 7352
rect 2148 7002 2176 7346
rect 2136 6996 2188 7002
rect 2136 6938 2188 6944
rect 2332 6390 2360 7890
rect 2424 6914 2452 9318
rect 2608 8090 2636 21286
rect 2792 20942 2820 23598
rect 2872 23112 2924 23118
rect 2872 23054 2924 23060
rect 2884 22642 2912 23054
rect 3056 22976 3108 22982
rect 3056 22918 3108 22924
rect 2872 22636 2924 22642
rect 2872 22578 2924 22584
rect 2884 21622 2912 22578
rect 3068 22098 3096 22918
rect 3056 22094 3108 22098
rect 2976 22092 3108 22094
rect 2976 22066 3056 22092
rect 2872 21616 2924 21622
rect 2872 21558 2924 21564
rect 2780 20936 2832 20942
rect 2780 20878 2832 20884
rect 2792 19922 2820 20878
rect 2884 20534 2912 21558
rect 2872 20528 2924 20534
rect 2872 20470 2924 20476
rect 2780 19916 2832 19922
rect 2780 19858 2832 19864
rect 2688 19508 2740 19514
rect 2688 19450 2740 19456
rect 2700 18290 2728 19450
rect 2976 19334 3004 22066
rect 3056 22034 3108 22040
rect 3068 21983 3096 22034
rect 3160 21690 3188 28018
rect 3344 27538 3372 28086
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 3332 27532 3384 27538
rect 3332 27474 3384 27480
rect 3344 26994 3372 27474
rect 5092 27470 5120 28086
rect 5080 27464 5132 27470
rect 5080 27406 5132 27412
rect 5448 27464 5500 27470
rect 5448 27406 5500 27412
rect 4436 27328 4488 27334
rect 4436 27270 4488 27276
rect 4448 27062 4476 27270
rect 4436 27056 4488 27062
rect 4436 26998 4488 27004
rect 3332 26988 3384 26994
rect 3332 26930 3384 26936
rect 3608 26920 3660 26926
rect 3608 26862 3660 26868
rect 4068 26920 4120 26926
rect 4068 26862 4120 26868
rect 3240 24880 3292 24886
rect 3240 24822 3292 24828
rect 3252 23730 3280 24822
rect 3332 24336 3384 24342
rect 3332 24278 3384 24284
rect 3344 23730 3372 24278
rect 3620 24274 3648 26862
rect 4080 26466 4108 26862
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4080 26438 4292 26466
rect 4264 26382 4292 26438
rect 3884 26376 3936 26382
rect 3884 26318 3936 26324
rect 4252 26376 4304 26382
rect 4252 26318 4304 26324
rect 3700 24812 3752 24818
rect 3700 24754 3752 24760
rect 3712 24410 3740 24754
rect 3700 24404 3752 24410
rect 3700 24346 3752 24352
rect 3608 24268 3660 24274
rect 3608 24210 3660 24216
rect 3240 23724 3292 23730
rect 3240 23666 3292 23672
rect 3332 23724 3384 23730
rect 3332 23666 3384 23672
rect 3344 23186 3372 23666
rect 3712 23594 3740 24346
rect 3896 24138 3924 26318
rect 4264 25906 4292 26318
rect 4252 25900 4304 25906
rect 4252 25842 4304 25848
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4068 24812 4120 24818
rect 4068 24754 4120 24760
rect 3976 24268 4028 24274
rect 3976 24210 4028 24216
rect 3884 24132 3936 24138
rect 3884 24074 3936 24080
rect 3700 23588 3752 23594
rect 3700 23530 3752 23536
rect 3884 23520 3936 23526
rect 3884 23462 3936 23468
rect 3332 23180 3384 23186
rect 3332 23122 3384 23128
rect 3896 22982 3924 23462
rect 3884 22976 3936 22982
rect 3884 22918 3936 22924
rect 3988 22710 4016 24210
rect 4080 23866 4108 24754
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4068 23860 4120 23866
rect 4068 23802 4120 23808
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 3976 22704 4028 22710
rect 3976 22646 4028 22652
rect 3884 21888 3936 21894
rect 3884 21830 3936 21836
rect 3148 21684 3200 21690
rect 3148 21626 3200 21632
rect 3056 20460 3108 20466
rect 3056 20402 3108 20408
rect 3068 20058 3096 20402
rect 3160 20058 3188 21626
rect 3896 21554 3924 21830
rect 3988 21690 4016 22646
rect 4618 22536 4674 22545
rect 4618 22471 4620 22480
rect 4672 22471 4674 22480
rect 4620 22442 4672 22448
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4632 22030 4660 22442
rect 4712 22432 4764 22438
rect 4712 22374 4764 22380
rect 4620 22024 4672 22030
rect 4620 21966 4672 21972
rect 3976 21684 4028 21690
rect 3976 21626 4028 21632
rect 4724 21622 4752 22374
rect 5092 22137 5120 27406
rect 5356 26988 5408 26994
rect 5356 26930 5408 26936
rect 5172 24200 5224 24206
rect 5172 24142 5224 24148
rect 5184 23089 5212 24142
rect 5368 23882 5396 26930
rect 5460 26382 5488 27406
rect 5448 26376 5500 26382
rect 5448 26318 5500 26324
rect 5460 25294 5488 26318
rect 5448 25288 5500 25294
rect 5448 25230 5500 25236
rect 5460 24886 5488 25230
rect 5448 24880 5500 24886
rect 5448 24822 5500 24828
rect 5540 24880 5592 24886
rect 5540 24822 5592 24828
rect 5276 23866 5396 23882
rect 5276 23860 5408 23866
rect 5276 23854 5356 23860
rect 5170 23080 5226 23089
rect 5170 23015 5226 23024
rect 5184 22982 5212 23015
rect 5172 22976 5224 22982
rect 5172 22918 5224 22924
rect 5172 22636 5224 22642
rect 5172 22578 5224 22584
rect 5184 22234 5212 22578
rect 5172 22228 5224 22234
rect 5172 22170 5224 22176
rect 5078 22128 5134 22137
rect 5276 22098 5304 23854
rect 5356 23802 5408 23808
rect 5552 23798 5580 24822
rect 5540 23792 5592 23798
rect 5540 23734 5592 23740
rect 5644 23254 5672 28562
rect 6840 28422 6868 29106
rect 7012 29028 7064 29034
rect 7012 28970 7064 28976
rect 7024 28626 7052 28970
rect 7012 28620 7064 28626
rect 7012 28562 7064 28568
rect 7208 28558 7236 29174
rect 7380 29096 7432 29102
rect 7380 29038 7432 29044
rect 7196 28552 7248 28558
rect 7196 28494 7248 28500
rect 7012 28484 7064 28490
rect 7012 28426 7064 28432
rect 5908 28416 5960 28422
rect 5908 28358 5960 28364
rect 6828 28416 6880 28422
rect 6828 28358 6880 28364
rect 5816 26580 5868 26586
rect 5816 26522 5868 26528
rect 5828 25974 5856 26522
rect 5816 25968 5868 25974
rect 5816 25910 5868 25916
rect 5724 24064 5776 24070
rect 5724 24006 5776 24012
rect 5736 23730 5764 24006
rect 5724 23724 5776 23730
rect 5724 23666 5776 23672
rect 5632 23248 5684 23254
rect 5632 23190 5684 23196
rect 5356 22636 5408 22642
rect 5356 22578 5408 22584
rect 5078 22063 5134 22072
rect 5264 22092 5316 22098
rect 4712 21616 4764 21622
rect 4712 21558 4764 21564
rect 3332 21548 3384 21554
rect 3332 21490 3384 21496
rect 3884 21548 3936 21554
rect 3884 21490 3936 21496
rect 4068 21548 4120 21554
rect 4068 21490 4120 21496
rect 3240 21344 3292 21350
rect 3240 21286 3292 21292
rect 3056 20052 3108 20058
rect 3056 19994 3108 20000
rect 3148 20052 3200 20058
rect 3148 19994 3200 20000
rect 3056 19916 3108 19922
rect 3056 19858 3108 19864
rect 2884 19306 3004 19334
rect 2688 18284 2740 18290
rect 2688 18226 2740 18232
rect 2700 17882 2728 18226
rect 2688 17876 2740 17882
rect 2688 17818 2740 17824
rect 2700 16114 2728 17818
rect 2688 16108 2740 16114
rect 2688 16050 2740 16056
rect 2688 15904 2740 15910
rect 2688 15846 2740 15852
rect 2700 15570 2728 15846
rect 2688 15564 2740 15570
rect 2688 15506 2740 15512
rect 2780 14272 2832 14278
rect 2780 14214 2832 14220
rect 2792 13938 2820 14214
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 2884 13682 2912 19306
rect 3068 13734 3096 19858
rect 3252 19378 3280 21286
rect 3344 20806 3372 21490
rect 3332 20800 3384 20806
rect 3332 20742 3384 20748
rect 3240 19372 3292 19378
rect 3240 19314 3292 19320
rect 3252 18970 3280 19314
rect 3240 18964 3292 18970
rect 3240 18906 3292 18912
rect 3252 16794 3280 18906
rect 3240 16788 3292 16794
rect 3240 16730 3292 16736
rect 3252 16590 3280 16730
rect 3240 16584 3292 16590
rect 3240 16526 3292 16532
rect 3148 15496 3200 15502
rect 3148 15438 3200 15444
rect 3160 14006 3188 15438
rect 3148 14000 3200 14006
rect 3148 13942 3200 13948
rect 2792 13654 2912 13682
rect 3056 13728 3108 13734
rect 3056 13670 3108 13676
rect 2792 12170 2820 13654
rect 3068 13530 3096 13670
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 3056 13524 3108 13530
rect 3056 13466 3108 13472
rect 2884 12434 2912 13466
rect 3160 13394 3188 13942
rect 3148 13388 3200 13394
rect 3148 13330 3200 13336
rect 3160 12850 3188 13330
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 3240 12844 3292 12850
rect 3240 12786 3292 12792
rect 3252 12442 3280 12786
rect 3240 12436 3292 12442
rect 2884 12406 3004 12434
rect 2780 12164 2832 12170
rect 2780 12106 2832 12112
rect 2792 11762 2820 12106
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2792 11354 2820 11698
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2976 9674 3004 12406
rect 3240 12378 3292 12384
rect 3148 11688 3200 11694
rect 3148 11630 3200 11636
rect 3160 11150 3188 11630
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 3160 10674 3188 11086
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3240 10668 3292 10674
rect 3240 10610 3292 10616
rect 2976 9646 3188 9674
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 2700 8566 2728 9318
rect 3160 8786 3188 9646
rect 3252 9178 3280 10610
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 3160 8758 3280 8786
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 2688 8560 2740 8566
rect 2688 8502 2740 8508
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2596 8084 2648 8090
rect 2596 8026 2648 8032
rect 2872 8084 2924 8090
rect 2872 8026 2924 8032
rect 2608 7886 2636 8026
rect 2688 8016 2740 8022
rect 2688 7958 2740 7964
rect 2596 7880 2648 7886
rect 2596 7822 2648 7828
rect 2700 7342 2728 7958
rect 2884 7750 2912 8026
rect 2872 7744 2924 7750
rect 2872 7686 2924 7692
rect 2976 7342 3004 8230
rect 2688 7336 2740 7342
rect 2688 7278 2740 7284
rect 2964 7336 3016 7342
rect 2964 7278 3016 7284
rect 2424 6886 2544 6914
rect 2320 6384 2372 6390
rect 2320 6326 2372 6332
rect 2228 5228 2280 5234
rect 2228 5170 2280 5176
rect 2240 4282 2268 5170
rect 2332 4690 2360 6326
rect 2320 4684 2372 4690
rect 2320 4626 2372 4632
rect 2228 4276 2280 4282
rect 2228 4218 2280 4224
rect 1952 4140 2004 4146
rect 2056 4134 2268 4162
rect 1952 4082 2004 4088
rect 1768 4072 1820 4078
rect 1768 4014 1820 4020
rect 1952 3936 2004 3942
rect 1952 3878 2004 3884
rect 1768 3392 1820 3398
rect 1768 3334 1820 3340
rect 1400 3188 1452 3194
rect 1400 3130 1452 3136
rect 1780 3058 1808 3334
rect 1964 3058 1992 3878
rect 2240 3398 2268 4134
rect 2332 3602 2360 4626
rect 2412 4480 2464 4486
rect 2412 4422 2464 4428
rect 2320 3596 2372 3602
rect 2320 3538 2372 3544
rect 2228 3392 2280 3398
rect 2226 3360 2228 3369
rect 2280 3360 2282 3369
rect 2226 3295 2282 3304
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 1952 3052 2004 3058
rect 1952 2994 2004 3000
rect 1768 2440 1820 2446
rect 2424 2417 2452 4422
rect 2516 2446 2544 6886
rect 2700 4486 2728 7278
rect 2976 6390 3004 7278
rect 2964 6384 3016 6390
rect 2964 6326 3016 6332
rect 3056 6316 3108 6322
rect 3056 6258 3108 6264
rect 3068 5914 3096 6258
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 2964 5024 3016 5030
rect 2964 4966 3016 4972
rect 2780 4752 2832 4758
rect 2780 4694 2832 4700
rect 2688 4480 2740 4486
rect 2688 4422 2740 4428
rect 2792 3074 2820 4694
rect 2976 4214 3004 4966
rect 2964 4208 3016 4214
rect 2964 4150 3016 4156
rect 2872 4072 2924 4078
rect 2924 4032 3004 4060
rect 2872 4014 2924 4020
rect 2976 3126 3004 4032
rect 3056 3936 3108 3942
rect 3056 3878 3108 3884
rect 3068 3534 3096 3878
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 2964 3120 3016 3126
rect 2792 3058 2912 3074
rect 2964 3062 3016 3068
rect 2792 3052 2924 3058
rect 2792 3046 2872 3052
rect 2872 2994 2924 3000
rect 3160 2774 3188 8570
rect 3252 5914 3280 8758
rect 3344 8022 3372 20742
rect 3424 19372 3476 19378
rect 3424 19314 3476 19320
rect 3436 18358 3464 19314
rect 3424 18352 3476 18358
rect 3424 18294 3476 18300
rect 3792 16584 3844 16590
rect 3792 16526 3844 16532
rect 3804 15502 3832 16526
rect 3792 15496 3844 15502
rect 3792 15438 3844 15444
rect 3804 15162 3832 15438
rect 3792 15156 3844 15162
rect 3792 15098 3844 15104
rect 3792 14408 3844 14414
rect 3792 14350 3844 14356
rect 3804 12918 3832 14350
rect 3792 12912 3844 12918
rect 3792 12854 3844 12860
rect 3792 10056 3844 10062
rect 3792 9998 3844 10004
rect 3804 8906 3832 9998
rect 3792 8900 3844 8906
rect 3792 8842 3844 8848
rect 3896 8498 3924 21490
rect 4080 21010 4108 21490
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4068 21004 4120 21010
rect 4068 20946 4120 20952
rect 4080 19922 4108 20946
rect 4712 20460 4764 20466
rect 4764 20420 4844 20448
rect 4712 20402 4764 20408
rect 4158 20360 4214 20369
rect 4158 20295 4160 20304
rect 4212 20295 4214 20304
rect 4160 20266 4212 20272
rect 4620 20256 4672 20262
rect 4620 20198 4672 20204
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4344 19984 4396 19990
rect 4344 19926 4396 19932
rect 4068 19916 4120 19922
rect 4068 19858 4120 19864
rect 4080 19378 4108 19858
rect 4356 19854 4384 19926
rect 4344 19848 4396 19854
rect 4344 19790 4396 19796
rect 4528 19848 4580 19854
rect 4632 19836 4660 20198
rect 4580 19808 4660 19836
rect 4528 19790 4580 19796
rect 4816 19417 4844 20420
rect 5092 19854 5120 22063
rect 5264 22034 5316 22040
rect 5264 20324 5316 20330
rect 5264 20266 5316 20272
rect 5080 19848 5132 19854
rect 5080 19790 5132 19796
rect 4802 19408 4858 19417
rect 4068 19372 4120 19378
rect 4802 19343 4858 19352
rect 4068 19314 4120 19320
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4620 18080 4672 18086
rect 4620 18022 4672 18028
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4632 17678 4660 18022
rect 4620 17672 4672 17678
rect 4620 17614 4672 17620
rect 4816 17610 4844 19343
rect 5172 19168 5224 19174
rect 5172 19110 5224 19116
rect 4988 18760 5040 18766
rect 4988 18702 5040 18708
rect 4804 17604 4856 17610
rect 4804 17546 4856 17552
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4816 15094 4844 17546
rect 5000 17134 5028 18702
rect 5184 18698 5212 19110
rect 5172 18692 5224 18698
rect 5172 18634 5224 18640
rect 5080 17196 5132 17202
rect 5080 17138 5132 17144
rect 4988 17128 5040 17134
rect 4908 17088 4988 17116
rect 4908 15978 4936 17088
rect 4988 17070 5040 17076
rect 5092 16794 5120 17138
rect 5080 16788 5132 16794
rect 5080 16730 5132 16736
rect 4988 16108 5040 16114
rect 5092 16096 5120 16730
rect 5184 16182 5212 18634
rect 5276 16454 5304 20266
rect 5368 19990 5396 22578
rect 5644 20534 5672 23190
rect 5920 22094 5948 28358
rect 6828 28212 6880 28218
rect 6828 28154 6880 28160
rect 6840 27334 6868 28154
rect 7024 28014 7052 28426
rect 7012 28008 7064 28014
rect 7012 27950 7064 27956
rect 6828 27328 6880 27334
rect 6828 27270 6880 27276
rect 7024 26450 7052 27950
rect 7208 27878 7236 28494
rect 7392 28490 7420 29038
rect 7668 28558 7696 29446
rect 7760 29170 7788 30058
rect 8128 29617 8156 30534
rect 8114 29608 8170 29617
rect 9232 29578 9260 30602
rect 9772 30592 9824 30598
rect 9772 30534 9824 30540
rect 9312 30252 9364 30258
rect 9312 30194 9364 30200
rect 8114 29543 8170 29552
rect 9220 29572 9272 29578
rect 9220 29514 9272 29520
rect 9128 29504 9180 29510
rect 9128 29446 9180 29452
rect 7748 29164 7800 29170
rect 7748 29106 7800 29112
rect 8024 29164 8076 29170
rect 8024 29106 8076 29112
rect 8036 28762 8064 29106
rect 9140 29034 9168 29446
rect 9128 29028 9180 29034
rect 9128 28970 9180 28976
rect 8024 28756 8076 28762
rect 8024 28698 8076 28704
rect 7656 28552 7708 28558
rect 7656 28494 7708 28500
rect 7380 28484 7432 28490
rect 7380 28426 7432 28432
rect 7656 28076 7708 28082
rect 7656 28018 7708 28024
rect 7564 28008 7616 28014
rect 7564 27950 7616 27956
rect 7196 27872 7248 27878
rect 7196 27814 7248 27820
rect 7104 26920 7156 26926
rect 7104 26862 7156 26868
rect 7012 26444 7064 26450
rect 7012 26386 7064 26392
rect 7012 25220 7064 25226
rect 7012 25162 7064 25168
rect 6276 24744 6328 24750
rect 6276 24686 6328 24692
rect 6288 24138 6316 24686
rect 7024 24410 7052 25162
rect 7116 24410 7144 26862
rect 7012 24404 7064 24410
rect 7012 24346 7064 24352
rect 7104 24404 7156 24410
rect 7104 24346 7156 24352
rect 6276 24132 6328 24138
rect 6276 24074 6328 24080
rect 7012 24132 7064 24138
rect 7012 24074 7064 24080
rect 6092 23044 6144 23050
rect 6092 22986 6144 22992
rect 5736 22066 5948 22094
rect 5736 21350 5764 22066
rect 5816 21956 5868 21962
rect 5816 21898 5868 21904
rect 5828 21418 5856 21898
rect 6104 21894 6132 22986
rect 6288 22098 6316 24074
rect 6828 23792 6880 23798
rect 6828 23734 6880 23740
rect 6460 23656 6512 23662
rect 6460 23598 6512 23604
rect 6368 23112 6420 23118
rect 6368 23054 6420 23060
rect 6276 22092 6328 22098
rect 6276 22034 6328 22040
rect 6092 21888 6144 21894
rect 6092 21830 6144 21836
rect 5816 21412 5868 21418
rect 5816 21354 5868 21360
rect 5724 21344 5776 21350
rect 5724 21286 5776 21292
rect 5736 21146 5764 21286
rect 5724 21140 5776 21146
rect 5724 21082 5776 21088
rect 5632 20528 5684 20534
rect 5632 20470 5684 20476
rect 5356 19984 5408 19990
rect 5356 19926 5408 19932
rect 5644 19514 5672 20470
rect 5632 19508 5684 19514
rect 5632 19450 5684 19456
rect 5356 17672 5408 17678
rect 5356 17614 5408 17620
rect 5264 16448 5316 16454
rect 5264 16390 5316 16396
rect 5172 16176 5224 16182
rect 5172 16118 5224 16124
rect 5040 16068 5120 16096
rect 4988 16050 5040 16056
rect 4896 15972 4948 15978
rect 4896 15914 4948 15920
rect 5264 15972 5316 15978
rect 5264 15914 5316 15920
rect 4804 15088 4856 15094
rect 4804 15030 4856 15036
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 4080 14822 4108 14962
rect 4068 14816 4120 14822
rect 4068 14758 4120 14764
rect 4080 14074 4108 14758
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 4620 14000 4672 14006
rect 4620 13942 4672 13948
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4632 13326 4660 13942
rect 4816 13938 4844 15030
rect 4908 14414 4936 15914
rect 5080 15428 5132 15434
rect 5080 15370 5132 15376
rect 5092 15026 5120 15370
rect 5276 15366 5304 15914
rect 5264 15360 5316 15366
rect 5264 15302 5316 15308
rect 5276 15026 5304 15302
rect 5368 15094 5396 17614
rect 5446 16008 5502 16017
rect 5446 15943 5448 15952
rect 5500 15943 5502 15952
rect 5448 15914 5500 15920
rect 5356 15088 5408 15094
rect 5356 15030 5408 15036
rect 5080 15020 5132 15026
rect 5080 14962 5132 14968
rect 5264 15020 5316 15026
rect 5264 14962 5316 14968
rect 5630 14920 5686 14929
rect 5630 14855 5632 14864
rect 5684 14855 5686 14864
rect 5724 14884 5776 14890
rect 5632 14826 5684 14832
rect 5724 14826 5776 14832
rect 5736 14414 5764 14826
rect 4896 14408 4948 14414
rect 4896 14350 4948 14356
rect 5264 14408 5316 14414
rect 5264 14350 5316 14356
rect 5724 14408 5776 14414
rect 5724 14350 5776 14356
rect 4804 13932 4856 13938
rect 4804 13874 4856 13880
rect 5276 13530 5304 14350
rect 5724 14272 5776 14278
rect 5724 14214 5776 14220
rect 5264 13524 5316 13530
rect 5264 13466 5316 13472
rect 5736 13326 5764 14214
rect 5908 13728 5960 13734
rect 5908 13670 5960 13676
rect 4620 13320 4672 13326
rect 4620 13262 4672 13268
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4632 12238 4660 13262
rect 5264 13184 5316 13190
rect 5264 13126 5316 13132
rect 5276 12986 5304 13126
rect 5264 12980 5316 12986
rect 5264 12922 5316 12928
rect 5816 12980 5868 12986
rect 5816 12922 5868 12928
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 5172 11824 5224 11830
rect 5172 11766 5224 11772
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 5184 11354 5212 11766
rect 5828 11762 5856 12922
rect 5920 12442 5948 13670
rect 5908 12436 5960 12442
rect 5908 12378 5960 12384
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 4528 10804 4580 10810
rect 4528 10746 4580 10752
rect 4540 10470 4568 10746
rect 5828 10742 5856 11698
rect 5816 10736 5868 10742
rect 5816 10678 5868 10684
rect 4528 10464 4580 10470
rect 4528 10406 4580 10412
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 5828 10062 5856 10678
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 3976 9988 4028 9994
rect 3976 9930 4028 9936
rect 3988 8634 4016 9930
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 5448 9920 5500 9926
rect 5448 9862 5500 9868
rect 4172 9722 4200 9862
rect 4160 9716 4212 9722
rect 4160 9658 4212 9664
rect 5172 9686 5224 9692
rect 4620 9648 4672 9654
rect 5264 9648 5316 9654
rect 5224 9634 5264 9636
rect 5172 9628 5264 9634
rect 4620 9590 4672 9596
rect 5184 9608 5264 9628
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 4080 8838 4108 9522
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4632 8974 4660 9590
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 3976 8424 4028 8430
rect 3976 8366 4028 8372
rect 3332 8016 3384 8022
rect 3332 7958 3384 7964
rect 3332 7744 3384 7750
rect 3332 7686 3384 7692
rect 3240 5908 3292 5914
rect 3240 5850 3292 5856
rect 3252 5817 3280 5850
rect 3238 5808 3294 5817
rect 3238 5743 3294 5752
rect 2976 2746 3188 2774
rect 2976 2446 3004 2746
rect 2504 2440 2556 2446
rect 1768 2382 1820 2388
rect 2410 2408 2466 2417
rect 1780 1358 1808 2382
rect 2504 2382 2556 2388
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 2410 2343 2466 2352
rect 1768 1352 1820 1358
rect 1768 1294 1820 1300
rect 2516 202 2544 2382
rect 2976 1698 3004 2382
rect 3240 2304 3292 2310
rect 3344 2281 3372 7686
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 3804 4162 3832 5510
rect 3884 4616 3936 4622
rect 3884 4558 3936 4564
rect 3712 4146 3832 4162
rect 3700 4140 3832 4146
rect 3752 4134 3832 4140
rect 3700 4082 3752 4088
rect 3804 3602 3832 4134
rect 3896 3738 3924 4558
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3792 3596 3844 3602
rect 3792 3538 3844 3544
rect 3884 3528 3936 3534
rect 3988 3516 4016 8366
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 7886 4660 8910
rect 5184 8906 5212 9608
rect 5264 9590 5316 9596
rect 5460 8906 5488 9862
rect 5828 9586 5856 9998
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 5172 8900 5224 8906
rect 5172 8842 5224 8848
rect 5448 8900 5500 8906
rect 5448 8842 5500 8848
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4436 7812 4488 7818
rect 4436 7754 4488 7760
rect 4448 7546 4476 7754
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4632 6662 4660 7822
rect 4816 7546 4844 8434
rect 5092 8378 5120 8774
rect 5724 8560 5776 8566
rect 5724 8502 5776 8508
rect 5092 8350 5212 8378
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 5092 7886 5120 8230
rect 5080 7880 5132 7886
rect 5080 7822 5132 7828
rect 4896 7744 4948 7750
rect 4896 7686 4948 7692
rect 4804 7540 4856 7546
rect 4804 7482 4856 7488
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 4080 6254 4108 6394
rect 4632 6390 4660 6598
rect 4620 6384 4672 6390
rect 4620 6326 4672 6332
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4632 4554 4660 6326
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4724 4622 4752 4966
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4252 4548 4304 4554
rect 4252 4490 4304 4496
rect 4620 4548 4672 4554
rect 4620 4490 4672 4496
rect 4264 4049 4292 4490
rect 4250 4040 4306 4049
rect 4250 3975 4306 3984
rect 4264 3942 4292 3975
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 3936 3488 4016 3516
rect 3884 3470 3936 3476
rect 3988 3194 4016 3488
rect 4632 3194 4660 4490
rect 4712 4480 4764 4486
rect 4712 4422 4764 4428
rect 3976 3188 4028 3194
rect 3976 3130 4028 3136
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4724 3126 4752 4422
rect 4712 3120 4764 3126
rect 4712 3062 4764 3068
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4908 2446 4936 7686
rect 5080 6792 5132 6798
rect 5080 6734 5132 6740
rect 5092 4146 5120 6734
rect 5080 4140 5132 4146
rect 5080 4082 5132 4088
rect 5092 3777 5120 4082
rect 5078 3768 5134 3777
rect 5078 3703 5134 3712
rect 5184 2514 5212 8350
rect 5540 6724 5592 6730
rect 5540 6666 5592 6672
rect 5448 6384 5500 6390
rect 5448 6326 5500 6332
rect 5264 5840 5316 5846
rect 5264 5782 5316 5788
rect 5276 3398 5304 5782
rect 5264 3392 5316 3398
rect 5264 3334 5316 3340
rect 5356 3392 5408 3398
rect 5356 3334 5408 3340
rect 5276 3097 5304 3334
rect 5368 3194 5396 3334
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 5262 3088 5318 3097
rect 5262 3023 5318 3032
rect 5460 2553 5488 6326
rect 5552 5914 5580 6666
rect 5736 6390 5764 8502
rect 5816 7268 5868 7274
rect 5816 7210 5868 7216
rect 5828 6458 5856 7210
rect 6104 7206 6132 21830
rect 6380 21554 6408 23054
rect 6368 21548 6420 21554
rect 6368 21490 6420 21496
rect 6380 20806 6408 21490
rect 6368 20800 6420 20806
rect 6368 20742 6420 20748
rect 6368 18080 6420 18086
rect 6368 18022 6420 18028
rect 6380 17270 6408 18022
rect 6368 17264 6420 17270
rect 6274 17232 6330 17241
rect 6368 17206 6420 17212
rect 6274 17167 6276 17176
rect 6328 17167 6330 17176
rect 6276 17138 6328 17144
rect 6380 16590 6408 17206
rect 6368 16584 6420 16590
rect 6368 16526 6420 16532
rect 6276 16516 6328 16522
rect 6276 16458 6328 16464
rect 6288 15366 6316 16458
rect 6472 15994 6500 23598
rect 6840 21894 6868 23734
rect 6920 23724 6972 23730
rect 6920 23666 6972 23672
rect 6932 23322 6960 23666
rect 7024 23594 7052 24074
rect 7208 24070 7236 27814
rect 7472 27464 7524 27470
rect 7576 27446 7604 27950
rect 7668 27470 7696 28018
rect 7748 27532 7800 27538
rect 7748 27474 7800 27480
rect 7656 27464 7708 27470
rect 7472 27406 7524 27412
rect 7564 27440 7616 27446
rect 7484 27130 7512 27406
rect 7656 27406 7708 27412
rect 7564 27382 7616 27388
rect 7472 27124 7524 27130
rect 7472 27066 7524 27072
rect 7472 26784 7524 26790
rect 7472 26726 7524 26732
rect 7484 26450 7512 26726
rect 7472 26444 7524 26450
rect 7472 26386 7524 26392
rect 7288 26376 7340 26382
rect 7288 26318 7340 26324
rect 7196 24064 7248 24070
rect 7196 24006 7248 24012
rect 7300 23730 7328 26318
rect 7472 26240 7524 26246
rect 7472 26182 7524 26188
rect 7380 24336 7432 24342
rect 7380 24278 7432 24284
rect 7392 23730 7420 24278
rect 7484 24206 7512 26182
rect 7760 25294 7788 27474
rect 9232 27402 9260 29514
rect 9324 29102 9352 30194
rect 9404 29776 9456 29782
rect 9404 29718 9456 29724
rect 9312 29096 9364 29102
rect 9312 29038 9364 29044
rect 9220 27396 9272 27402
rect 9220 27338 9272 27344
rect 7932 27328 7984 27334
rect 7932 27270 7984 27276
rect 7944 27062 7972 27270
rect 7932 27056 7984 27062
rect 7932 26998 7984 27004
rect 9232 26926 9260 27338
rect 9220 26920 9272 26926
rect 9220 26862 9272 26868
rect 8208 26784 8260 26790
rect 8260 26732 8340 26738
rect 8208 26726 8340 26732
rect 8220 26710 8340 26726
rect 7932 26376 7984 26382
rect 7932 26318 7984 26324
rect 7944 25498 7972 26318
rect 8312 25906 8340 26710
rect 9232 26450 9260 26862
rect 9220 26444 9272 26450
rect 9220 26386 9272 26392
rect 8852 26376 8904 26382
rect 8852 26318 8904 26324
rect 8392 26308 8444 26314
rect 8392 26250 8444 26256
rect 8404 25974 8432 26250
rect 8484 26240 8536 26246
rect 8484 26182 8536 26188
rect 8392 25968 8444 25974
rect 8392 25910 8444 25916
rect 8300 25900 8352 25906
rect 8300 25842 8352 25848
rect 7932 25492 7984 25498
rect 7932 25434 7984 25440
rect 8312 25362 8340 25842
rect 8300 25356 8352 25362
rect 8300 25298 8352 25304
rect 7564 25288 7616 25294
rect 7564 25230 7616 25236
rect 7748 25288 7800 25294
rect 7748 25230 7800 25236
rect 7912 25288 7964 25294
rect 8011 25285 8063 25291
rect 7964 25236 7972 25276
rect 7912 25230 7972 25236
rect 7576 24954 7604 25230
rect 7564 24948 7616 24954
rect 7564 24890 7616 24896
rect 7472 24200 7524 24206
rect 7472 24142 7524 24148
rect 7288 23724 7340 23730
rect 7288 23666 7340 23672
rect 7380 23724 7432 23730
rect 7380 23666 7432 23672
rect 7012 23588 7064 23594
rect 7012 23530 7064 23536
rect 6920 23316 6972 23322
rect 6920 23258 6972 23264
rect 6932 22710 6960 23258
rect 7288 23112 7340 23118
rect 7288 23054 7340 23060
rect 6920 22704 6972 22710
rect 6920 22646 6972 22652
rect 6920 22432 6972 22438
rect 6920 22374 6972 22380
rect 6552 21888 6604 21894
rect 6552 21830 6604 21836
rect 6828 21888 6880 21894
rect 6828 21830 6880 21836
rect 6564 21554 6592 21830
rect 6552 21548 6604 21554
rect 6552 21490 6604 21496
rect 6644 21480 6696 21486
rect 6644 21422 6696 21428
rect 6656 21010 6684 21422
rect 6644 21004 6696 21010
rect 6644 20946 6696 20952
rect 6932 20874 6960 22374
rect 7300 22234 7328 23054
rect 7380 22500 7432 22506
rect 7380 22442 7432 22448
rect 7472 22500 7524 22506
rect 7472 22442 7524 22448
rect 7288 22228 7340 22234
rect 7288 22170 7340 22176
rect 7104 22092 7156 22098
rect 7104 22034 7156 22040
rect 6920 20868 6972 20874
rect 6920 20810 6972 20816
rect 6736 20596 6788 20602
rect 6736 20538 6788 20544
rect 6748 19718 6776 20538
rect 6736 19712 6788 19718
rect 6736 19654 6788 19660
rect 6644 17536 6696 17542
rect 6644 17478 6696 17484
rect 6656 17270 6684 17478
rect 6644 17264 6696 17270
rect 6644 17206 6696 17212
rect 6656 16658 6684 17206
rect 6644 16652 6696 16658
rect 6644 16594 6696 16600
rect 6552 16584 6604 16590
rect 6748 16538 6776 19654
rect 7116 19378 7144 22034
rect 7300 21690 7328 22170
rect 7288 21684 7340 21690
rect 7288 21626 7340 21632
rect 7288 20256 7340 20262
rect 7288 20198 7340 20204
rect 7300 19786 7328 20198
rect 7288 19780 7340 19786
rect 7288 19722 7340 19728
rect 7104 19372 7156 19378
rect 7104 19314 7156 19320
rect 7012 19304 7064 19310
rect 7012 19246 7064 19252
rect 7024 18970 7052 19246
rect 7012 18964 7064 18970
rect 7012 18906 7064 18912
rect 7116 18834 7144 19314
rect 7104 18828 7156 18834
rect 7104 18770 7156 18776
rect 6920 18284 6972 18290
rect 6920 18226 6972 18232
rect 6932 17338 6960 18226
rect 7116 17746 7144 18770
rect 7104 17740 7156 17746
rect 7104 17682 7156 17688
rect 7104 17604 7156 17610
rect 7104 17546 7156 17552
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 7116 17202 7144 17546
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 7104 17196 7156 17202
rect 7104 17138 7156 17144
rect 6552 16526 6604 16532
rect 6564 16114 6592 16526
rect 6656 16510 6776 16538
rect 6932 16522 6960 17138
rect 7010 16552 7066 16561
rect 6920 16516 6972 16522
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 6380 15978 6500 15994
rect 6368 15972 6500 15978
rect 6420 15966 6500 15972
rect 6368 15914 6420 15920
rect 6380 15570 6408 15914
rect 6460 15904 6512 15910
rect 6460 15846 6512 15852
rect 6368 15564 6420 15570
rect 6368 15506 6420 15512
rect 6276 15360 6328 15366
rect 6276 15302 6328 15308
rect 6472 14482 6500 15846
rect 6564 15026 6592 16050
rect 6552 15020 6604 15026
rect 6552 14962 6604 14968
rect 6460 14476 6512 14482
rect 6460 14418 6512 14424
rect 6656 14362 6684 16510
rect 7010 16487 7066 16496
rect 6920 16458 6972 16464
rect 6828 16244 6880 16250
rect 6828 16186 6880 16192
rect 6840 15094 6868 16186
rect 6932 15706 6960 16458
rect 7024 16454 7052 16487
rect 7012 16448 7064 16454
rect 7012 16390 7064 16396
rect 7012 16040 7064 16046
rect 7012 15982 7064 15988
rect 6920 15700 6972 15706
rect 6920 15642 6972 15648
rect 7024 15638 7052 15982
rect 7012 15632 7064 15638
rect 7012 15574 7064 15580
rect 6920 15360 6972 15366
rect 6920 15302 6972 15308
rect 6828 15088 6880 15094
rect 6472 14334 6684 14362
rect 6748 15048 6828 15076
rect 6368 12232 6420 12238
rect 6368 12174 6420 12180
rect 6184 12096 6236 12102
rect 6184 12038 6236 12044
rect 6196 11082 6224 12038
rect 6380 11694 6408 12174
rect 6472 12102 6500 14334
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 6564 12986 6592 13262
rect 6552 12980 6604 12986
rect 6552 12922 6604 12928
rect 6656 12850 6684 14010
rect 6644 12844 6696 12850
rect 6644 12786 6696 12792
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 6460 12096 6512 12102
rect 6460 12038 6512 12044
rect 6656 11898 6684 12174
rect 6644 11892 6696 11898
rect 6644 11834 6696 11840
rect 6748 11762 6776 15048
rect 6828 15030 6880 15036
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6840 14414 6868 14894
rect 6828 14408 6880 14414
rect 6828 14350 6880 14356
rect 6828 13932 6880 13938
rect 6932 13920 6960 15302
rect 7012 14272 7064 14278
rect 7116 14260 7144 17138
rect 7300 16674 7328 19722
rect 7392 17746 7420 22442
rect 7484 20602 7512 22442
rect 7576 20874 7604 24890
rect 7760 24818 7788 25230
rect 7944 25158 7972 25230
rect 8208 25288 8260 25294
rect 8063 25233 8064 25276
rect 8011 25227 8064 25233
rect 8208 25230 8260 25236
rect 7932 25152 7984 25158
rect 7932 25094 7984 25100
rect 7748 24812 7800 24818
rect 7748 24754 7800 24760
rect 7760 24206 7788 24754
rect 8036 24750 8064 25227
rect 8220 24954 8248 25230
rect 8208 24948 8260 24954
rect 8208 24890 8260 24896
rect 8024 24744 8076 24750
rect 8024 24686 8076 24692
rect 8116 24404 8168 24410
rect 8116 24346 8168 24352
rect 8128 24206 8156 24346
rect 7748 24200 7800 24206
rect 7748 24142 7800 24148
rect 8116 24200 8168 24206
rect 8116 24142 8168 24148
rect 7656 24064 7708 24070
rect 7656 24006 7708 24012
rect 7564 20868 7616 20874
rect 7564 20810 7616 20816
rect 7472 20596 7524 20602
rect 7472 20538 7524 20544
rect 7564 19780 7616 19786
rect 7564 19722 7616 19728
rect 7472 19304 7524 19310
rect 7472 19246 7524 19252
rect 7380 17740 7432 17746
rect 7380 17682 7432 17688
rect 7380 17196 7432 17202
rect 7380 17138 7432 17144
rect 7392 16794 7420 17138
rect 7380 16788 7432 16794
rect 7380 16730 7432 16736
rect 7300 16646 7420 16674
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 7208 14958 7236 15846
rect 7288 15496 7340 15502
rect 7288 15438 7340 15444
rect 7196 14952 7248 14958
rect 7196 14894 7248 14900
rect 7196 14340 7248 14346
rect 7196 14282 7248 14288
rect 7064 14232 7144 14260
rect 7012 14214 7064 14220
rect 6880 13892 6960 13920
rect 6828 13874 6880 13880
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 6368 11688 6420 11694
rect 6368 11630 6420 11636
rect 6184 11076 6236 11082
rect 6184 11018 6236 11024
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 6380 8974 6408 10406
rect 6368 8968 6420 8974
rect 6368 8910 6420 8916
rect 6748 8634 6776 11698
rect 7024 11082 7052 14214
rect 7102 13424 7158 13433
rect 7102 13359 7104 13368
rect 7156 13359 7158 13368
rect 7104 13330 7156 13336
rect 7208 12238 7236 14282
rect 7300 14074 7328 15438
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 7012 11076 7064 11082
rect 7012 11018 7064 11024
rect 7024 10674 7052 11018
rect 6828 10668 6880 10674
rect 6828 10610 6880 10616
rect 7012 10668 7064 10674
rect 7012 10610 7064 10616
rect 6840 10266 6868 10610
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 7024 10062 7052 10610
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 6920 9988 6972 9994
rect 6920 9930 6972 9936
rect 6932 9178 6960 9930
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 7116 9382 7144 9862
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6368 7404 6420 7410
rect 6368 7346 6420 7352
rect 6092 7200 6144 7206
rect 6092 7142 6144 7148
rect 6380 7002 6408 7346
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6368 6996 6420 7002
rect 6368 6938 6420 6944
rect 5908 6860 5960 6866
rect 5908 6802 5960 6808
rect 5920 6458 5948 6802
rect 6472 6662 6500 7142
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 6460 6656 6512 6662
rect 6460 6598 6512 6604
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 5724 6384 5776 6390
rect 5724 6326 5776 6332
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5920 5794 5948 6394
rect 6460 6384 6512 6390
rect 6460 6326 6512 6332
rect 5828 5766 5948 5794
rect 5828 5710 5856 5766
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 6472 5574 6500 6326
rect 6656 6254 6684 6734
rect 6644 6248 6696 6254
rect 6644 6190 6696 6196
rect 6368 5568 6420 5574
rect 6368 5510 6420 5516
rect 6460 5568 6512 5574
rect 6460 5510 6512 5516
rect 5540 5160 5592 5166
rect 5592 5108 5672 5114
rect 5540 5102 5672 5108
rect 5552 5086 5672 5102
rect 5644 4146 5672 5086
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5644 2825 5672 4082
rect 6380 3534 6408 5510
rect 6656 4758 6684 6190
rect 6748 5914 6776 8570
rect 6828 8016 6880 8022
rect 6828 7958 6880 7964
rect 6840 6866 6868 7958
rect 7196 7744 7248 7750
rect 7196 7686 7248 7692
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 6932 6730 6960 7278
rect 7208 7274 7236 7686
rect 7196 7268 7248 7274
rect 7196 7210 7248 7216
rect 6920 6724 6972 6730
rect 6920 6666 6972 6672
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6840 6254 6868 6598
rect 6932 6322 6960 6666
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 6734 5808 6790 5817
rect 6734 5743 6790 5752
rect 6748 5574 6776 5743
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6828 5296 6880 5302
rect 6828 5238 6880 5244
rect 6644 4752 6696 4758
rect 6644 4694 6696 4700
rect 6736 4072 6788 4078
rect 6736 4014 6788 4020
rect 6748 3913 6776 4014
rect 6734 3904 6790 3913
rect 6734 3839 6790 3848
rect 6368 3528 6420 3534
rect 6368 3470 6420 3476
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6460 3392 6512 3398
rect 6460 3334 6512 3340
rect 6472 3058 6500 3334
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 6564 2961 6592 3470
rect 6550 2952 6606 2961
rect 6550 2887 6606 2896
rect 6368 2848 6420 2854
rect 5630 2816 5686 2825
rect 6368 2790 6420 2796
rect 5630 2751 5686 2760
rect 5446 2544 5502 2553
rect 5172 2508 5224 2514
rect 5446 2479 5502 2488
rect 5172 2450 5224 2456
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 4344 2372 4396 2378
rect 4344 2314 4396 2320
rect 3240 2246 3292 2252
rect 3330 2272 3386 2281
rect 3252 1766 3280 2246
rect 3330 2207 3386 2216
rect 4356 1834 4384 2314
rect 4344 1828 4396 1834
rect 4344 1770 4396 1776
rect 3240 1760 3292 1766
rect 3240 1702 3292 1708
rect 2964 1692 3016 1698
rect 2964 1634 3016 1640
rect 4908 1018 4936 2382
rect 5080 2304 5132 2310
rect 5080 2246 5132 2252
rect 5092 2038 5120 2246
rect 5080 2032 5132 2038
rect 5080 1974 5132 1980
rect 5184 1290 5212 2450
rect 6380 2446 6408 2790
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 6736 2304 6788 2310
rect 6736 2246 6788 2252
rect 6748 2106 6776 2246
rect 6840 2145 6868 5238
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 6932 4826 6960 5102
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 7024 3194 7052 6598
rect 7208 6458 7236 7210
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 7208 5642 7236 6394
rect 7196 5636 7248 5642
rect 7196 5578 7248 5584
rect 7196 5092 7248 5098
rect 7196 5034 7248 5040
rect 7208 3913 7236 5034
rect 7194 3904 7250 3913
rect 7194 3839 7250 3848
rect 7300 3534 7328 8774
rect 7392 8634 7420 16646
rect 7484 14550 7512 19246
rect 7576 17202 7604 19722
rect 7564 17196 7616 17202
rect 7564 17138 7616 17144
rect 7668 16726 7696 24006
rect 7932 23792 7984 23798
rect 7932 23734 7984 23740
rect 7944 23526 7972 23734
rect 8024 23656 8076 23662
rect 8024 23598 8076 23604
rect 7932 23520 7984 23526
rect 7932 23462 7984 23468
rect 8036 22710 8064 23598
rect 8128 22760 8156 24142
rect 8300 23724 8352 23730
rect 8300 23666 8352 23672
rect 8312 23322 8340 23666
rect 8300 23316 8352 23322
rect 8300 23258 8352 23264
rect 8128 22732 8248 22760
rect 8024 22704 8076 22710
rect 8024 22646 8076 22652
rect 8220 22642 8248 22732
rect 8116 22636 8168 22642
rect 8116 22578 8168 22584
rect 8208 22636 8260 22642
rect 8208 22578 8260 22584
rect 8128 22098 8156 22578
rect 8116 22092 8168 22098
rect 8116 22034 8168 22040
rect 8024 21684 8076 21690
rect 8024 21626 8076 21632
rect 7748 21548 7800 21554
rect 7748 21490 7800 21496
rect 7760 20602 7788 21490
rect 7840 20800 7892 20806
rect 7840 20742 7892 20748
rect 7748 20596 7800 20602
rect 7748 20538 7800 20544
rect 7852 18766 7880 20742
rect 7932 20324 7984 20330
rect 7932 20266 7984 20272
rect 7944 18766 7972 20266
rect 8036 19786 8064 21626
rect 8128 21146 8156 22034
rect 8300 21888 8352 21894
rect 8300 21830 8352 21836
rect 8116 21140 8168 21146
rect 8116 21082 8168 21088
rect 8116 20868 8168 20874
rect 8116 20810 8168 20816
rect 8024 19780 8076 19786
rect 8024 19722 8076 19728
rect 7840 18760 7892 18766
rect 7840 18702 7892 18708
rect 7932 18760 7984 18766
rect 7932 18702 7984 18708
rect 7852 17082 7880 18702
rect 7944 17610 7972 18702
rect 8036 18426 8064 19722
rect 8024 18420 8076 18426
rect 8024 18362 8076 18368
rect 8024 18284 8076 18290
rect 8024 18226 8076 18232
rect 7932 17604 7984 17610
rect 7932 17546 7984 17552
rect 8036 17202 8064 18226
rect 8128 17542 8156 20810
rect 8312 20466 8340 21830
rect 8404 20942 8432 25910
rect 8496 25226 8524 26182
rect 8864 25294 8892 26318
rect 9324 26314 9352 29038
rect 9416 28422 9444 29718
rect 9784 29170 9812 30534
rect 10980 29850 11008 30602
rect 11072 30122 11100 30670
rect 11060 30116 11112 30122
rect 11060 30058 11112 30064
rect 10968 29844 11020 29850
rect 10968 29786 11020 29792
rect 11072 29646 11100 30058
rect 11060 29640 11112 29646
rect 11060 29582 11112 29588
rect 10232 29572 10284 29578
rect 10232 29514 10284 29520
rect 10244 29306 10272 29514
rect 9956 29300 10008 29306
rect 9956 29242 10008 29248
rect 10232 29300 10284 29306
rect 10232 29242 10284 29248
rect 9496 29164 9548 29170
rect 9496 29106 9548 29112
rect 9772 29164 9824 29170
rect 9772 29106 9824 29112
rect 9404 28416 9456 28422
rect 9404 28358 9456 28364
rect 9416 26432 9444 28358
rect 9508 28082 9536 29106
rect 9496 28076 9548 28082
rect 9496 28018 9548 28024
rect 9680 28076 9732 28082
rect 9680 28018 9732 28024
rect 9508 27538 9536 28018
rect 9692 27674 9720 28018
rect 9968 28014 9996 29242
rect 10048 29164 10100 29170
rect 10048 29106 10100 29112
rect 10060 28422 10088 29106
rect 11072 28558 11100 29582
rect 12452 29578 12480 31282
rect 12636 30598 12664 31350
rect 15120 31346 15148 31690
rect 15108 31340 15160 31346
rect 15160 31300 15240 31328
rect 15108 31282 15160 31288
rect 15212 31142 15240 31300
rect 13636 31136 13688 31142
rect 13636 31078 13688 31084
rect 15108 31136 15160 31142
rect 15108 31078 15160 31084
rect 15200 31136 15252 31142
rect 15200 31078 15252 31084
rect 13176 30660 13228 30666
rect 13176 30602 13228 30608
rect 12624 30592 12676 30598
rect 12624 30534 12676 30540
rect 12440 29572 12492 29578
rect 12440 29514 12492 29520
rect 12532 29232 12584 29238
rect 12532 29174 12584 29180
rect 11060 28552 11112 28558
rect 11060 28494 11112 28500
rect 10232 28484 10284 28490
rect 10232 28426 10284 28432
rect 10048 28416 10100 28422
rect 10048 28358 10100 28364
rect 10244 28218 10272 28426
rect 10232 28212 10284 28218
rect 10232 28154 10284 28160
rect 9956 28008 10008 28014
rect 9956 27950 10008 27956
rect 9680 27668 9732 27674
rect 9680 27610 9732 27616
rect 11072 27538 11100 28494
rect 11152 28416 11204 28422
rect 11152 28358 11204 28364
rect 9496 27532 9548 27538
rect 9496 27474 9548 27480
rect 11060 27532 11112 27538
rect 11060 27474 11112 27480
rect 11164 27470 11192 28358
rect 12440 28144 12492 28150
rect 12440 28086 12492 28092
rect 11152 27464 11204 27470
rect 12452 27418 12480 28086
rect 11152 27406 11204 27412
rect 12360 27390 12480 27418
rect 12360 27062 12388 27390
rect 12544 27316 12572 29174
rect 12636 28082 12664 30534
rect 12900 30388 12952 30394
rect 12900 30330 12952 30336
rect 12912 29714 12940 30330
rect 13188 30326 13216 30602
rect 13176 30320 13228 30326
rect 13176 30262 13228 30268
rect 13648 30258 13676 31078
rect 13820 30728 13872 30734
rect 13820 30670 13872 30676
rect 13452 30252 13504 30258
rect 13452 30194 13504 30200
rect 13636 30252 13688 30258
rect 13636 30194 13688 30200
rect 13464 30122 13492 30194
rect 13452 30116 13504 30122
rect 13452 30058 13504 30064
rect 13268 29776 13320 29782
rect 13268 29718 13320 29724
rect 12900 29708 12952 29714
rect 12900 29650 12952 29656
rect 12992 29640 13044 29646
rect 12992 29582 13044 29588
rect 13084 29640 13136 29646
rect 13280 29628 13308 29718
rect 13452 29708 13504 29714
rect 13452 29650 13504 29656
rect 13360 29640 13412 29646
rect 13280 29600 13360 29628
rect 13084 29582 13136 29588
rect 13360 29582 13412 29588
rect 12808 29504 12860 29510
rect 12808 29446 12860 29452
rect 12820 29170 12848 29446
rect 13004 29306 13032 29582
rect 13096 29492 13124 29582
rect 13464 29492 13492 29650
rect 13096 29464 13492 29492
rect 12992 29300 13044 29306
rect 12992 29242 13044 29248
rect 12808 29164 12860 29170
rect 12808 29106 12860 29112
rect 13004 28558 13032 29242
rect 13832 29102 13860 30670
rect 15120 30666 15148 31078
rect 15108 30660 15160 30666
rect 15108 30602 15160 30608
rect 14096 30592 14148 30598
rect 14096 30534 14148 30540
rect 14108 30258 14136 30534
rect 14096 30252 14148 30258
rect 14096 30194 14148 30200
rect 14108 29646 14136 30194
rect 14096 29640 14148 29646
rect 14096 29582 14148 29588
rect 14740 29640 14792 29646
rect 14740 29582 14792 29588
rect 14464 29232 14516 29238
rect 14464 29174 14516 29180
rect 13820 29096 13872 29102
rect 13820 29038 13872 29044
rect 12992 28552 13044 28558
rect 12992 28494 13044 28500
rect 13360 28552 13412 28558
rect 13360 28494 13412 28500
rect 13176 28484 13228 28490
rect 13176 28426 13228 28432
rect 13268 28484 13320 28490
rect 13268 28426 13320 28432
rect 12624 28076 12676 28082
rect 12624 28018 12676 28024
rect 13188 28014 13216 28426
rect 13176 28008 13228 28014
rect 13176 27950 13228 27956
rect 13280 27402 13308 28426
rect 13372 28082 13400 28494
rect 13832 28150 13860 29038
rect 14476 28558 14504 29174
rect 14648 29164 14700 29170
rect 14648 29106 14700 29112
rect 14464 28552 14516 28558
rect 14464 28494 14516 28500
rect 13820 28144 13872 28150
rect 13820 28086 13872 28092
rect 13360 28076 13412 28082
rect 13360 28018 13412 28024
rect 13728 28076 13780 28082
rect 13728 28018 13780 28024
rect 13360 27940 13412 27946
rect 13360 27882 13412 27888
rect 13268 27396 13320 27402
rect 13268 27338 13320 27344
rect 12452 27288 12572 27316
rect 12624 27328 12676 27334
rect 12348 27056 12400 27062
rect 12348 26998 12400 27004
rect 9588 26988 9640 26994
rect 9588 26930 9640 26936
rect 9600 26897 9628 26930
rect 9586 26888 9642 26897
rect 9586 26823 9588 26832
rect 9640 26823 9642 26832
rect 9680 26852 9732 26858
rect 9588 26794 9640 26800
rect 9680 26794 9732 26800
rect 9600 26763 9628 26794
rect 9692 26586 9720 26794
rect 9680 26580 9732 26586
rect 9680 26522 9732 26528
rect 9416 26404 9628 26432
rect 9312 26308 9364 26314
rect 9312 26250 9364 26256
rect 9404 25968 9456 25974
rect 9404 25910 9456 25916
rect 9036 25900 9088 25906
rect 9036 25842 9088 25848
rect 9048 25498 9076 25842
rect 9128 25696 9180 25702
rect 9128 25638 9180 25644
rect 9036 25492 9088 25498
rect 9036 25434 9088 25440
rect 9140 25294 9168 25638
rect 8852 25288 8904 25294
rect 8852 25230 8904 25236
rect 9128 25288 9180 25294
rect 9128 25230 9180 25236
rect 8484 25220 8536 25226
rect 8484 25162 8536 25168
rect 8484 24812 8536 24818
rect 8484 24754 8536 24760
rect 8668 24812 8720 24818
rect 8668 24754 8720 24760
rect 8496 22710 8524 24754
rect 8576 24744 8628 24750
rect 8576 24686 8628 24692
rect 8588 23866 8616 24686
rect 8576 23860 8628 23866
rect 8576 23802 8628 23808
rect 8484 22704 8536 22710
rect 8484 22646 8536 22652
rect 8588 22574 8616 23802
rect 8680 23322 8708 24754
rect 8864 24410 8892 25230
rect 9416 24750 9444 25910
rect 9404 24744 9456 24750
rect 9404 24686 9456 24692
rect 8852 24404 8904 24410
rect 8852 24346 8904 24352
rect 9036 24404 9088 24410
rect 9036 24346 9088 24352
rect 8864 24256 8892 24346
rect 8864 24228 8984 24256
rect 8852 24132 8904 24138
rect 8852 24074 8904 24080
rect 8864 23866 8892 24074
rect 8852 23860 8904 23866
rect 8852 23802 8904 23808
rect 8668 23316 8720 23322
rect 8668 23258 8720 23264
rect 8956 23118 8984 24228
rect 9048 23118 9076 24346
rect 9416 24206 9444 24686
rect 9404 24200 9456 24206
rect 9404 24142 9456 24148
rect 9312 24064 9364 24070
rect 9312 24006 9364 24012
rect 9324 23186 9352 24006
rect 9416 23186 9444 24142
rect 9312 23180 9364 23186
rect 9312 23122 9364 23128
rect 9404 23180 9456 23186
rect 9404 23122 9456 23128
rect 8944 23112 8996 23118
rect 8944 23054 8996 23060
rect 9036 23112 9088 23118
rect 9036 23054 9088 23060
rect 9496 23044 9548 23050
rect 9496 22986 9548 22992
rect 9036 22976 9088 22982
rect 9036 22918 9088 22924
rect 9048 22642 9076 22918
rect 9508 22778 9536 22986
rect 9496 22772 9548 22778
rect 9496 22714 9548 22720
rect 8852 22636 8904 22642
rect 8852 22578 8904 22584
rect 9036 22636 9088 22642
rect 9036 22578 9088 22584
rect 8576 22568 8628 22574
rect 8576 22510 8628 22516
rect 8864 22030 8892 22578
rect 8852 22024 8904 22030
rect 8852 21966 8904 21972
rect 8392 20936 8444 20942
rect 8392 20878 8444 20884
rect 8864 20466 8892 21966
rect 9036 21956 9088 21962
rect 9036 21898 9088 21904
rect 9312 21956 9364 21962
rect 9312 21898 9364 21904
rect 9048 21350 9076 21898
rect 9324 21690 9352 21898
rect 9312 21684 9364 21690
rect 9312 21626 9364 21632
rect 9220 21480 9272 21486
rect 9220 21422 9272 21428
rect 9036 21344 9088 21350
rect 9036 21286 9088 21292
rect 9048 20505 9076 21286
rect 9034 20496 9090 20505
rect 8300 20460 8352 20466
rect 8300 20402 8352 20408
rect 8852 20460 8904 20466
rect 9034 20431 9090 20440
rect 8852 20402 8904 20408
rect 8760 20392 8812 20398
rect 8760 20334 8812 20340
rect 8392 20052 8444 20058
rect 8392 19994 8444 20000
rect 8300 19848 8352 19854
rect 8300 19790 8352 19796
rect 8312 18290 8340 19790
rect 8404 19310 8432 19994
rect 8484 19712 8536 19718
rect 8484 19654 8536 19660
rect 8496 19514 8524 19654
rect 8484 19508 8536 19514
rect 8484 19450 8536 19456
rect 8482 19408 8538 19417
rect 8772 19378 8800 20334
rect 9232 19854 9260 21422
rect 9600 20874 9628 26404
rect 11796 26376 11848 26382
rect 11796 26318 11848 26324
rect 10416 26240 10468 26246
rect 10416 26182 10468 26188
rect 9864 25152 9916 25158
rect 9864 25094 9916 25100
rect 9876 24954 9904 25094
rect 9864 24948 9916 24954
rect 9864 24890 9916 24896
rect 9876 23866 9904 24890
rect 10428 24818 10456 26182
rect 11808 25906 11836 26318
rect 11796 25900 11848 25906
rect 11796 25842 11848 25848
rect 10416 24812 10468 24818
rect 10416 24754 10468 24760
rect 12072 24812 12124 24818
rect 12072 24754 12124 24760
rect 10968 24608 11020 24614
rect 10968 24550 11020 24556
rect 10980 24410 11008 24550
rect 10968 24404 11020 24410
rect 10968 24346 11020 24352
rect 12084 24206 12112 24754
rect 10692 24200 10744 24206
rect 12072 24200 12124 24206
rect 10744 24160 10824 24188
rect 10692 24142 10744 24148
rect 9864 23860 9916 23866
rect 9864 23802 9916 23808
rect 10140 21888 10192 21894
rect 10140 21830 10192 21836
rect 9680 21548 9732 21554
rect 9680 21490 9732 21496
rect 9692 21146 9720 21490
rect 9680 21140 9732 21146
rect 9680 21082 9732 21088
rect 10152 21010 10180 21830
rect 10600 21072 10652 21078
rect 10600 21014 10652 21020
rect 10140 21004 10192 21010
rect 10140 20946 10192 20952
rect 10324 20936 10376 20942
rect 10324 20878 10376 20884
rect 9588 20868 9640 20874
rect 9588 20810 9640 20816
rect 10336 20466 10364 20878
rect 10612 20466 10640 21014
rect 10324 20460 10376 20466
rect 10324 20402 10376 20408
rect 10600 20460 10652 20466
rect 10600 20402 10652 20408
rect 9220 19848 9272 19854
rect 9220 19790 9272 19796
rect 9128 19780 9180 19786
rect 9128 19722 9180 19728
rect 9140 19514 9168 19722
rect 9128 19508 9180 19514
rect 9128 19450 9180 19456
rect 10336 19446 10364 20402
rect 9220 19440 9272 19446
rect 9218 19408 9220 19417
rect 10324 19440 10376 19446
rect 9272 19408 9274 19417
rect 8482 19343 8484 19352
rect 8536 19343 8538 19352
rect 8760 19372 8812 19378
rect 8484 19314 8536 19320
rect 10324 19382 10376 19388
rect 9218 19343 9274 19352
rect 8760 19314 8812 19320
rect 8392 19304 8444 19310
rect 8392 19246 8444 19252
rect 8772 18766 8800 19314
rect 9036 19236 9088 19242
rect 9036 19178 9088 19184
rect 8760 18760 8812 18766
rect 8760 18702 8812 18708
rect 8852 18692 8904 18698
rect 8852 18634 8904 18640
rect 8864 18358 8892 18634
rect 9048 18630 9076 19178
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 9036 18624 9088 18630
rect 9036 18566 9088 18572
rect 8852 18352 8904 18358
rect 8852 18294 8904 18300
rect 9692 18290 9720 18770
rect 10508 18624 10560 18630
rect 10508 18566 10560 18572
rect 8300 18284 8352 18290
rect 8300 18226 8352 18232
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 9496 18080 9548 18086
rect 9496 18022 9548 18028
rect 8208 17740 8260 17746
rect 8208 17682 8260 17688
rect 8116 17536 8168 17542
rect 8116 17478 8168 17484
rect 8024 17196 8076 17202
rect 8024 17138 8076 17144
rect 7760 17054 7880 17082
rect 7656 16720 7708 16726
rect 7656 16662 7708 16668
rect 7564 16516 7616 16522
rect 7564 16458 7616 16464
rect 7576 16114 7604 16458
rect 7564 16108 7616 16114
rect 7564 16050 7616 16056
rect 7564 15972 7616 15978
rect 7564 15914 7616 15920
rect 7472 14544 7524 14550
rect 7472 14486 7524 14492
rect 7484 14414 7512 14486
rect 7472 14408 7524 14414
rect 7472 14350 7524 14356
rect 7484 12782 7512 14350
rect 7472 12776 7524 12782
rect 7472 12718 7524 12724
rect 7576 12209 7604 15914
rect 7668 14414 7696 16662
rect 7760 16046 7788 17054
rect 7840 16992 7892 16998
rect 7840 16934 7892 16940
rect 7748 16040 7800 16046
rect 7748 15982 7800 15988
rect 7760 15434 7788 15982
rect 7852 15502 7880 16934
rect 8128 16658 8156 17478
rect 8116 16652 8168 16658
rect 8116 16594 8168 16600
rect 8024 15564 8076 15570
rect 8024 15506 8076 15512
rect 7840 15496 7892 15502
rect 7840 15438 7892 15444
rect 7748 15428 7800 15434
rect 7748 15370 7800 15376
rect 7748 15020 7800 15026
rect 7748 14962 7800 14968
rect 7656 14408 7708 14414
rect 7656 14350 7708 14356
rect 7760 13938 7788 14962
rect 7852 14482 7880 15438
rect 7840 14476 7892 14482
rect 7840 14418 7892 14424
rect 8036 14278 8064 15506
rect 8220 14890 8248 17682
rect 9508 17678 9536 18022
rect 9692 17678 9720 18226
rect 9404 17672 9456 17678
rect 9404 17614 9456 17620
rect 9496 17672 9548 17678
rect 9496 17614 9548 17620
rect 9680 17672 9732 17678
rect 9680 17614 9732 17620
rect 8300 17604 8352 17610
rect 8300 17546 8352 17552
rect 8208 14884 8260 14890
rect 8208 14826 8260 14832
rect 8220 14414 8248 14826
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 8024 14272 8076 14278
rect 8024 14214 8076 14220
rect 8116 14272 8168 14278
rect 8116 14214 8168 14220
rect 7748 13932 7800 13938
rect 7748 13874 7800 13880
rect 7840 13728 7892 13734
rect 7840 13670 7892 13676
rect 7852 13394 7880 13670
rect 7840 13388 7892 13394
rect 7840 13330 7892 13336
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 7760 12374 7788 12718
rect 7852 12434 7880 13330
rect 8036 12850 8064 14214
rect 8128 14074 8156 14214
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 8220 13530 8248 14350
rect 8312 13802 8340 17546
rect 9416 16658 9444 17614
rect 10520 17202 10548 18566
rect 10600 18216 10652 18222
rect 10600 18158 10652 18164
rect 10508 17196 10560 17202
rect 10508 17138 10560 17144
rect 9864 16992 9916 16998
rect 9864 16934 9916 16940
rect 10416 16992 10468 16998
rect 10416 16934 10468 16940
rect 8760 16652 8812 16658
rect 8760 16594 8812 16600
rect 9404 16652 9456 16658
rect 9404 16594 9456 16600
rect 8392 14272 8444 14278
rect 8392 14214 8444 14220
rect 8404 14006 8432 14214
rect 8392 14000 8444 14006
rect 8392 13942 8444 13948
rect 8300 13796 8352 13802
rect 8300 13738 8352 13744
rect 8208 13524 8260 13530
rect 8208 13466 8260 13472
rect 8576 13252 8628 13258
rect 8576 13194 8628 13200
rect 8668 13252 8720 13258
rect 8668 13194 8720 13200
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 8024 12844 8076 12850
rect 8024 12786 8076 12792
rect 8208 12844 8260 12850
rect 8208 12786 8260 12792
rect 8220 12442 8248 12786
rect 8208 12436 8260 12442
rect 7852 12406 7972 12434
rect 7748 12368 7800 12374
rect 7800 12328 7880 12356
rect 7748 12310 7800 12316
rect 7760 12245 7788 12310
rect 7562 12200 7618 12209
rect 7562 12135 7618 12144
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7576 11150 7604 11494
rect 7564 11144 7616 11150
rect 7564 11086 7616 11092
rect 7748 11144 7800 11150
rect 7852 11132 7880 12328
rect 7944 12238 7972 12406
rect 8208 12378 8260 12384
rect 8312 12306 8340 13126
rect 8588 12986 8616 13194
rect 8576 12980 8628 12986
rect 8576 12922 8628 12928
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 7932 12232 7984 12238
rect 7932 12174 7984 12180
rect 7944 11354 7972 12174
rect 7932 11348 7984 11354
rect 7932 11290 7984 11296
rect 8404 11218 8432 12718
rect 8392 11212 8444 11218
rect 8392 11154 8444 11160
rect 7932 11144 7984 11150
rect 7852 11104 7932 11132
rect 7748 11086 7800 11092
rect 7932 11086 7984 11092
rect 7576 9586 7604 11086
rect 7760 10810 7788 11086
rect 7748 10804 7800 10810
rect 7748 10746 7800 10752
rect 7944 10606 7972 11086
rect 7932 10600 7984 10606
rect 7932 10542 7984 10548
rect 7944 10130 7972 10542
rect 7932 10124 7984 10130
rect 7932 10066 7984 10072
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7840 10056 7892 10062
rect 7840 9998 7892 10004
rect 7668 9722 7696 9998
rect 7852 9926 7880 9998
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 8300 9920 8352 9926
rect 8300 9862 8352 9868
rect 7656 9716 7708 9722
rect 7656 9658 7708 9664
rect 8312 9654 8340 9862
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 8116 9104 8168 9110
rect 8116 9046 8168 9052
rect 7380 8628 7432 8634
rect 7380 8570 7432 8576
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7668 7818 7696 8434
rect 7840 8424 7892 8430
rect 7838 8392 7840 8401
rect 7892 8392 7894 8401
rect 7748 8356 7800 8362
rect 7838 8327 7894 8336
rect 7748 8298 7800 8304
rect 7760 8090 7788 8298
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7656 7812 7708 7818
rect 7656 7754 7708 7760
rect 7668 7342 7696 7754
rect 7656 7336 7708 7342
rect 7656 7278 7708 7284
rect 7668 6798 7696 7278
rect 8128 6866 8156 9046
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 8220 7886 8248 8434
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8220 7732 8248 7822
rect 8392 7744 8444 7750
rect 8220 7704 8392 7732
rect 8392 7686 8444 7692
rect 8300 7472 8352 7478
rect 8300 7414 8352 7420
rect 8116 6860 8168 6866
rect 8116 6802 8168 6808
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 7932 6792 7984 6798
rect 7932 6734 7984 6740
rect 7656 6248 7708 6254
rect 7656 6190 7708 6196
rect 7564 5568 7616 5574
rect 7564 5510 7616 5516
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 7484 4729 7512 5102
rect 7470 4720 7526 4729
rect 7470 4655 7472 4664
rect 7524 4655 7526 4664
rect 7472 4626 7524 4632
rect 7484 3738 7512 4626
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 7104 3392 7156 3398
rect 7104 3334 7156 3340
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 7116 3058 7144 3334
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 7208 2378 7236 3334
rect 7300 3233 7328 3470
rect 7576 3466 7604 5510
rect 7668 5234 7696 6190
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 7760 3738 7788 5646
rect 7852 5114 7880 5646
rect 7944 5574 7972 6734
rect 8312 6390 8340 7414
rect 8404 7410 8432 7686
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8300 6384 8352 6390
rect 8300 6326 8352 6332
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 7932 5568 7984 5574
rect 7932 5510 7984 5516
rect 7944 5234 7972 5510
rect 7932 5228 7984 5234
rect 7932 5170 7984 5176
rect 7852 5086 7972 5114
rect 7840 5024 7892 5030
rect 7840 4966 7892 4972
rect 7852 4554 7880 4966
rect 7840 4548 7892 4554
rect 7840 4490 7892 4496
rect 7852 4078 7880 4490
rect 7840 4072 7892 4078
rect 7840 4014 7892 4020
rect 7944 3913 7972 5086
rect 8036 4146 8064 6258
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 8128 5370 8156 6054
rect 8208 5772 8260 5778
rect 8208 5714 8260 5720
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 8220 4622 8248 5714
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 8220 4214 8248 4558
rect 8392 4480 8444 4486
rect 8390 4448 8392 4457
rect 8444 4448 8446 4457
rect 8390 4383 8446 4392
rect 8208 4208 8260 4214
rect 8208 4150 8260 4156
rect 8024 4140 8076 4146
rect 8024 4082 8076 4088
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 7930 3904 7986 3913
rect 7930 3839 7986 3848
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 7932 3664 7984 3670
rect 7930 3632 7932 3641
rect 7984 3632 7986 3641
rect 7930 3567 7986 3576
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 7564 3460 7616 3466
rect 7564 3402 7616 3408
rect 7286 3224 7342 3233
rect 7286 3159 7342 3168
rect 7944 3074 7972 3470
rect 8036 3194 8064 4082
rect 8208 4004 8260 4010
rect 8208 3946 8260 3952
rect 8220 3602 8248 3946
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 8128 3074 8156 3130
rect 7944 3046 8156 3074
rect 7654 2680 7710 2689
rect 8312 2650 8340 4082
rect 8392 3664 8444 3670
rect 8390 3632 8392 3641
rect 8444 3632 8446 3641
rect 8390 3567 8446 3576
rect 7654 2615 7710 2624
rect 8300 2644 8352 2650
rect 7668 2446 7696 2615
rect 8300 2586 8352 2592
rect 8496 2514 8524 8774
rect 8680 8430 8708 13194
rect 8772 11150 8800 16594
rect 9876 16522 9904 16934
rect 10428 16590 10456 16934
rect 10612 16674 10640 18158
rect 10796 16794 10824 24160
rect 12072 24142 12124 24148
rect 12452 23202 12480 27288
rect 12624 27270 12676 27276
rect 12636 27062 12664 27270
rect 13372 27062 13400 27882
rect 13452 27872 13504 27878
rect 13452 27814 13504 27820
rect 13464 27674 13492 27814
rect 13452 27668 13504 27674
rect 13452 27610 13504 27616
rect 12624 27056 12676 27062
rect 12624 26998 12676 27004
rect 13360 27056 13412 27062
rect 13360 26998 13412 27004
rect 12992 26988 13044 26994
rect 12992 26930 13044 26936
rect 13004 26314 13032 26930
rect 12900 26308 12952 26314
rect 12900 26250 12952 26256
rect 12992 26308 13044 26314
rect 12992 26250 13044 26256
rect 12912 25498 12940 26250
rect 13176 25696 13228 25702
rect 13176 25638 13228 25644
rect 12900 25492 12952 25498
rect 12900 25434 12952 25440
rect 13188 25294 13216 25638
rect 13176 25288 13228 25294
rect 12990 25256 13046 25265
rect 13176 25230 13228 25236
rect 13360 25288 13412 25294
rect 13360 25230 13412 25236
rect 12990 25191 12992 25200
rect 13044 25191 13046 25200
rect 12992 25162 13044 25168
rect 12624 24948 12676 24954
rect 12624 24890 12676 24896
rect 12636 24274 12664 24890
rect 13188 24886 13216 25230
rect 13176 24880 13228 24886
rect 13176 24822 13228 24828
rect 13372 24410 13400 25230
rect 13360 24404 13412 24410
rect 13360 24346 13412 24352
rect 12624 24268 12676 24274
rect 12624 24210 12676 24216
rect 12532 24064 12584 24070
rect 12532 24006 12584 24012
rect 13360 24064 13412 24070
rect 13360 24006 13412 24012
rect 12544 23730 12572 24006
rect 12900 23860 12952 23866
rect 12900 23802 12952 23808
rect 12532 23724 12584 23730
rect 12532 23666 12584 23672
rect 12360 23174 12480 23202
rect 11058 22128 11114 22137
rect 11058 22063 11114 22072
rect 11152 22092 11204 22098
rect 10968 21956 11020 21962
rect 10968 21898 11020 21904
rect 10980 21457 11008 21898
rect 10966 21448 11022 21457
rect 10966 21383 10968 21392
rect 11020 21383 11022 21392
rect 10968 21354 11020 21360
rect 11072 20466 11100 22063
rect 11152 22034 11204 22040
rect 11164 21622 11192 22034
rect 11152 21616 11204 21622
rect 11152 21558 11204 21564
rect 11612 21616 11664 21622
rect 11612 21558 11664 21564
rect 11624 20466 11652 21558
rect 11796 21344 11848 21350
rect 11796 21286 11848 21292
rect 11808 20874 11836 21286
rect 12164 20936 12216 20942
rect 12164 20878 12216 20884
rect 11796 20868 11848 20874
rect 11796 20810 11848 20816
rect 12176 20806 12204 20878
rect 12164 20800 12216 20806
rect 12164 20742 12216 20748
rect 11060 20460 11112 20466
rect 11060 20402 11112 20408
rect 11612 20460 11664 20466
rect 11612 20402 11664 20408
rect 12360 19854 12388 23174
rect 12440 23112 12492 23118
rect 12440 23054 12492 23060
rect 12452 21554 12480 23054
rect 12808 21888 12860 21894
rect 12808 21830 12860 21836
rect 12440 21548 12492 21554
rect 12440 21490 12492 21496
rect 12716 21548 12768 21554
rect 12716 21490 12768 21496
rect 12452 20398 12480 21490
rect 12728 21146 12756 21490
rect 12716 21140 12768 21146
rect 12716 21082 12768 21088
rect 12440 20392 12492 20398
rect 12440 20334 12492 20340
rect 12452 20058 12480 20334
rect 12820 20262 12848 21830
rect 12808 20256 12860 20262
rect 12808 20198 12860 20204
rect 12440 20052 12492 20058
rect 12440 19994 12492 20000
rect 11336 19848 11388 19854
rect 11336 19790 11388 19796
rect 12348 19848 12400 19854
rect 12348 19790 12400 19796
rect 10968 18760 11020 18766
rect 10968 18702 11020 18708
rect 10980 17270 11008 18702
rect 11058 17640 11114 17649
rect 11058 17575 11114 17584
rect 10968 17264 11020 17270
rect 10968 17206 11020 17212
rect 10784 16788 10836 16794
rect 10784 16730 10836 16736
rect 10520 16646 10640 16674
rect 10520 16590 10548 16646
rect 10796 16590 10824 16730
rect 10416 16584 10468 16590
rect 10416 16526 10468 16532
rect 10508 16584 10560 16590
rect 10508 16526 10560 16532
rect 10784 16584 10836 16590
rect 10836 16532 11008 16538
rect 10784 16526 11008 16532
rect 9864 16516 9916 16522
rect 10796 16510 11008 16526
rect 9864 16458 9916 16464
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9036 15020 9088 15026
rect 9036 14962 9088 14968
rect 9220 15020 9272 15026
rect 9220 14962 9272 14968
rect 9048 14482 9076 14962
rect 9232 14618 9260 14962
rect 9220 14612 9272 14618
rect 9220 14554 9272 14560
rect 9036 14476 9088 14482
rect 9036 14418 9088 14424
rect 9048 13938 9076 14418
rect 9220 14408 9272 14414
rect 9220 14350 9272 14356
rect 9128 14340 9180 14346
rect 9128 14282 9180 14288
rect 9140 14074 9168 14282
rect 9128 14068 9180 14074
rect 9128 14010 9180 14016
rect 9036 13932 9088 13938
rect 9036 13874 9088 13880
rect 9036 13796 9088 13802
rect 9036 13738 9088 13744
rect 9048 12102 9076 13738
rect 9036 12096 9088 12102
rect 9036 12038 9088 12044
rect 8760 11144 8812 11150
rect 8760 11086 8812 11092
rect 8772 10674 8800 11086
rect 9048 11014 9076 12038
rect 9036 11008 9088 11014
rect 9036 10950 9088 10956
rect 8760 10668 8812 10674
rect 8760 10610 8812 10616
rect 8772 10198 8800 10610
rect 8760 10192 8812 10198
rect 8760 10134 8812 10140
rect 8760 9580 8812 9586
rect 8760 9522 8812 9528
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8680 4282 8708 8366
rect 8668 4276 8720 4282
rect 8668 4218 8720 4224
rect 8484 2508 8536 2514
rect 8484 2450 8536 2456
rect 8772 2446 8800 9522
rect 9232 7478 9260 14350
rect 9692 13394 9720 15438
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 9404 13252 9456 13258
rect 9784 13240 9812 14554
rect 9456 13212 9812 13240
rect 9404 13194 9456 13200
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9784 12714 9812 12922
rect 9772 12708 9824 12714
rect 9772 12650 9824 12656
rect 9876 12374 9904 16458
rect 10324 16176 10376 16182
rect 10324 16118 10376 16124
rect 10336 15162 10364 16118
rect 10784 15632 10836 15638
rect 10784 15574 10836 15580
rect 10140 15156 10192 15162
rect 10140 15098 10192 15104
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 9954 13832 10010 13841
rect 9954 13767 10010 13776
rect 9864 12368 9916 12374
rect 9864 12310 9916 12316
rect 9496 11688 9548 11694
rect 9496 11630 9548 11636
rect 9508 11558 9536 11630
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9680 10192 9732 10198
rect 9680 10134 9732 10140
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 9416 9382 9444 9998
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 9692 8362 9720 10134
rect 9968 9738 9996 13767
rect 10152 12850 10180 15098
rect 10232 15088 10284 15094
rect 10232 15030 10284 15036
rect 10140 12844 10192 12850
rect 10140 12786 10192 12792
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 10060 10713 10088 12038
rect 10140 11008 10192 11014
rect 10140 10950 10192 10956
rect 10046 10704 10102 10713
rect 10152 10674 10180 10950
rect 10046 10639 10102 10648
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 9968 9710 10088 9738
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 9864 9512 9916 9518
rect 9770 9480 9826 9489
rect 9864 9454 9916 9460
rect 9770 9415 9826 9424
rect 9680 8356 9732 8362
rect 9680 8298 9732 8304
rect 9496 7880 9548 7886
rect 9324 7840 9496 7868
rect 9220 7472 9272 7478
rect 9220 7414 9272 7420
rect 9220 6724 9272 6730
rect 9220 6666 9272 6672
rect 9232 6458 9260 6666
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 9128 6384 9180 6390
rect 9128 6326 9180 6332
rect 8852 5296 8904 5302
rect 8852 5238 8904 5244
rect 7656 2440 7708 2446
rect 7656 2382 7708 2388
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 7196 2372 7248 2378
rect 7196 2314 7248 2320
rect 8484 2372 8536 2378
rect 8484 2314 8536 2320
rect 8208 2304 8260 2310
rect 8496 2258 8524 2314
rect 8260 2252 8524 2258
rect 8208 2246 8524 2252
rect 8220 2230 8524 2246
rect 6826 2136 6882 2145
rect 6736 2100 6788 2106
rect 6826 2071 6882 2080
rect 6736 2042 6788 2048
rect 8864 1970 8892 5238
rect 8944 5092 8996 5098
rect 8944 5034 8996 5040
rect 8956 4622 8984 5034
rect 8944 4616 8996 4622
rect 8944 4558 8996 4564
rect 8956 3194 8984 4558
rect 9036 4548 9088 4554
rect 9036 4490 9088 4496
rect 9048 3738 9076 4490
rect 9140 4146 9168 6326
rect 9324 6322 9352 7840
rect 9496 7822 9548 7828
rect 9680 7812 9732 7818
rect 9680 7754 9732 7760
rect 9692 7410 9720 7754
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9784 6866 9812 9415
rect 9876 9110 9904 9454
rect 9968 9178 9996 9522
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 9864 9104 9916 9110
rect 9864 9046 9916 9052
rect 9864 6928 9916 6934
rect 9864 6870 9916 6876
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9508 6458 9536 6734
rect 9692 6633 9720 6734
rect 9678 6624 9734 6633
rect 9678 6559 9734 6568
rect 9496 6452 9548 6458
rect 9496 6394 9548 6400
rect 9312 6316 9364 6322
rect 9312 6258 9364 6264
rect 9220 5840 9272 5846
rect 9220 5782 9272 5788
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 9140 3534 9168 3878
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 9232 3058 9260 5782
rect 9324 5710 9352 6258
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9324 4486 9352 5646
rect 9508 5370 9536 6394
rect 9588 6248 9640 6254
rect 9588 6190 9640 6196
rect 9600 5914 9628 6190
rect 9588 5908 9640 5914
rect 9588 5850 9640 5856
rect 9876 5778 9904 6870
rect 10060 6730 10088 9710
rect 10152 9586 10180 10066
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 10048 6724 10100 6730
rect 10048 6666 10100 6672
rect 10152 6322 10180 7346
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 9956 6248 10008 6254
rect 9956 6190 10008 6196
rect 9864 5772 9916 5778
rect 9864 5714 9916 5720
rect 9968 5642 9996 6190
rect 9956 5636 10008 5642
rect 9956 5578 10008 5584
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 9496 5228 9548 5234
rect 9496 5170 9548 5176
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 9508 4622 9536 5170
rect 9784 4826 9812 5170
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9496 4616 9548 4622
rect 9496 4558 9548 4564
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 9508 4282 9536 4558
rect 9404 4276 9456 4282
rect 9404 4218 9456 4224
rect 9496 4276 9548 4282
rect 9496 4218 9548 4224
rect 9416 4162 9444 4218
rect 9770 4176 9826 4185
rect 9416 4134 9720 4162
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 9324 3738 9352 4014
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 9692 3641 9720 4134
rect 9770 4111 9772 4120
rect 9824 4111 9826 4120
rect 9772 4082 9824 4088
rect 9678 3632 9734 3641
rect 9678 3567 9734 3576
rect 9680 3392 9732 3398
rect 9784 3380 9812 4082
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9732 3352 9812 3380
rect 9680 3334 9732 3340
rect 9220 3052 9272 3058
rect 9220 2994 9272 3000
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 8852 1964 8904 1970
rect 8852 1906 8904 1912
rect 9140 1902 9168 2382
rect 9128 1896 9180 1902
rect 9128 1838 9180 1844
rect 9876 1834 9904 3674
rect 9968 3126 9996 5578
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 10060 4758 10088 5170
rect 10048 4752 10100 4758
rect 10048 4694 10100 4700
rect 10060 4622 10088 4694
rect 10048 4616 10100 4622
rect 10048 4558 10100 4564
rect 10152 4486 10180 6258
rect 10140 4480 10192 4486
rect 10140 4422 10192 4428
rect 10140 3392 10192 3398
rect 10046 3360 10102 3369
rect 10140 3334 10192 3340
rect 10046 3295 10102 3304
rect 10060 3126 10088 3295
rect 10152 3194 10180 3334
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 9956 3120 10008 3126
rect 9956 3062 10008 3068
rect 10048 3120 10100 3126
rect 10048 3062 10100 3068
rect 10048 2508 10100 2514
rect 10048 2450 10100 2456
rect 9956 2372 10008 2378
rect 9956 2314 10008 2320
rect 9968 1970 9996 2314
rect 10060 2281 10088 2450
rect 10046 2272 10102 2281
rect 10046 2207 10102 2216
rect 9956 1964 10008 1970
rect 9956 1906 10008 1912
rect 9864 1828 9916 1834
rect 9864 1770 9916 1776
rect 5172 1284 5224 1290
rect 5172 1226 5224 1232
rect 4896 1012 4948 1018
rect 4896 954 4948 960
rect 9680 944 9732 950
rect 9680 886 9732 892
rect 9692 202 9720 886
rect 10244 762 10272 15030
rect 10508 14816 10560 14822
rect 10508 14758 10560 14764
rect 10520 12918 10548 14758
rect 10796 14618 10824 15574
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 10508 12912 10560 12918
rect 10508 12854 10560 12860
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 10600 12844 10652 12850
rect 10600 12786 10652 12792
rect 10428 12170 10456 12786
rect 10612 12238 10640 12786
rect 10784 12640 10836 12646
rect 10784 12582 10836 12588
rect 10796 12345 10824 12582
rect 10782 12336 10838 12345
rect 10782 12271 10838 12280
rect 10600 12232 10652 12238
rect 10600 12174 10652 12180
rect 10416 12164 10468 12170
rect 10416 12106 10468 12112
rect 10428 11762 10456 12106
rect 10416 11756 10468 11762
rect 10416 11698 10468 11704
rect 10428 10810 10456 11698
rect 10416 10804 10468 10810
rect 10416 10746 10468 10752
rect 10428 10130 10456 10746
rect 10612 10674 10640 12174
rect 10980 12102 11008 16510
rect 11072 15094 11100 17575
rect 11348 16250 11376 19790
rect 12164 19440 12216 19446
rect 12164 19382 12216 19388
rect 11520 18692 11572 18698
rect 11520 18634 11572 18640
rect 11532 18426 11560 18634
rect 11520 18420 11572 18426
rect 11520 18362 11572 18368
rect 12176 18290 12204 19382
rect 12452 18766 12480 19994
rect 12440 18760 12492 18766
rect 12440 18702 12492 18708
rect 11796 18284 11848 18290
rect 11796 18226 11848 18232
rect 12164 18284 12216 18290
rect 12164 18226 12216 18232
rect 12256 18284 12308 18290
rect 12256 18226 12308 18232
rect 11808 17542 11836 18226
rect 12268 17882 12296 18226
rect 12452 18222 12480 18702
rect 12624 18692 12676 18698
rect 12624 18634 12676 18640
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 12256 17876 12308 17882
rect 12256 17818 12308 17824
rect 12452 17746 12480 18158
rect 12440 17740 12492 17746
rect 12440 17682 12492 17688
rect 11796 17536 11848 17542
rect 11796 17478 11848 17484
rect 12452 17270 12480 17682
rect 12636 17610 12664 18634
rect 12716 18080 12768 18086
rect 12716 18022 12768 18028
rect 12624 17604 12676 17610
rect 12624 17546 12676 17552
rect 12440 17264 12492 17270
rect 12440 17206 12492 17212
rect 11612 17196 11664 17202
rect 11612 17138 11664 17144
rect 11624 16522 11652 17138
rect 11612 16516 11664 16522
rect 11612 16458 11664 16464
rect 11336 16244 11388 16250
rect 11336 16186 11388 16192
rect 11348 15706 11376 16186
rect 12636 16114 12664 17546
rect 12728 17134 12756 18022
rect 12716 17128 12768 17134
rect 12716 17070 12768 17076
rect 12440 16108 12492 16114
rect 12440 16050 12492 16056
rect 12624 16108 12676 16114
rect 12624 16050 12676 16056
rect 12164 15904 12216 15910
rect 12164 15846 12216 15852
rect 11336 15700 11388 15706
rect 11336 15642 11388 15648
rect 11060 15088 11112 15094
rect 11060 15030 11112 15036
rect 11348 14346 11376 15642
rect 12176 15502 12204 15846
rect 12164 15496 12216 15502
rect 12162 15464 12164 15473
rect 12216 15464 12218 15473
rect 12162 15399 12218 15408
rect 12452 15094 12480 16050
rect 12728 15570 12756 17070
rect 12716 15564 12768 15570
rect 12716 15506 12768 15512
rect 12624 15360 12676 15366
rect 12624 15302 12676 15308
rect 12532 15156 12584 15162
rect 12532 15098 12584 15104
rect 12440 15088 12492 15094
rect 12440 15030 12492 15036
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 11900 14618 11928 14962
rect 12544 14958 12572 15098
rect 12636 15094 12664 15302
rect 12624 15088 12676 15094
rect 12624 15030 12676 15036
rect 12532 14952 12584 14958
rect 12532 14894 12584 14900
rect 11980 14816 12032 14822
rect 11980 14758 12032 14764
rect 11888 14612 11940 14618
rect 11888 14554 11940 14560
rect 11244 14340 11296 14346
rect 11244 14282 11296 14288
rect 11336 14340 11388 14346
rect 11336 14282 11388 14288
rect 11256 14074 11284 14282
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 11244 14068 11296 14074
rect 11244 14010 11296 14016
rect 11164 13326 11192 14010
rect 11992 13938 12020 14758
rect 12256 14340 12308 14346
rect 12256 14282 12308 14288
rect 11796 13932 11848 13938
rect 11796 13874 11848 13880
rect 11980 13932 12032 13938
rect 11980 13874 12032 13880
rect 11808 13734 11836 13874
rect 11888 13796 11940 13802
rect 11888 13738 11940 13744
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 11808 13530 11836 13670
rect 11796 13524 11848 13530
rect 11796 13466 11848 13472
rect 11900 13326 11928 13738
rect 11152 13320 11204 13326
rect 11152 13262 11204 13268
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 12070 13288 12126 13297
rect 11704 13252 11756 13258
rect 11704 13194 11756 13200
rect 11716 12918 11744 13194
rect 11704 12912 11756 12918
rect 11704 12854 11756 12860
rect 11520 12844 11572 12850
rect 11520 12786 11572 12792
rect 11532 12714 11560 12786
rect 11520 12708 11572 12714
rect 11520 12650 11572 12656
rect 11060 12640 11112 12646
rect 11060 12582 11112 12588
rect 11072 12306 11100 12582
rect 11716 12442 11744 12854
rect 11900 12850 11928 13262
rect 12070 13223 12126 13232
rect 12084 13190 12112 13223
rect 12072 13184 12124 13190
rect 12072 13126 12124 13132
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 11900 12646 11928 12786
rect 12070 12744 12126 12753
rect 12070 12679 12072 12688
rect 12124 12679 12126 12688
rect 12072 12650 12124 12656
rect 11888 12640 11940 12646
rect 11888 12582 11940 12588
rect 11704 12436 11756 12442
rect 11704 12378 11756 12384
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 10968 12096 11020 12102
rect 10968 12038 11020 12044
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 10612 10062 10640 10610
rect 10690 10568 10746 10577
rect 10690 10503 10692 10512
rect 10744 10503 10746 10512
rect 10692 10474 10744 10480
rect 10980 10266 11008 12038
rect 11716 11762 11744 12378
rect 11900 11762 11928 12582
rect 11704 11756 11756 11762
rect 11704 11698 11756 11704
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 12070 11656 12126 11665
rect 12070 11591 12072 11600
rect 12124 11591 12126 11600
rect 12072 11562 12124 11568
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 11428 10668 11480 10674
rect 11428 10610 11480 10616
rect 11440 10266 11468 10610
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 11428 10260 11480 10266
rect 11428 10202 11480 10208
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10600 10056 10652 10062
rect 10600 9998 10652 10004
rect 10416 9648 10468 9654
rect 10416 9590 10468 9596
rect 10324 8900 10376 8906
rect 10324 8842 10376 8848
rect 10336 4570 10364 8842
rect 10428 8566 10456 9590
rect 10612 9586 10640 9998
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10508 9376 10560 9382
rect 10506 9344 10508 9353
rect 10560 9344 10562 9353
rect 10506 9279 10562 9288
rect 10416 8560 10468 8566
rect 10416 8502 10468 8508
rect 10704 7546 10732 10066
rect 11532 10044 11560 10406
rect 12176 10062 12204 10746
rect 11612 10056 11664 10062
rect 10966 10024 11022 10033
rect 11532 10016 11612 10044
rect 11612 9998 11664 10004
rect 12164 10056 12216 10062
rect 12164 9998 12216 10004
rect 10966 9959 11022 9968
rect 10980 9926 11008 9959
rect 10968 9920 11020 9926
rect 10968 9862 11020 9868
rect 10968 9716 11020 9722
rect 10968 9658 11020 9664
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 10784 8356 10836 8362
rect 10784 8298 10836 8304
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 10600 6860 10652 6866
rect 10600 6802 10652 6808
rect 10508 6180 10560 6186
rect 10508 6122 10560 6128
rect 10336 4542 10456 4570
rect 10324 4480 10376 4486
rect 10324 4422 10376 4428
rect 10336 4214 10364 4422
rect 10324 4208 10376 4214
rect 10324 4150 10376 4156
rect 10428 3584 10456 4542
rect 10336 3556 10456 3584
rect 10336 1358 10364 3556
rect 10414 3496 10470 3505
rect 10414 3431 10416 3440
rect 10468 3431 10470 3440
rect 10416 3402 10468 3408
rect 10520 3346 10548 6122
rect 10612 6118 10640 6802
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10704 6458 10732 6734
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 10600 6112 10652 6118
rect 10600 6054 10652 6060
rect 10600 4820 10652 4826
rect 10600 4762 10652 4768
rect 10612 4282 10640 4762
rect 10600 4276 10652 4282
rect 10600 4218 10652 4224
rect 10692 4140 10744 4146
rect 10692 4082 10744 4088
rect 10704 4010 10732 4082
rect 10692 4004 10744 4010
rect 10692 3946 10744 3952
rect 10796 3738 10824 8298
rect 10888 6254 10916 8910
rect 10876 6248 10928 6254
rect 10876 6190 10928 6196
rect 10980 5234 11008 9658
rect 11624 9625 11652 9998
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 11610 9616 11666 9625
rect 11610 9551 11666 9560
rect 11520 9376 11572 9382
rect 11520 9318 11572 9324
rect 11152 8560 11204 8566
rect 11152 8502 11204 8508
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 11072 7410 11100 7686
rect 11060 7404 11112 7410
rect 11060 7346 11112 7352
rect 11164 6662 11192 8502
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11072 6390 11100 6598
rect 11060 6384 11112 6390
rect 11060 6326 11112 6332
rect 11256 5370 11284 8366
rect 11428 8356 11480 8362
rect 11428 8298 11480 8304
rect 11336 6112 11388 6118
rect 11336 6054 11388 6060
rect 11244 5364 11296 5370
rect 11244 5306 11296 5312
rect 11060 5296 11112 5302
rect 11060 5238 11112 5244
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 10876 5160 10928 5166
rect 10876 5102 10928 5108
rect 10888 3738 10916 5102
rect 10968 5024 11020 5030
rect 10968 4966 11020 4972
rect 10980 3942 11008 4966
rect 10968 3936 11020 3942
rect 10968 3878 11020 3884
rect 10966 3768 11022 3777
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 10876 3732 10928 3738
rect 10966 3703 11022 3712
rect 10876 3674 10928 3680
rect 10600 3460 10652 3466
rect 10600 3402 10652 3408
rect 10428 3318 10548 3346
rect 10428 2650 10456 3318
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 10508 2644 10560 2650
rect 10508 2586 10560 2592
rect 10428 2281 10456 2586
rect 10520 2446 10548 2586
rect 10508 2440 10560 2446
rect 10508 2382 10560 2388
rect 10414 2272 10470 2281
rect 10414 2207 10470 2216
rect 10612 1766 10640 3402
rect 10784 2576 10836 2582
rect 10784 2518 10836 2524
rect 10600 1760 10652 1766
rect 10600 1702 10652 1708
rect 10324 1352 10376 1358
rect 10324 1294 10376 1300
rect 10692 1352 10744 1358
rect 10692 1294 10744 1300
rect 10520 870 10640 898
rect 10520 762 10548 870
rect 10612 800 10640 870
rect 10704 800 10732 1294
rect 10796 800 10824 2518
rect 10876 944 10928 950
rect 10876 886 10928 892
rect 10888 800 10916 886
rect 10980 800 11008 3703
rect 11072 2774 11100 5238
rect 11152 4548 11204 4554
rect 11152 4490 11204 4496
rect 11164 4162 11192 4490
rect 11164 4134 11284 4162
rect 11256 4010 11284 4134
rect 11244 4004 11296 4010
rect 11244 3946 11296 3952
rect 11256 3602 11284 3946
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 11256 2990 11284 3538
rect 11244 2984 11296 2990
rect 11244 2926 11296 2932
rect 11072 2746 11192 2774
rect 11060 2576 11112 2582
rect 11060 2518 11112 2524
rect 11072 2310 11100 2518
rect 11164 2446 11192 2746
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 11060 2304 11112 2310
rect 11060 2246 11112 2252
rect 11060 1692 11112 1698
rect 11060 1634 11112 1640
rect 11072 800 11100 1634
rect 11164 800 11192 2382
rect 11244 1964 11296 1970
rect 11244 1906 11296 1912
rect 11256 800 11284 1906
rect 11348 800 11376 6054
rect 11440 800 11468 8298
rect 11532 3040 11560 9318
rect 11992 9042 12020 9862
rect 12176 9586 12204 9998
rect 12164 9580 12216 9586
rect 12164 9522 12216 9528
rect 12072 9104 12124 9110
rect 12072 9046 12124 9052
rect 11980 9036 12032 9042
rect 11980 8978 12032 8984
rect 11992 8430 12020 8978
rect 12084 8498 12112 9046
rect 12072 8492 12124 8498
rect 12072 8434 12124 8440
rect 12164 8492 12216 8498
rect 12164 8434 12216 8440
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 11888 8356 11940 8362
rect 11888 8298 11940 8304
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11612 7336 11664 7342
rect 11612 7278 11664 7284
rect 11624 6730 11652 7278
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11612 6724 11664 6730
rect 11612 6666 11664 6672
rect 11716 6118 11744 6734
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11808 5930 11836 7822
rect 11624 5902 11836 5930
rect 11624 4457 11652 5902
rect 11900 5642 11928 8298
rect 11992 7410 12020 8366
rect 12084 7478 12112 8434
rect 12176 8090 12204 8434
rect 12268 8362 12296 14282
rect 12438 12200 12494 12209
rect 12438 12135 12494 12144
rect 12452 11286 12480 12135
rect 12440 11280 12492 11286
rect 12440 11222 12492 11228
rect 12544 10742 12572 14894
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 12636 13938 12664 14214
rect 12624 13932 12676 13938
rect 12624 13874 12676 13880
rect 12636 12238 12664 13874
rect 12728 13870 12756 15506
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 12820 12714 12848 20198
rect 12912 17270 12940 23802
rect 13372 23798 13400 24006
rect 13360 23792 13412 23798
rect 13360 23734 13412 23740
rect 12992 23724 13044 23730
rect 12992 23666 13044 23672
rect 13004 23322 13032 23666
rect 13268 23520 13320 23526
rect 13268 23462 13320 23468
rect 12992 23316 13044 23322
rect 12992 23258 13044 23264
rect 13004 22642 13032 23258
rect 13280 23050 13308 23462
rect 13268 23044 13320 23050
rect 13268 22986 13320 22992
rect 12992 22636 13044 22642
rect 12992 22578 13044 22584
rect 13464 20233 13492 27610
rect 13740 26994 13768 28018
rect 13728 26988 13780 26994
rect 13728 26930 13780 26936
rect 13740 26450 13768 26930
rect 13728 26444 13780 26450
rect 13728 26386 13780 26392
rect 13740 24818 13768 26386
rect 13832 26382 13860 28086
rect 14096 27872 14148 27878
rect 14096 27814 14148 27820
rect 14108 27470 14136 27814
rect 14096 27464 14148 27470
rect 14096 27406 14148 27412
rect 14280 27056 14332 27062
rect 14280 26998 14332 27004
rect 13912 26784 13964 26790
rect 13912 26726 13964 26732
rect 13820 26376 13872 26382
rect 13820 26318 13872 26324
rect 13820 26240 13872 26246
rect 13820 26182 13872 26188
rect 13728 24812 13780 24818
rect 13728 24754 13780 24760
rect 13832 24138 13860 26182
rect 13924 25294 13952 26726
rect 14096 26580 14148 26586
rect 14096 26522 14148 26528
rect 14108 26382 14136 26522
rect 14096 26376 14148 26382
rect 14096 26318 14148 26324
rect 14108 26042 14136 26318
rect 14292 26314 14320 26998
rect 14280 26308 14332 26314
rect 14280 26250 14332 26256
rect 14372 26308 14424 26314
rect 14372 26250 14424 26256
rect 14096 26036 14148 26042
rect 14096 25978 14148 25984
rect 14096 25832 14148 25838
rect 14096 25774 14148 25780
rect 14108 25362 14136 25774
rect 14096 25356 14148 25362
rect 14096 25298 14148 25304
rect 13912 25288 13964 25294
rect 13912 25230 13964 25236
rect 14292 25242 14320 26250
rect 14384 25430 14412 26250
rect 14476 26042 14504 28494
rect 14556 27464 14608 27470
rect 14556 27406 14608 27412
rect 14568 27130 14596 27406
rect 14660 27402 14688 29106
rect 14752 27470 14780 29582
rect 15212 29306 15240 31078
rect 15304 30938 15332 31690
rect 15568 31680 15620 31686
rect 15568 31622 15620 31628
rect 18512 31680 18564 31686
rect 18512 31622 18564 31628
rect 15580 31346 15608 31622
rect 15936 31408 15988 31414
rect 15936 31350 15988 31356
rect 15568 31340 15620 31346
rect 15568 31282 15620 31288
rect 15752 31340 15804 31346
rect 15752 31282 15804 31288
rect 15660 31204 15712 31210
rect 15660 31146 15712 31152
rect 15292 30932 15344 30938
rect 15292 30874 15344 30880
rect 15304 30258 15332 30874
rect 15672 30258 15700 31146
rect 15764 30598 15792 31282
rect 15752 30592 15804 30598
rect 15752 30534 15804 30540
rect 15948 30394 15976 31350
rect 18524 31346 18552 31622
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 17408 31340 17460 31346
rect 17408 31282 17460 31288
rect 17592 31340 17644 31346
rect 17592 31282 17644 31288
rect 18512 31340 18564 31346
rect 18512 31282 18564 31288
rect 19524 31340 19576 31346
rect 19524 31282 19576 31288
rect 17420 31142 17448 31282
rect 17408 31136 17460 31142
rect 17408 31078 17460 31084
rect 17420 30802 17448 31078
rect 17408 30796 17460 30802
rect 17408 30738 17460 30744
rect 17604 30598 17632 31282
rect 18236 31136 18288 31142
rect 18236 31078 18288 31084
rect 18248 30734 18276 31078
rect 19536 30938 19564 31282
rect 20076 31272 20128 31278
rect 20076 31214 20128 31220
rect 19984 31136 20036 31142
rect 19984 31078 20036 31084
rect 19524 30932 19576 30938
rect 19524 30874 19576 30880
rect 18236 30728 18288 30734
rect 18236 30670 18288 30676
rect 19432 30660 19484 30666
rect 19432 30602 19484 30608
rect 17408 30592 17460 30598
rect 17408 30534 17460 30540
rect 17592 30592 17644 30598
rect 17592 30534 17644 30540
rect 15936 30388 15988 30394
rect 15936 30330 15988 30336
rect 15292 30252 15344 30258
rect 15292 30194 15344 30200
rect 15660 30252 15712 30258
rect 15660 30194 15712 30200
rect 15948 29306 15976 30330
rect 17132 30320 17184 30326
rect 17132 30262 17184 30268
rect 16580 30184 16632 30190
rect 16580 30126 16632 30132
rect 16592 29510 16620 30126
rect 17040 29708 17092 29714
rect 17040 29650 17092 29656
rect 16580 29504 16632 29510
rect 16580 29446 16632 29452
rect 15200 29300 15252 29306
rect 15200 29242 15252 29248
rect 15936 29300 15988 29306
rect 15936 29242 15988 29248
rect 16592 29170 16620 29446
rect 16304 29164 16356 29170
rect 16304 29106 16356 29112
rect 16580 29164 16632 29170
rect 16580 29106 16632 29112
rect 15108 28416 15160 28422
rect 15108 28358 15160 28364
rect 15120 28150 15148 28358
rect 15108 28144 15160 28150
rect 15108 28086 15160 28092
rect 15384 28076 15436 28082
rect 15384 28018 15436 28024
rect 14832 27872 14884 27878
rect 14832 27814 14884 27820
rect 15108 27872 15160 27878
rect 15108 27814 15160 27820
rect 14740 27464 14792 27470
rect 14740 27406 14792 27412
rect 14648 27396 14700 27402
rect 14648 27338 14700 27344
rect 14660 27130 14688 27338
rect 14556 27124 14608 27130
rect 14556 27066 14608 27072
rect 14648 27124 14700 27130
rect 14648 27066 14700 27072
rect 14464 26036 14516 26042
rect 14464 25978 14516 25984
rect 14660 25906 14688 27066
rect 14752 26382 14780 27406
rect 14740 26376 14792 26382
rect 14740 26318 14792 26324
rect 14740 26240 14792 26246
rect 14740 26182 14792 26188
rect 14648 25900 14700 25906
rect 14648 25842 14700 25848
rect 14752 25702 14780 26182
rect 14740 25696 14792 25702
rect 14740 25638 14792 25644
rect 14372 25424 14424 25430
rect 14372 25366 14424 25372
rect 14372 25288 14424 25294
rect 14292 25236 14372 25242
rect 14292 25230 14424 25236
rect 13820 24132 13872 24138
rect 13820 24074 13872 24080
rect 13544 23724 13596 23730
rect 13544 23666 13596 23672
rect 13556 23254 13584 23666
rect 13544 23248 13596 23254
rect 13544 23190 13596 23196
rect 13832 23202 13860 24074
rect 13924 23730 13952 25230
rect 14292 25214 14412 25230
rect 14384 24818 14412 25214
rect 14372 24812 14424 24818
rect 14372 24754 14424 24760
rect 14280 24744 14332 24750
rect 14280 24686 14332 24692
rect 14292 24206 14320 24686
rect 14740 24608 14792 24614
rect 14740 24550 14792 24556
rect 14280 24200 14332 24206
rect 14280 24142 14332 24148
rect 13912 23724 13964 23730
rect 13912 23666 13964 23672
rect 13832 23174 13952 23202
rect 14292 23186 14320 24142
rect 13820 23112 13872 23118
rect 13820 23054 13872 23060
rect 13832 22710 13860 23054
rect 13924 23050 13952 23174
rect 14280 23180 14332 23186
rect 14280 23122 14332 23128
rect 13912 23044 13964 23050
rect 13912 22986 13964 22992
rect 13820 22704 13872 22710
rect 13820 22646 13872 22652
rect 13912 22704 13964 22710
rect 13912 22646 13964 22652
rect 13924 22545 13952 22646
rect 14292 22574 14320 23122
rect 14752 23118 14780 24550
rect 14740 23112 14792 23118
rect 14740 23054 14792 23060
rect 14280 22568 14332 22574
rect 13910 22536 13966 22545
rect 14280 22510 14332 22516
rect 13910 22471 13966 22480
rect 14292 22166 14320 22510
rect 14280 22160 14332 22166
rect 14280 22102 14332 22108
rect 13450 20224 13506 20233
rect 13450 20159 13506 20168
rect 12992 19236 13044 19242
rect 12992 19178 13044 19184
rect 13004 18970 13032 19178
rect 13084 19168 13136 19174
rect 13084 19110 13136 19116
rect 12992 18964 13044 18970
rect 12992 18906 13044 18912
rect 12900 17264 12952 17270
rect 12900 17206 12952 17212
rect 13096 16522 13124 19110
rect 13176 18624 13228 18630
rect 13176 18566 13228 18572
rect 13188 18358 13216 18566
rect 13464 18442 13492 20159
rect 13464 18414 13676 18442
rect 13176 18352 13228 18358
rect 13176 18294 13228 18300
rect 13544 17536 13596 17542
rect 13544 17478 13596 17484
rect 13452 17264 13504 17270
rect 13452 17206 13504 17212
rect 13268 17196 13320 17202
rect 13268 17138 13320 17144
rect 13280 16590 13308 17138
rect 13268 16584 13320 16590
rect 13268 16526 13320 16532
rect 13084 16516 13136 16522
rect 13084 16458 13136 16464
rect 13084 15904 13136 15910
rect 13084 15846 13136 15852
rect 13096 15502 13124 15846
rect 13280 15502 13308 16526
rect 13084 15496 13136 15502
rect 13084 15438 13136 15444
rect 13268 15496 13320 15502
rect 13268 15438 13320 15444
rect 13280 14006 13308 15438
rect 13360 15428 13412 15434
rect 13360 15370 13412 15376
rect 13372 14278 13400 15370
rect 13360 14272 13412 14278
rect 13360 14214 13412 14220
rect 13268 14000 13320 14006
rect 13268 13942 13320 13948
rect 13176 13252 13228 13258
rect 13176 13194 13228 13200
rect 12808 12708 12860 12714
rect 12808 12650 12860 12656
rect 12624 12232 12676 12238
rect 12622 12200 12624 12209
rect 13084 12232 13136 12238
rect 12676 12200 12678 12209
rect 13084 12174 13136 12180
rect 12622 12135 12678 12144
rect 12900 12164 12952 12170
rect 12900 12106 12952 12112
rect 12912 11762 12940 12106
rect 12900 11756 12952 11762
rect 12900 11698 12952 11704
rect 12532 10736 12584 10742
rect 12532 10678 12584 10684
rect 12624 10192 12676 10198
rect 12624 10134 12676 10140
rect 12636 9586 12664 10134
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12532 9512 12584 9518
rect 12532 9454 12584 9460
rect 12544 9178 12572 9454
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12440 9036 12492 9042
rect 12440 8978 12492 8984
rect 12452 8634 12480 8978
rect 12544 8650 12572 9114
rect 12440 8628 12492 8634
rect 12544 8622 12664 8650
rect 12440 8570 12492 8576
rect 12532 8492 12584 8498
rect 12452 8452 12532 8480
rect 12256 8356 12308 8362
rect 12256 8298 12308 8304
rect 12164 8084 12216 8090
rect 12164 8026 12216 8032
rect 12164 7948 12216 7954
rect 12164 7890 12216 7896
rect 12072 7472 12124 7478
rect 12072 7414 12124 7420
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 11888 5636 11940 5642
rect 11888 5578 11940 5584
rect 11980 5160 12032 5166
rect 11980 5102 12032 5108
rect 11992 4826 12020 5102
rect 11980 4820 12032 4826
rect 11980 4762 12032 4768
rect 11704 4752 11756 4758
rect 11704 4694 11756 4700
rect 11796 4752 11848 4758
rect 11848 4712 11928 4740
rect 11796 4694 11848 4700
rect 11716 4604 11744 4694
rect 11716 4576 11836 4604
rect 11610 4448 11666 4457
rect 11610 4383 11666 4392
rect 11624 3194 11652 4383
rect 11704 4208 11756 4214
rect 11704 4150 11756 4156
rect 11612 3188 11664 3194
rect 11612 3130 11664 3136
rect 11612 3052 11664 3058
rect 11532 3012 11612 3040
rect 11612 2994 11664 3000
rect 11518 2816 11574 2825
rect 11518 2751 11574 2760
rect 11532 800 11560 2751
rect 11624 800 11652 2994
rect 11716 2854 11744 4150
rect 11808 4010 11836 4576
rect 11900 4214 11928 4712
rect 11992 4554 12020 4762
rect 12072 4752 12124 4758
rect 12072 4694 12124 4700
rect 11980 4548 12032 4554
rect 11980 4490 12032 4496
rect 12084 4282 12112 4694
rect 12072 4276 12124 4282
rect 12072 4218 12124 4224
rect 11888 4208 11940 4214
rect 11888 4150 11940 4156
rect 11900 4010 11928 4150
rect 12084 4078 12112 4218
rect 12072 4072 12124 4078
rect 12072 4014 12124 4020
rect 12176 4026 12204 7890
rect 12452 7750 12480 8452
rect 12532 8434 12584 8440
rect 12532 8016 12584 8022
rect 12532 7958 12584 7964
rect 12440 7744 12492 7750
rect 12440 7686 12492 7692
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12360 5574 12388 6598
rect 12452 6390 12480 7686
rect 12440 6384 12492 6390
rect 12440 6326 12492 6332
rect 12348 5568 12400 5574
rect 12348 5510 12400 5516
rect 12348 5228 12400 5234
rect 12348 5170 12400 5176
rect 12360 4214 12388 5170
rect 12544 5030 12572 7958
rect 12636 6866 12664 8622
rect 12624 6860 12676 6866
rect 12624 6802 12676 6808
rect 12636 6390 12664 6802
rect 12624 6384 12676 6390
rect 12624 6326 12676 6332
rect 12624 5568 12676 5574
rect 12624 5510 12676 5516
rect 12532 5024 12584 5030
rect 12532 4966 12584 4972
rect 12544 4758 12572 4966
rect 12532 4752 12584 4758
rect 12532 4694 12584 4700
rect 12440 4616 12492 4622
rect 12440 4558 12492 4564
rect 12348 4208 12400 4214
rect 12348 4150 12400 4156
rect 12348 4072 12400 4078
rect 11796 4004 11848 4010
rect 11796 3946 11848 3952
rect 11888 4004 11940 4010
rect 12176 3998 12296 4026
rect 12348 4014 12400 4020
rect 11888 3946 11940 3952
rect 11808 3738 11836 3946
rect 11900 3738 11928 3946
rect 12072 3936 12124 3942
rect 12072 3878 12124 3884
rect 12164 3936 12216 3942
rect 12164 3878 12216 3884
rect 11796 3732 11848 3738
rect 11796 3674 11848 3680
rect 11888 3732 11940 3738
rect 11888 3674 11940 3680
rect 11808 3466 11836 3674
rect 11796 3460 11848 3466
rect 11796 3402 11848 3408
rect 11808 3058 11836 3402
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 11980 3188 12032 3194
rect 11980 3130 12032 3136
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 11808 2922 11836 2994
rect 11900 2922 11928 3130
rect 11796 2916 11848 2922
rect 11796 2858 11848 2864
rect 11888 2916 11940 2922
rect 11888 2858 11940 2864
rect 11704 2848 11756 2854
rect 11704 2790 11756 2796
rect 11716 2514 11744 2790
rect 11992 2632 12020 3130
rect 11900 2604 12020 2632
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 11900 2378 11928 2604
rect 11888 2372 11940 2378
rect 11888 2314 11940 2320
rect 11704 2100 11756 2106
rect 11704 2042 11756 2048
rect 11716 800 11744 2042
rect 11900 1850 11928 2314
rect 11900 1822 12020 1850
rect 11888 1284 11940 1290
rect 11888 1226 11940 1232
rect 11900 800 11928 1226
rect 11992 800 12020 1822
rect 12084 800 12112 3878
rect 12176 3058 12204 3878
rect 12268 3194 12296 3998
rect 12360 3602 12388 4014
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12256 3188 12308 3194
rect 12256 3130 12308 3136
rect 12360 3058 12388 3538
rect 12452 3398 12480 4558
rect 12532 4480 12584 4486
rect 12532 4422 12584 4428
rect 12440 3392 12492 3398
rect 12440 3334 12492 3340
rect 12164 3052 12216 3058
rect 12164 2994 12216 3000
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 12452 2990 12480 3334
rect 12440 2984 12492 2990
rect 12254 2952 12310 2961
rect 12440 2926 12492 2932
rect 12254 2887 12310 2896
rect 12164 2508 12216 2514
rect 12164 2450 12216 2456
rect 12176 2038 12204 2450
rect 12164 2032 12216 2038
rect 12164 1974 12216 1980
rect 12268 800 12296 2887
rect 12440 2576 12492 2582
rect 12440 2518 12492 2524
rect 12348 2032 12400 2038
rect 12348 1974 12400 1980
rect 12360 800 12388 1974
rect 12452 800 12480 2518
rect 12544 898 12572 4422
rect 12636 1426 12664 5510
rect 12728 2378 12756 9862
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 12820 7886 12848 8230
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12808 6996 12860 7002
rect 12808 6938 12860 6944
rect 12820 4078 12848 6938
rect 12912 5098 12940 11698
rect 13096 6882 13124 12174
rect 13188 12102 13216 13194
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 13188 11694 13216 12038
rect 13372 11898 13400 14214
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 13176 11688 13228 11694
rect 13176 11630 13228 11636
rect 13188 7002 13216 11630
rect 13372 11558 13400 11834
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 13464 11354 13492 17206
rect 13556 17202 13584 17478
rect 13544 17196 13596 17202
rect 13544 17138 13596 17144
rect 13544 16516 13596 16522
rect 13544 16458 13596 16464
rect 13556 15910 13584 16458
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13556 15434 13584 15846
rect 13544 15428 13596 15434
rect 13544 15370 13596 15376
rect 13648 13870 13676 18414
rect 14004 16992 14056 16998
rect 14004 16934 14056 16940
rect 14016 16590 14044 16934
rect 14004 16584 14056 16590
rect 14004 16526 14056 16532
rect 13912 16176 13964 16182
rect 13912 16118 13964 16124
rect 13924 14890 13952 16118
rect 14188 15496 14240 15502
rect 14188 15438 14240 15444
rect 13912 14884 13964 14890
rect 13912 14826 13964 14832
rect 14096 14408 14148 14414
rect 14096 14350 14148 14356
rect 14108 13938 14136 14350
rect 14200 14074 14228 15438
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 13820 13252 13872 13258
rect 13820 13194 13872 13200
rect 13832 12850 13860 13194
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 14188 12844 14240 12850
rect 14188 12786 14240 12792
rect 14200 12646 14228 12786
rect 14188 12640 14240 12646
rect 14186 12608 14188 12617
rect 14240 12608 14242 12617
rect 14186 12543 14242 12552
rect 14292 12374 14320 22102
rect 14844 22030 14872 27814
rect 15016 27464 15068 27470
rect 15016 27406 15068 27412
rect 14924 26512 14976 26518
rect 14924 26454 14976 26460
rect 14936 26246 14964 26454
rect 15028 26314 15056 27406
rect 15120 26994 15148 27814
rect 15396 27130 15424 28018
rect 16212 27872 16264 27878
rect 16212 27814 16264 27820
rect 15936 27328 15988 27334
rect 15936 27270 15988 27276
rect 16028 27328 16080 27334
rect 16028 27270 16080 27276
rect 15384 27124 15436 27130
rect 15384 27066 15436 27072
rect 15568 27056 15620 27062
rect 15568 26998 15620 27004
rect 15108 26988 15160 26994
rect 15108 26930 15160 26936
rect 15200 26920 15252 26926
rect 15200 26862 15252 26868
rect 15212 26586 15240 26862
rect 15476 26784 15528 26790
rect 15476 26726 15528 26732
rect 15488 26586 15516 26726
rect 15200 26580 15252 26586
rect 15200 26522 15252 26528
rect 15476 26580 15528 26586
rect 15476 26522 15528 26528
rect 15120 26382 15148 26413
rect 15108 26376 15160 26382
rect 15384 26376 15436 26382
rect 15160 26324 15332 26330
rect 15108 26318 15332 26324
rect 15384 26318 15436 26324
rect 15016 26308 15068 26314
rect 15016 26250 15068 26256
rect 15120 26302 15332 26318
rect 14924 26240 14976 26246
rect 14924 26182 14976 26188
rect 14924 25832 14976 25838
rect 14924 25774 14976 25780
rect 14936 23050 14964 25774
rect 15028 25226 15056 26250
rect 15016 25220 15068 25226
rect 15016 25162 15068 25168
rect 15028 23866 15056 25162
rect 15120 24206 15148 26302
rect 15304 26246 15332 26302
rect 15200 26240 15252 26246
rect 15200 26182 15252 26188
rect 15292 26240 15344 26246
rect 15292 26182 15344 26188
rect 15212 25974 15240 26182
rect 15200 25968 15252 25974
rect 15200 25910 15252 25916
rect 15396 25158 15424 26318
rect 15580 25906 15608 26998
rect 15948 26994 15976 27270
rect 15752 26988 15804 26994
rect 15752 26930 15804 26936
rect 15936 26988 15988 26994
rect 15936 26930 15988 26936
rect 15764 26874 15792 26930
rect 16040 26874 16068 27270
rect 16120 26988 16172 26994
rect 16120 26930 16172 26936
rect 15764 26846 16068 26874
rect 15660 26784 15712 26790
rect 15660 26726 15712 26732
rect 15672 26382 15700 26726
rect 15660 26376 15712 26382
rect 15660 26318 15712 26324
rect 15568 25900 15620 25906
rect 15568 25842 15620 25848
rect 15384 25152 15436 25158
rect 15384 25094 15436 25100
rect 15476 24812 15528 24818
rect 15476 24754 15528 24760
rect 15108 24200 15160 24206
rect 15108 24142 15160 24148
rect 15488 23866 15516 24754
rect 15568 24336 15620 24342
rect 15568 24278 15620 24284
rect 15580 23866 15608 24278
rect 15016 23860 15068 23866
rect 15016 23802 15068 23808
rect 15476 23860 15528 23866
rect 15476 23802 15528 23808
rect 15568 23860 15620 23866
rect 15568 23802 15620 23808
rect 15016 23724 15068 23730
rect 15016 23666 15068 23672
rect 15660 23724 15712 23730
rect 15660 23666 15712 23672
rect 15028 23322 15056 23666
rect 15672 23322 15700 23666
rect 15764 23322 15792 26846
rect 16132 26586 16160 26930
rect 16120 26580 16172 26586
rect 16120 26522 16172 26528
rect 15936 25152 15988 25158
rect 15936 25094 15988 25100
rect 15948 24954 15976 25094
rect 15936 24948 15988 24954
rect 15936 24890 15988 24896
rect 16120 24948 16172 24954
rect 16120 24890 16172 24896
rect 16028 24880 16080 24886
rect 16028 24822 16080 24828
rect 15016 23316 15068 23322
rect 15016 23258 15068 23264
rect 15660 23316 15712 23322
rect 15660 23258 15712 23264
rect 15752 23316 15804 23322
rect 15752 23258 15804 23264
rect 15382 23080 15438 23089
rect 14924 23044 14976 23050
rect 15382 23015 15384 23024
rect 14924 22986 14976 22992
rect 15436 23015 15438 23024
rect 15384 22986 15436 22992
rect 15016 22976 15068 22982
rect 15016 22918 15068 22924
rect 15108 22976 15160 22982
rect 15108 22918 15160 22924
rect 15028 22710 15056 22918
rect 15016 22704 15068 22710
rect 15016 22646 15068 22652
rect 14924 22636 14976 22642
rect 14924 22578 14976 22584
rect 14936 22094 14964 22578
rect 14936 22066 15056 22094
rect 14832 22024 14884 22030
rect 14832 21966 14884 21972
rect 14740 21956 14792 21962
rect 14740 21898 14792 21904
rect 14372 21888 14424 21894
rect 14372 21830 14424 21836
rect 14384 21554 14412 21830
rect 14372 21548 14424 21554
rect 14372 21490 14424 21496
rect 14372 20868 14424 20874
rect 14372 20810 14424 20816
rect 14384 18902 14412 20810
rect 14464 19372 14516 19378
rect 14464 19314 14516 19320
rect 14372 18896 14424 18902
rect 14372 18838 14424 18844
rect 14384 16250 14412 18838
rect 14476 18630 14504 19314
rect 14464 18624 14516 18630
rect 14464 18566 14516 18572
rect 14372 16244 14424 16250
rect 14372 16186 14424 16192
rect 14384 15502 14412 16186
rect 14372 15496 14424 15502
rect 14372 15438 14424 15444
rect 14372 15020 14424 15026
rect 14372 14962 14424 14968
rect 14384 14346 14412 14962
rect 14476 14414 14504 18566
rect 14556 17332 14608 17338
rect 14556 17274 14608 17280
rect 14464 14408 14516 14414
rect 14464 14350 14516 14356
rect 14372 14340 14424 14346
rect 14372 14282 14424 14288
rect 14568 14226 14596 17274
rect 14476 14198 14596 14226
rect 14280 12368 14332 12374
rect 14280 12310 14332 12316
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 14186 11928 14242 11937
rect 14186 11863 14188 11872
rect 14240 11863 14242 11872
rect 14188 11834 14240 11840
rect 13728 11756 13780 11762
rect 13728 11698 13780 11704
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13268 11076 13320 11082
rect 13268 11018 13320 11024
rect 13280 10538 13308 11018
rect 13268 10532 13320 10538
rect 13268 10474 13320 10480
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 13004 6854 13124 6882
rect 12900 5092 12952 5098
rect 12900 5034 12952 5040
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 12898 4040 12954 4049
rect 12898 3975 12954 3984
rect 12912 3738 12940 3975
rect 12900 3732 12952 3738
rect 12900 3674 12952 3680
rect 12900 3528 12952 3534
rect 12900 3470 12952 3476
rect 12912 3126 12940 3470
rect 13004 3194 13032 6854
rect 13176 5704 13228 5710
rect 13176 5646 13228 5652
rect 13084 5364 13136 5370
rect 13084 5306 13136 5312
rect 12992 3188 13044 3194
rect 12992 3130 13044 3136
rect 13096 3126 13124 5306
rect 12900 3120 12952 3126
rect 12900 3062 12952 3068
rect 13084 3120 13136 3126
rect 13084 3062 13136 3068
rect 13188 2774 13216 5646
rect 13280 5302 13308 10474
rect 13464 10470 13492 11290
rect 13740 11150 13768 11698
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13820 11008 13872 11014
rect 13820 10950 13872 10956
rect 14280 11008 14332 11014
rect 14280 10950 14332 10956
rect 13452 10464 13504 10470
rect 13452 10406 13504 10412
rect 13832 9994 13860 10950
rect 14292 10674 14320 10950
rect 13912 10668 13964 10674
rect 13912 10610 13964 10616
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 13924 10441 13952 10610
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 13910 10432 13966 10441
rect 13910 10367 13966 10376
rect 14016 10266 14044 10542
rect 14004 10260 14056 10266
rect 14004 10202 14056 10208
rect 14108 10062 14136 10542
rect 14096 10056 14148 10062
rect 14096 9998 14148 10004
rect 13820 9988 13872 9994
rect 13820 9930 13872 9936
rect 13544 9920 13596 9926
rect 13544 9862 13596 9868
rect 14188 9920 14240 9926
rect 14188 9862 14240 9868
rect 13360 9512 13412 9518
rect 13360 9454 13412 9460
rect 13372 9382 13400 9454
rect 13360 9376 13412 9382
rect 13360 9318 13412 9324
rect 13372 8294 13400 9318
rect 13556 8401 13584 9862
rect 13636 9104 13688 9110
rect 13636 9046 13688 9052
rect 13648 8430 13676 9046
rect 13636 8424 13688 8430
rect 13542 8392 13598 8401
rect 13636 8366 13688 8372
rect 13542 8327 13598 8336
rect 13360 8288 13412 8294
rect 13360 8230 13412 8236
rect 13452 7880 13504 7886
rect 13452 7822 13504 7828
rect 13360 6792 13412 6798
rect 13360 6734 13412 6740
rect 13268 5296 13320 5302
rect 13268 5238 13320 5244
rect 13372 4865 13400 6734
rect 13464 6322 13492 7822
rect 13544 7336 13596 7342
rect 13648 7324 13676 8366
rect 13820 7472 13872 7478
rect 13820 7414 13872 7420
rect 13596 7296 13676 7324
rect 13544 7278 13596 7284
rect 13542 6624 13598 6633
rect 13542 6559 13598 6568
rect 13452 6316 13504 6322
rect 13452 6258 13504 6264
rect 13556 5681 13584 6559
rect 13648 6225 13676 7296
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13634 6216 13690 6225
rect 13634 6151 13690 6160
rect 13636 5840 13688 5846
rect 13636 5782 13688 5788
rect 13542 5672 13598 5681
rect 13542 5607 13598 5616
rect 13556 5574 13584 5607
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 13648 5386 13676 5782
rect 13556 5358 13676 5386
rect 13358 4856 13414 4865
rect 13358 4791 13414 4800
rect 13452 4752 13504 4758
rect 13452 4694 13504 4700
rect 13268 4276 13320 4282
rect 13268 4218 13320 4224
rect 13280 3097 13308 4218
rect 13358 4176 13414 4185
rect 13358 4111 13414 4120
rect 13372 3398 13400 4111
rect 13464 4078 13492 4694
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 13360 3392 13412 3398
rect 13360 3334 13412 3340
rect 13450 3224 13506 3233
rect 13360 3188 13412 3194
rect 13450 3159 13506 3168
rect 13360 3130 13412 3136
rect 13266 3088 13322 3097
rect 13266 3023 13322 3032
rect 13266 2952 13322 2961
rect 13266 2887 13268 2896
rect 13320 2887 13322 2896
rect 13268 2858 13320 2864
rect 13096 2746 13216 2774
rect 13266 2816 13322 2825
rect 13266 2751 13322 2760
rect 12808 2644 12860 2650
rect 12808 2586 12860 2592
rect 12716 2372 12768 2378
rect 12716 2314 12768 2320
rect 12624 1420 12676 1426
rect 12624 1362 12676 1368
rect 12544 870 12664 898
rect 12636 800 12664 870
rect 12728 800 12756 2314
rect 12820 800 12848 2586
rect 12990 2408 13046 2417
rect 12990 2343 13046 2352
rect 13004 2310 13032 2343
rect 12992 2304 13044 2310
rect 12992 2246 13044 2252
rect 13096 1442 13124 2746
rect 13176 2440 13228 2446
rect 13176 2382 13228 2388
rect 13188 2106 13216 2382
rect 13176 2100 13228 2106
rect 13176 2042 13228 2048
rect 13004 1414 13124 1442
rect 13176 1420 13228 1426
rect 12900 944 12952 950
rect 12900 886 12952 892
rect 12912 800 12940 886
rect 13004 800 13032 1414
rect 13176 1362 13228 1368
rect 13084 1352 13136 1358
rect 13084 1294 13136 1300
rect 13096 800 13124 1294
rect 13188 800 13216 1362
rect 13280 800 13308 2751
rect 13372 800 13400 3130
rect 13464 800 13492 3159
rect 13556 3058 13584 5358
rect 13636 5092 13688 5098
rect 13636 5034 13688 5040
rect 13648 4690 13676 5034
rect 13740 5001 13768 6734
rect 13832 5846 13860 7414
rect 14004 7404 14056 7410
rect 14004 7346 14056 7352
rect 14016 7206 14044 7346
rect 13912 7200 13964 7206
rect 13912 7142 13964 7148
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 13820 5840 13872 5846
rect 13820 5782 13872 5788
rect 13924 5302 13952 7142
rect 14200 5710 14228 9862
rect 14292 9722 14320 10610
rect 14280 9716 14332 9722
rect 14280 9658 14332 9664
rect 14384 9625 14412 12174
rect 14370 9616 14426 9625
rect 14370 9551 14426 9560
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 14292 8634 14320 8910
rect 14280 8628 14332 8634
rect 14280 8570 14332 8576
rect 14292 7410 14320 8570
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14476 6474 14504 14198
rect 14752 13530 14780 21898
rect 15028 21690 15056 22066
rect 15120 21962 15148 22918
rect 15292 22432 15344 22438
rect 15292 22374 15344 22380
rect 15304 22273 15332 22374
rect 15290 22264 15346 22273
rect 15290 22199 15346 22208
rect 15764 22094 15792 23258
rect 16040 23050 16068 24822
rect 16028 23044 16080 23050
rect 16028 22986 16080 22992
rect 15844 22976 15896 22982
rect 15844 22918 15896 22924
rect 15856 22642 15884 22918
rect 15844 22636 15896 22642
rect 15844 22578 15896 22584
rect 15856 22166 15884 22578
rect 15936 22432 15988 22438
rect 15936 22374 15988 22380
rect 15948 22234 15976 22374
rect 15936 22228 15988 22234
rect 15936 22170 15988 22176
rect 15844 22160 15896 22166
rect 15844 22102 15896 22108
rect 15672 22066 15792 22094
rect 15108 21956 15160 21962
rect 15108 21898 15160 21904
rect 15016 21684 15068 21690
rect 15016 21626 15068 21632
rect 15028 20890 15056 21626
rect 14844 20862 15056 20890
rect 15476 20936 15528 20942
rect 15476 20878 15528 20884
rect 15384 20868 15436 20874
rect 14740 13524 14792 13530
rect 14740 13466 14792 13472
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14568 12238 14596 13262
rect 14844 13190 14872 20862
rect 15384 20810 15436 20816
rect 15016 20800 15068 20806
rect 15016 20742 15068 20748
rect 15028 19854 15056 20742
rect 15396 20602 15424 20810
rect 15384 20596 15436 20602
rect 15384 20538 15436 20544
rect 15488 19922 15516 20878
rect 15568 20392 15620 20398
rect 15568 20334 15620 20340
rect 15476 19916 15528 19922
rect 15476 19858 15528 19864
rect 15016 19848 15068 19854
rect 15016 19790 15068 19796
rect 14924 19780 14976 19786
rect 14924 19722 14976 19728
rect 14936 19446 14964 19722
rect 14924 19440 14976 19446
rect 14924 19382 14976 19388
rect 15028 16114 15056 19790
rect 15384 19168 15436 19174
rect 15384 19110 15436 19116
rect 15396 18698 15424 19110
rect 15488 18766 15516 19858
rect 15580 19310 15608 20334
rect 15568 19304 15620 19310
rect 15568 19246 15620 19252
rect 15476 18760 15528 18766
rect 15476 18702 15528 18708
rect 15384 18692 15436 18698
rect 15384 18634 15436 18640
rect 15292 18284 15344 18290
rect 15292 18226 15344 18232
rect 15200 16788 15252 16794
rect 15200 16730 15252 16736
rect 15016 16108 15068 16114
rect 15016 16050 15068 16056
rect 15212 15162 15240 16730
rect 15304 16046 15332 18226
rect 15292 16040 15344 16046
rect 15292 15982 15344 15988
rect 15200 15156 15252 15162
rect 15200 15098 15252 15104
rect 15304 14414 15332 15982
rect 15384 15972 15436 15978
rect 15384 15914 15436 15920
rect 15396 14482 15424 15914
rect 15672 15706 15700 22066
rect 15856 21554 15884 22102
rect 15844 21548 15896 21554
rect 15844 21490 15896 21496
rect 16028 20528 16080 20534
rect 16028 20470 16080 20476
rect 15752 20460 15804 20466
rect 15752 20402 15804 20408
rect 15764 20262 15792 20402
rect 15844 20324 15896 20330
rect 15844 20266 15896 20272
rect 15752 20256 15804 20262
rect 15752 20198 15804 20204
rect 15856 20097 15884 20266
rect 15842 20088 15898 20097
rect 16040 20058 16068 20470
rect 16132 20058 16160 24890
rect 16224 24886 16252 27814
rect 16316 27538 16344 29106
rect 16396 28756 16448 28762
rect 16396 28698 16448 28704
rect 16304 27532 16356 27538
rect 16304 27474 16356 27480
rect 16316 27062 16344 27474
rect 16304 27056 16356 27062
rect 16304 26998 16356 27004
rect 16212 24880 16264 24886
rect 16212 24822 16264 24828
rect 16212 23656 16264 23662
rect 16212 23598 16264 23604
rect 16224 20262 16252 23598
rect 16408 22438 16436 28698
rect 16488 28484 16540 28490
rect 16488 28426 16540 28432
rect 16500 27470 16528 28426
rect 16592 27878 16620 29106
rect 16764 28552 16816 28558
rect 16764 28494 16816 28500
rect 16948 28552 17000 28558
rect 16948 28494 17000 28500
rect 16776 28218 16804 28494
rect 16764 28212 16816 28218
rect 16764 28154 16816 28160
rect 16960 28150 16988 28494
rect 16948 28144 17000 28150
rect 16948 28086 17000 28092
rect 16580 27872 16632 27878
rect 16580 27814 16632 27820
rect 16488 27464 16540 27470
rect 16488 27406 16540 27412
rect 16592 24070 16620 27814
rect 17052 27674 17080 29650
rect 17144 29578 17172 30262
rect 17314 30152 17370 30161
rect 17314 30087 17370 30096
rect 17328 29646 17356 30087
rect 17316 29640 17368 29646
rect 17316 29582 17368 29588
rect 17132 29572 17184 29578
rect 17132 29514 17184 29520
rect 17144 29458 17172 29514
rect 17144 29430 17264 29458
rect 17236 29238 17264 29430
rect 17224 29232 17276 29238
rect 17224 29174 17276 29180
rect 17420 29170 17448 30534
rect 18236 30388 18288 30394
rect 18236 30330 18288 30336
rect 18052 30048 18104 30054
rect 18052 29990 18104 29996
rect 18064 29646 18092 29990
rect 18248 29646 18276 30330
rect 19444 30036 19472 30602
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19996 30326 20024 31078
rect 19984 30320 20036 30326
rect 19984 30262 20036 30268
rect 20088 30138 20116 31214
rect 21376 30598 21404 31690
rect 21364 30592 21416 30598
rect 21364 30534 21416 30540
rect 19996 30110 20116 30138
rect 19524 30048 19576 30054
rect 19444 30008 19524 30036
rect 19524 29990 19576 29996
rect 19536 29850 19564 29990
rect 19524 29844 19576 29850
rect 19524 29786 19576 29792
rect 18052 29640 18104 29646
rect 18052 29582 18104 29588
rect 18236 29640 18288 29646
rect 18236 29582 18288 29588
rect 18512 29640 18564 29646
rect 18512 29582 18564 29588
rect 19248 29640 19300 29646
rect 19248 29582 19300 29588
rect 19614 29608 19670 29617
rect 17500 29232 17552 29238
rect 17500 29174 17552 29180
rect 17132 29164 17184 29170
rect 17132 29106 17184 29112
rect 17408 29164 17460 29170
rect 17408 29106 17460 29112
rect 17144 29073 17172 29106
rect 17130 29064 17186 29073
rect 17130 28999 17186 29008
rect 17408 28416 17460 28422
rect 17408 28358 17460 28364
rect 17040 27668 17092 27674
rect 17040 27610 17092 27616
rect 17224 27464 17276 27470
rect 17224 27406 17276 27412
rect 17040 27396 17092 27402
rect 17040 27338 17092 27344
rect 17132 27396 17184 27402
rect 17132 27338 17184 27344
rect 16672 26988 16724 26994
rect 16672 26930 16724 26936
rect 16684 26518 16712 26930
rect 16948 26852 17000 26858
rect 16948 26794 17000 26800
rect 16672 26512 16724 26518
rect 16672 26454 16724 26460
rect 16672 26240 16724 26246
rect 16672 26182 16724 26188
rect 16684 25838 16712 26182
rect 16672 25832 16724 25838
rect 16672 25774 16724 25780
rect 16580 24064 16632 24070
rect 16580 24006 16632 24012
rect 16396 22432 16448 22438
rect 16396 22374 16448 22380
rect 16684 22094 16712 25774
rect 16960 25294 16988 26794
rect 17052 26382 17080 27338
rect 17144 26897 17172 27338
rect 17130 26888 17186 26897
rect 17130 26823 17186 26832
rect 17236 26382 17264 27406
rect 17420 26790 17448 28358
rect 17512 27130 17540 29174
rect 18524 28966 18552 29582
rect 19064 29572 19116 29578
rect 19064 29514 19116 29520
rect 18604 29504 18656 29510
rect 18604 29446 18656 29452
rect 18616 29170 18644 29446
rect 18604 29164 18656 29170
rect 18604 29106 18656 29112
rect 18880 29096 18932 29102
rect 19076 29050 19104 29514
rect 19156 29504 19208 29510
rect 19156 29446 19208 29452
rect 18932 29044 19104 29050
rect 18880 29038 19104 29044
rect 18892 29022 19104 29038
rect 17960 28960 18012 28966
rect 17960 28902 18012 28908
rect 18512 28960 18564 28966
rect 18512 28902 18564 28908
rect 17972 28558 18000 28902
rect 17960 28552 18012 28558
rect 17960 28494 18012 28500
rect 19076 28490 19104 29022
rect 19064 28484 19116 28490
rect 19064 28426 19116 28432
rect 18972 28076 19024 28082
rect 18972 28018 19024 28024
rect 17960 27872 18012 27878
rect 17960 27814 18012 27820
rect 17684 27668 17736 27674
rect 17684 27610 17736 27616
rect 17500 27124 17552 27130
rect 17500 27066 17552 27072
rect 17512 26994 17540 27066
rect 17500 26988 17552 26994
rect 17500 26930 17552 26936
rect 17408 26784 17460 26790
rect 17408 26726 17460 26732
rect 17408 26512 17460 26518
rect 17408 26454 17460 26460
rect 17040 26376 17092 26382
rect 17040 26318 17092 26324
rect 17224 26376 17276 26382
rect 17420 26353 17448 26454
rect 17224 26318 17276 26324
rect 17406 26344 17462 26353
rect 17052 25906 17080 26318
rect 17132 26308 17184 26314
rect 17132 26250 17184 26256
rect 17040 25900 17092 25906
rect 17040 25842 17092 25848
rect 17144 25770 17172 26250
rect 17132 25764 17184 25770
rect 17132 25706 17184 25712
rect 17236 25362 17264 26318
rect 17406 26279 17462 26288
rect 17696 26234 17724 27610
rect 17776 27328 17828 27334
rect 17828 27288 17908 27316
rect 17776 27270 17828 27276
rect 17776 26376 17828 26382
rect 17776 26318 17828 26324
rect 17604 26206 17724 26234
rect 17316 25900 17368 25906
rect 17316 25842 17368 25848
rect 17224 25356 17276 25362
rect 17144 25316 17224 25344
rect 16948 25288 17000 25294
rect 16948 25230 17000 25236
rect 17040 24608 17092 24614
rect 17040 24550 17092 24556
rect 17052 24206 17080 24550
rect 17144 24206 17172 25316
rect 17224 25298 17276 25304
rect 17328 25294 17356 25842
rect 17316 25288 17368 25294
rect 17316 25230 17368 25236
rect 17406 25256 17462 25265
rect 17224 24336 17276 24342
rect 17224 24278 17276 24284
rect 17040 24200 17092 24206
rect 17040 24142 17092 24148
rect 17132 24200 17184 24206
rect 17132 24142 17184 24148
rect 17236 23526 17264 24278
rect 17328 24154 17356 25230
rect 17406 25191 17408 25200
rect 17460 25191 17462 25200
rect 17408 25162 17460 25168
rect 17604 24290 17632 26206
rect 17788 25362 17816 26318
rect 17776 25356 17828 25362
rect 17776 25298 17828 25304
rect 17684 25152 17736 25158
rect 17684 25094 17736 25100
rect 17696 24993 17724 25094
rect 17682 24984 17738 24993
rect 17682 24919 17738 24928
rect 17604 24262 17724 24290
rect 17592 24200 17644 24206
rect 17328 24138 17448 24154
rect 17592 24142 17644 24148
rect 17328 24132 17460 24138
rect 17328 24126 17408 24132
rect 17408 24074 17460 24080
rect 17500 24132 17552 24138
rect 17500 24074 17552 24080
rect 17314 23760 17370 23769
rect 17420 23730 17448 24074
rect 17314 23695 17316 23704
rect 17368 23695 17370 23704
rect 17408 23724 17460 23730
rect 17316 23666 17368 23672
rect 17408 23666 17460 23672
rect 17512 23594 17540 24074
rect 17604 23730 17632 24142
rect 17592 23724 17644 23730
rect 17592 23666 17644 23672
rect 17500 23588 17552 23594
rect 17500 23530 17552 23536
rect 17224 23520 17276 23526
rect 17224 23462 17276 23468
rect 17040 23044 17092 23050
rect 17040 22986 17092 22992
rect 16592 22066 16712 22094
rect 16592 21962 16620 22066
rect 16580 21956 16632 21962
rect 16580 21898 16632 21904
rect 16592 21690 16620 21898
rect 16580 21684 16632 21690
rect 16580 21626 16632 21632
rect 16948 21548 17000 21554
rect 16948 21490 17000 21496
rect 16960 21146 16988 21490
rect 16948 21140 17000 21146
rect 16948 21082 17000 21088
rect 17052 21078 17080 22986
rect 17236 22094 17264 23462
rect 17604 23254 17632 23666
rect 17500 23248 17552 23254
rect 17500 23190 17552 23196
rect 17592 23248 17644 23254
rect 17592 23190 17644 23196
rect 17512 22642 17540 23190
rect 17592 23112 17644 23118
rect 17592 23054 17644 23060
rect 17500 22636 17552 22642
rect 17500 22578 17552 22584
rect 17236 22066 17356 22094
rect 17224 21888 17276 21894
rect 17224 21830 17276 21836
rect 17040 21072 17092 21078
rect 17040 21014 17092 21020
rect 16304 20868 16356 20874
rect 16304 20810 16356 20816
rect 16212 20256 16264 20262
rect 16212 20198 16264 20204
rect 15842 20023 15898 20032
rect 16028 20052 16080 20058
rect 16028 19994 16080 20000
rect 16120 20052 16172 20058
rect 16120 19994 16172 20000
rect 16132 19258 16160 19994
rect 16224 19854 16252 20198
rect 16212 19848 16264 19854
rect 16212 19790 16264 19796
rect 15948 19230 16160 19258
rect 15844 18964 15896 18970
rect 15844 18906 15896 18912
rect 15752 18692 15804 18698
rect 15752 18634 15804 18640
rect 15764 16046 15792 18634
rect 15856 18358 15884 18906
rect 15844 18352 15896 18358
rect 15844 18294 15896 18300
rect 15948 18170 15976 19230
rect 16120 18352 16172 18358
rect 16120 18294 16172 18300
rect 15856 18142 15976 18170
rect 15856 17338 15884 18142
rect 16028 17672 16080 17678
rect 16028 17614 16080 17620
rect 16040 17542 16068 17614
rect 15936 17536 15988 17542
rect 15936 17478 15988 17484
rect 16028 17536 16080 17542
rect 16028 17478 16080 17484
rect 15844 17332 15896 17338
rect 15844 17274 15896 17280
rect 15948 17270 15976 17478
rect 15936 17264 15988 17270
rect 15842 17232 15898 17241
rect 15936 17206 15988 17212
rect 15842 17167 15844 17176
rect 15896 17167 15898 17176
rect 15844 17138 15896 17144
rect 15844 16652 15896 16658
rect 15844 16594 15896 16600
rect 15752 16040 15804 16046
rect 15752 15982 15804 15988
rect 15660 15700 15712 15706
rect 15660 15642 15712 15648
rect 15476 15428 15528 15434
rect 15476 15370 15528 15376
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 15108 13456 15160 13462
rect 15108 13398 15160 13404
rect 14832 13184 14884 13190
rect 14832 13126 14884 13132
rect 15120 12714 15148 13398
rect 15212 13326 15240 13806
rect 15304 13394 15332 14350
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 15200 13320 15252 13326
rect 15200 13262 15252 13268
rect 15212 12918 15240 13262
rect 15396 13002 15424 14418
rect 15304 12974 15424 13002
rect 15200 12912 15252 12918
rect 15200 12854 15252 12860
rect 14648 12708 14700 12714
rect 14648 12650 14700 12656
rect 15108 12708 15160 12714
rect 15108 12650 15160 12656
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 14384 6446 14504 6474
rect 14188 5704 14240 5710
rect 14188 5646 14240 5652
rect 14384 5574 14412 6446
rect 14556 6112 14608 6118
rect 14556 6054 14608 6060
rect 14372 5568 14424 5574
rect 14372 5510 14424 5516
rect 13912 5296 13964 5302
rect 13912 5238 13964 5244
rect 14096 5228 14148 5234
rect 14096 5170 14148 5176
rect 13912 5160 13964 5166
rect 13912 5102 13964 5108
rect 13820 5092 13872 5098
rect 13820 5034 13872 5040
rect 13726 4992 13782 5001
rect 13726 4927 13782 4936
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 13636 4684 13688 4690
rect 13636 4626 13688 4632
rect 13648 4554 13676 4626
rect 13636 4548 13688 4554
rect 13636 4490 13688 4496
rect 13740 4146 13768 4762
rect 13832 4758 13860 5034
rect 13820 4752 13872 4758
rect 13820 4694 13872 4700
rect 13924 4622 13952 5102
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 13912 4616 13964 4622
rect 13912 4558 13964 4564
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 13726 4040 13782 4049
rect 13924 4010 13952 4558
rect 13726 3975 13782 3984
rect 13912 4004 13964 4010
rect 13544 3052 13596 3058
rect 13544 2994 13596 3000
rect 13556 2514 13584 2994
rect 13636 2916 13688 2922
rect 13636 2858 13688 2864
rect 13544 2508 13596 2514
rect 13544 2450 13596 2456
rect 13544 2372 13596 2378
rect 13544 2314 13596 2320
rect 13556 1426 13584 2314
rect 13544 1420 13596 1426
rect 13544 1362 13596 1368
rect 13544 1284 13596 1290
rect 13544 1226 13596 1232
rect 13556 800 13584 1226
rect 13648 800 13676 2858
rect 13740 2378 13768 3975
rect 13912 3946 13964 3952
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 13832 3210 13860 3878
rect 13832 3182 13952 3210
rect 13820 3120 13872 3126
rect 13820 3062 13872 3068
rect 13728 2372 13780 2378
rect 13728 2314 13780 2320
rect 13740 2038 13768 2314
rect 13728 2032 13780 2038
rect 13728 1974 13780 1980
rect 13832 800 13860 3062
rect 13924 3058 13952 3182
rect 13912 3052 13964 3058
rect 13912 2994 13964 3000
rect 14016 2774 14044 4966
rect 14108 4758 14136 5170
rect 14384 5166 14412 5510
rect 14372 5160 14424 5166
rect 14372 5102 14424 5108
rect 14096 4752 14148 4758
rect 14096 4694 14148 4700
rect 14108 4078 14136 4694
rect 14384 4282 14412 5102
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 14372 4276 14424 4282
rect 14372 4218 14424 4224
rect 14096 4072 14148 4078
rect 14096 4014 14148 4020
rect 14108 3738 14136 4014
rect 14096 3732 14148 3738
rect 14096 3674 14148 3680
rect 14372 3732 14424 3738
rect 14372 3674 14424 3680
rect 14384 3641 14412 3674
rect 14370 3632 14426 3641
rect 14370 3567 14426 3576
rect 14476 3534 14504 4558
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14280 3460 14332 3466
rect 14280 3402 14332 3408
rect 14292 2990 14320 3402
rect 14372 3392 14424 3398
rect 14372 3334 14424 3340
rect 14280 2984 14332 2990
rect 14280 2926 14332 2932
rect 14188 2848 14240 2854
rect 14188 2790 14240 2796
rect 13924 2746 14044 2774
rect 13924 800 13952 2746
rect 14096 2304 14148 2310
rect 14096 2246 14148 2252
rect 14108 800 14136 2246
rect 14200 800 14228 2790
rect 14384 800 14412 3334
rect 14568 3058 14596 6054
rect 14660 5370 14688 12650
rect 15212 12594 15240 12854
rect 15120 12566 15240 12594
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 14752 8974 14780 9454
rect 15016 9036 15068 9042
rect 15016 8978 15068 8984
rect 14740 8968 14792 8974
rect 14740 8910 14792 8916
rect 14924 7812 14976 7818
rect 14924 7754 14976 7760
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14752 7392 14780 7686
rect 14936 7546 14964 7754
rect 14924 7540 14976 7546
rect 14924 7482 14976 7488
rect 14832 7404 14884 7410
rect 14752 7364 14832 7392
rect 14832 7346 14884 7352
rect 14740 7200 14792 7206
rect 14740 7142 14792 7148
rect 14648 5364 14700 5370
rect 14648 5306 14700 5312
rect 14752 5250 14780 7142
rect 14660 5222 14780 5250
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 14464 2576 14516 2582
rect 14464 2518 14516 2524
rect 14476 800 14504 2518
rect 14660 800 14688 5222
rect 14740 5092 14792 5098
rect 14740 5034 14792 5040
rect 14752 4690 14780 5034
rect 14740 4684 14792 4690
rect 14740 4626 14792 4632
rect 14740 3664 14792 3670
rect 14740 3606 14792 3612
rect 14752 800 14780 3606
rect 14844 3466 14872 7346
rect 14922 5672 14978 5681
rect 14922 5607 14978 5616
rect 14832 3460 14884 3466
rect 14832 3402 14884 3408
rect 14832 2644 14884 2650
rect 14832 2586 14884 2592
rect 14844 2553 14872 2586
rect 14830 2544 14886 2553
rect 14830 2479 14886 2488
rect 14936 2446 14964 5607
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 15028 800 15056 8978
rect 15120 7478 15148 12566
rect 15304 12374 15332 12974
rect 15384 12844 15436 12850
rect 15384 12786 15436 12792
rect 15292 12368 15344 12374
rect 15292 12310 15344 12316
rect 15396 12170 15424 12786
rect 15488 12374 15516 15370
rect 15752 14340 15804 14346
rect 15752 14282 15804 14288
rect 15568 13932 15620 13938
rect 15568 13874 15620 13880
rect 15580 12850 15608 13874
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 15764 12714 15792 14282
rect 15752 12708 15804 12714
rect 15752 12650 15804 12656
rect 15476 12368 15528 12374
rect 15476 12310 15528 12316
rect 15384 12164 15436 12170
rect 15384 12106 15436 12112
rect 15856 11830 15884 16594
rect 15948 14414 15976 17206
rect 16040 16794 16068 17478
rect 16028 16788 16080 16794
rect 16028 16730 16080 16736
rect 16132 14482 16160 18294
rect 16224 16658 16252 19790
rect 16212 16652 16264 16658
rect 16212 16594 16264 16600
rect 16120 14476 16172 14482
rect 16120 14418 16172 14424
rect 15936 14408 15988 14414
rect 15936 14350 15988 14356
rect 16132 14006 16160 14418
rect 16120 14000 16172 14006
rect 16120 13942 16172 13948
rect 16316 13376 16344 20810
rect 16396 20596 16448 20602
rect 16396 20538 16448 20544
rect 16408 20398 16436 20538
rect 16948 20460 17000 20466
rect 17052 20448 17080 21014
rect 17000 20420 17080 20448
rect 16948 20402 17000 20408
rect 16396 20392 16448 20398
rect 16396 20334 16448 20340
rect 16408 19378 16436 20334
rect 16672 20256 16724 20262
rect 16672 20198 16724 20204
rect 16488 19984 16540 19990
rect 16488 19926 16540 19932
rect 16500 19446 16528 19926
rect 16684 19854 16712 20198
rect 16672 19848 16724 19854
rect 16672 19790 16724 19796
rect 16856 19508 16908 19514
rect 16856 19450 16908 19456
rect 16488 19440 16540 19446
rect 16488 19382 16540 19388
rect 16396 19372 16448 19378
rect 16396 19314 16448 19320
rect 16396 19236 16448 19242
rect 16396 19178 16448 19184
rect 16408 18766 16436 19178
rect 16396 18760 16448 18766
rect 16396 18702 16448 18708
rect 16672 18760 16724 18766
rect 16672 18702 16724 18708
rect 16764 18760 16816 18766
rect 16764 18702 16816 18708
rect 16684 18426 16712 18702
rect 16672 18420 16724 18426
rect 16672 18362 16724 18368
rect 16776 18306 16804 18702
rect 16500 18290 16804 18306
rect 16488 18284 16804 18290
rect 16540 18278 16804 18284
rect 16488 18226 16540 18232
rect 16396 18216 16448 18222
rect 16396 18158 16448 18164
rect 16408 16046 16436 18158
rect 16776 18154 16804 18278
rect 16764 18148 16816 18154
rect 16764 18090 16816 18096
rect 16868 17678 16896 19450
rect 16948 18624 17000 18630
rect 16948 18566 17000 18572
rect 16960 18358 16988 18566
rect 16948 18352 17000 18358
rect 16948 18294 17000 18300
rect 17130 18320 17186 18329
rect 17130 18255 17132 18264
rect 17184 18255 17186 18264
rect 17132 18226 17184 18232
rect 17132 18080 17184 18086
rect 17132 18022 17184 18028
rect 16856 17672 16908 17678
rect 16856 17614 16908 17620
rect 17040 17672 17092 17678
rect 17040 17614 17092 17620
rect 16672 17196 16724 17202
rect 16672 17138 16724 17144
rect 16684 16726 16712 17138
rect 16868 17134 16896 17614
rect 17052 17338 17080 17614
rect 17040 17332 17092 17338
rect 17040 17274 17092 17280
rect 16856 17128 16908 17134
rect 16856 17070 16908 17076
rect 16672 16720 16724 16726
rect 16672 16662 16724 16668
rect 16684 16182 16712 16662
rect 16764 16448 16816 16454
rect 16764 16390 16816 16396
rect 16672 16176 16724 16182
rect 16672 16118 16724 16124
rect 16396 16040 16448 16046
rect 16396 15982 16448 15988
rect 16408 14278 16436 15982
rect 16488 15496 16540 15502
rect 16488 15438 16540 15444
rect 16500 15026 16528 15438
rect 16776 15026 16804 16390
rect 16488 15020 16540 15026
rect 16488 14962 16540 14968
rect 16764 15020 16816 15026
rect 16764 14962 16816 14968
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 16672 14272 16724 14278
rect 16672 14214 16724 14220
rect 16684 13938 16712 14214
rect 16672 13932 16724 13938
rect 16672 13874 16724 13880
rect 16580 13864 16632 13870
rect 16578 13832 16580 13841
rect 16632 13832 16634 13841
rect 16578 13767 16634 13776
rect 16672 13728 16724 13734
rect 16670 13696 16672 13705
rect 16724 13696 16726 13705
rect 16670 13631 16726 13640
rect 16764 13456 16816 13462
rect 16762 13424 16764 13433
rect 16816 13424 16818 13433
rect 16316 13348 16436 13376
rect 16762 13359 16818 13368
rect 16304 13252 16356 13258
rect 16304 13194 16356 13200
rect 16316 12986 16344 13194
rect 16304 12980 16356 12986
rect 16304 12922 16356 12928
rect 16212 12436 16264 12442
rect 16212 12378 16264 12384
rect 16224 12238 16252 12378
rect 16212 12232 16264 12238
rect 16212 12174 16264 12180
rect 16408 11898 16436 13348
rect 16868 12782 16896 17070
rect 17040 16584 17092 16590
rect 17040 16526 17092 16532
rect 17052 16250 17080 16526
rect 17040 16244 17092 16250
rect 17040 16186 17092 16192
rect 17144 14414 17172 18022
rect 17236 14618 17264 21830
rect 17328 19310 17356 22066
rect 17512 19514 17540 22578
rect 17604 22030 17632 23054
rect 17592 22024 17644 22030
rect 17592 21966 17644 21972
rect 17696 21690 17724 24262
rect 17776 24064 17828 24070
rect 17776 24006 17828 24012
rect 17684 21684 17736 21690
rect 17684 21626 17736 21632
rect 17592 21548 17644 21554
rect 17592 21490 17644 21496
rect 17604 20874 17632 21490
rect 17684 21140 17736 21146
rect 17684 21082 17736 21088
rect 17592 20868 17644 20874
rect 17592 20810 17644 20816
rect 17592 20460 17644 20466
rect 17592 20402 17644 20408
rect 17604 19786 17632 20402
rect 17592 19780 17644 19786
rect 17592 19722 17644 19728
rect 17500 19508 17552 19514
rect 17500 19450 17552 19456
rect 17316 19304 17368 19310
rect 17316 19246 17368 19252
rect 17328 18766 17356 19246
rect 17316 18760 17368 18766
rect 17316 18702 17368 18708
rect 17500 18760 17552 18766
rect 17500 18702 17552 18708
rect 17408 18624 17460 18630
rect 17408 18566 17460 18572
rect 17316 18284 17368 18290
rect 17316 18226 17368 18232
rect 17328 18193 17356 18226
rect 17314 18184 17370 18193
rect 17314 18119 17370 18128
rect 17420 18034 17448 18566
rect 17328 18006 17448 18034
rect 17328 17678 17356 18006
rect 17408 17740 17460 17746
rect 17408 17682 17460 17688
rect 17316 17672 17368 17678
rect 17316 17614 17368 17620
rect 17328 16658 17356 17614
rect 17316 16652 17368 16658
rect 17316 16594 17368 16600
rect 17420 16522 17448 17682
rect 17408 16516 17460 16522
rect 17408 16458 17460 16464
rect 17224 14612 17276 14618
rect 17224 14554 17276 14560
rect 17132 14408 17184 14414
rect 17132 14350 17184 14356
rect 17132 14272 17184 14278
rect 17132 14214 17184 14220
rect 16856 12776 16908 12782
rect 16856 12718 16908 12724
rect 17144 12434 17172 14214
rect 17512 13734 17540 18702
rect 17592 15088 17644 15094
rect 17592 15030 17644 15036
rect 17500 13728 17552 13734
rect 17500 13670 17552 13676
rect 17512 13530 17540 13670
rect 17500 13524 17552 13530
rect 17500 13466 17552 13472
rect 17500 12776 17552 12782
rect 17500 12718 17552 12724
rect 17224 12640 17276 12646
rect 17224 12582 17276 12588
rect 16868 12406 17172 12434
rect 16396 11892 16448 11898
rect 16396 11834 16448 11840
rect 15844 11824 15896 11830
rect 15844 11766 15896 11772
rect 15844 11552 15896 11558
rect 15844 11494 15896 11500
rect 15200 11076 15252 11082
rect 15200 11018 15252 11024
rect 15212 10810 15240 11018
rect 15200 10804 15252 10810
rect 15200 10746 15252 10752
rect 15856 10062 15884 11494
rect 16408 11354 16436 11834
rect 16396 11348 16448 11354
rect 16396 11290 16448 11296
rect 16396 10736 16448 10742
rect 16396 10678 16448 10684
rect 16304 10668 16356 10674
rect 16304 10610 16356 10616
rect 16316 10062 16344 10610
rect 15844 10056 15896 10062
rect 15844 9998 15896 10004
rect 16304 10056 16356 10062
rect 16304 9998 16356 10004
rect 15476 9920 15528 9926
rect 15476 9862 15528 9868
rect 15292 9512 15344 9518
rect 15292 9454 15344 9460
rect 15304 9178 15332 9454
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 15396 8974 15424 9318
rect 15384 8968 15436 8974
rect 15384 8910 15436 8916
rect 15292 8424 15344 8430
rect 15292 8366 15344 8372
rect 15108 7472 15160 7478
rect 15108 7414 15160 7420
rect 15120 4214 15148 7414
rect 15200 6180 15252 6186
rect 15200 6122 15252 6128
rect 15212 5234 15240 6122
rect 15200 5228 15252 5234
rect 15200 5170 15252 5176
rect 15108 4208 15160 4214
rect 15108 4150 15160 4156
rect 15108 4072 15160 4078
rect 15108 4014 15160 4020
rect 15120 3913 15148 4014
rect 15200 3936 15252 3942
rect 15106 3904 15162 3913
rect 15200 3878 15252 3884
rect 15106 3839 15162 3848
rect 15212 3670 15240 3878
rect 15200 3664 15252 3670
rect 15200 3606 15252 3612
rect 15108 3460 15160 3466
rect 15108 3402 15160 3408
rect 15120 3126 15148 3402
rect 15108 3120 15160 3126
rect 15108 3062 15160 3068
rect 15304 800 15332 8366
rect 15488 7018 15516 9862
rect 15568 9580 15620 9586
rect 15568 9522 15620 9528
rect 15580 9178 15608 9522
rect 15568 9172 15620 9178
rect 15568 9114 15620 9120
rect 15856 8430 15884 9998
rect 16408 9586 16436 10678
rect 16396 9580 16448 9586
rect 16396 9522 16448 9528
rect 16408 8498 16436 9522
rect 16868 9489 16896 12406
rect 17040 11552 17092 11558
rect 17040 11494 17092 11500
rect 17052 10724 17080 11494
rect 17132 10736 17184 10742
rect 17052 10696 17132 10724
rect 16948 9512 17000 9518
rect 16854 9480 16910 9489
rect 16948 9454 17000 9460
rect 16854 9415 16910 9424
rect 16764 8900 16816 8906
rect 16764 8842 16816 8848
rect 16396 8492 16448 8498
rect 16396 8434 16448 8440
rect 15844 8424 15896 8430
rect 15844 8366 15896 8372
rect 15488 6990 15608 7018
rect 15476 6860 15528 6866
rect 15476 6802 15528 6808
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 15396 4146 15424 5646
rect 15384 4140 15436 4146
rect 15384 4082 15436 4088
rect 15488 2774 15516 6802
rect 15580 4570 15608 6990
rect 15752 6792 15804 6798
rect 15752 6734 15804 6740
rect 15660 6248 15712 6254
rect 15660 6190 15712 6196
rect 15672 5914 15700 6190
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 15580 4542 15700 4570
rect 15568 4480 15620 4486
rect 15568 4422 15620 4428
rect 15580 4146 15608 4422
rect 15568 4140 15620 4146
rect 15568 4082 15620 4088
rect 15672 3534 15700 4542
rect 15660 3528 15712 3534
rect 15660 3470 15712 3476
rect 15764 2774 15792 6734
rect 15856 4486 15884 8366
rect 16212 8288 16264 8294
rect 16212 8230 16264 8236
rect 16120 7200 16172 7206
rect 16120 7142 16172 7148
rect 15936 6724 15988 6730
rect 15936 6666 15988 6672
rect 15948 6322 15976 6666
rect 15936 6316 15988 6322
rect 15936 6258 15988 6264
rect 15936 5568 15988 5574
rect 15936 5510 15988 5516
rect 15948 4690 15976 5510
rect 16026 4720 16082 4729
rect 15936 4684 15988 4690
rect 16026 4655 16028 4664
rect 15936 4626 15988 4632
rect 16080 4655 16082 4664
rect 16028 4626 16080 4632
rect 15844 4480 15896 4486
rect 15844 4422 15896 4428
rect 15856 3738 15884 4422
rect 15948 4010 15976 4626
rect 15936 4004 15988 4010
rect 15936 3946 15988 3952
rect 15844 3732 15896 3738
rect 15844 3674 15896 3680
rect 15488 2746 15608 2774
rect 15764 2746 15884 2774
rect 15580 800 15608 2746
rect 15856 800 15884 2746
rect 16132 800 16160 7142
rect 16224 4282 16252 8230
rect 16408 7886 16436 8434
rect 16304 7880 16356 7886
rect 16304 7822 16356 7828
rect 16396 7880 16448 7886
rect 16396 7822 16448 7828
rect 16316 6866 16344 7822
rect 16672 7404 16724 7410
rect 16672 7346 16724 7352
rect 16684 7002 16712 7346
rect 16672 6996 16724 7002
rect 16672 6938 16724 6944
rect 16304 6860 16356 6866
rect 16304 6802 16356 6808
rect 16316 6458 16344 6802
rect 16396 6792 16448 6798
rect 16396 6734 16448 6740
rect 16304 6452 16356 6458
rect 16304 6394 16356 6400
rect 16212 4276 16264 4282
rect 16212 4218 16264 4224
rect 16408 800 16436 6734
rect 16672 6724 16724 6730
rect 16672 6666 16724 6672
rect 16684 5914 16712 6666
rect 16672 5908 16724 5914
rect 16672 5850 16724 5856
rect 16672 5704 16724 5710
rect 16672 5646 16724 5652
rect 16684 5302 16712 5646
rect 16672 5296 16724 5302
rect 16672 5238 16724 5244
rect 16488 3392 16540 3398
rect 16488 3334 16540 3340
rect 16500 3194 16528 3334
rect 16488 3188 16540 3194
rect 16488 3130 16540 3136
rect 16776 2774 16804 8842
rect 16960 7818 16988 9454
rect 17052 8362 17080 10696
rect 17132 10678 17184 10684
rect 17236 9654 17264 12582
rect 17512 12209 17540 12718
rect 17498 12200 17554 12209
rect 17498 12135 17554 12144
rect 17498 10976 17554 10985
rect 17498 10911 17554 10920
rect 17512 10266 17540 10911
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17604 10062 17632 15030
rect 17696 13569 17724 21082
rect 17682 13560 17738 13569
rect 17682 13495 17738 13504
rect 17592 10056 17644 10062
rect 17592 9998 17644 10004
rect 17224 9648 17276 9654
rect 17224 9590 17276 9596
rect 17682 9616 17738 9625
rect 17682 9551 17738 9560
rect 17132 9376 17184 9382
rect 17132 9318 17184 9324
rect 17316 9376 17368 9382
rect 17316 9318 17368 9324
rect 17144 9217 17172 9318
rect 17130 9208 17186 9217
rect 17130 9143 17186 9152
rect 17224 8832 17276 8838
rect 17224 8774 17276 8780
rect 17236 8362 17264 8774
rect 17040 8356 17092 8362
rect 17040 8298 17092 8304
rect 17224 8356 17276 8362
rect 17224 8298 17276 8304
rect 16948 7812 17000 7818
rect 16948 7754 17000 7760
rect 16856 6656 16908 6662
rect 16856 6598 16908 6604
rect 16868 5710 16896 6598
rect 16960 5760 16988 7754
rect 17052 6390 17080 8298
rect 17224 6724 17276 6730
rect 17224 6666 17276 6672
rect 17040 6384 17092 6390
rect 17040 6326 17092 6332
rect 16960 5732 17080 5760
rect 16856 5704 16908 5710
rect 16856 5646 16908 5652
rect 16868 3058 16896 5646
rect 17052 5642 17080 5732
rect 16948 5636 17000 5642
rect 16948 5578 17000 5584
rect 17040 5636 17092 5642
rect 17040 5578 17092 5584
rect 16960 5234 16988 5578
rect 17132 5568 17184 5574
rect 17132 5510 17184 5516
rect 17144 5370 17172 5510
rect 17132 5364 17184 5370
rect 17132 5306 17184 5312
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 17236 5114 17264 6666
rect 17328 5710 17356 9318
rect 17696 9178 17724 9551
rect 17788 9382 17816 24006
rect 17880 12646 17908 27288
rect 17972 27062 18000 27814
rect 18144 27464 18196 27470
rect 18144 27406 18196 27412
rect 18052 27396 18104 27402
rect 18052 27338 18104 27344
rect 17960 27056 18012 27062
rect 17960 26998 18012 27004
rect 17972 21962 18000 26998
rect 18064 26994 18092 27338
rect 18052 26988 18104 26994
rect 18052 26930 18104 26936
rect 18064 22098 18092 26930
rect 18156 26382 18184 27406
rect 18604 27328 18656 27334
rect 18604 27270 18656 27276
rect 18616 26994 18644 27270
rect 18984 27130 19012 28018
rect 19076 27470 19104 28426
rect 19064 27464 19116 27470
rect 19064 27406 19116 27412
rect 18972 27124 19024 27130
rect 18972 27066 19024 27072
rect 19064 27124 19116 27130
rect 19064 27066 19116 27072
rect 18604 26988 18656 26994
rect 18604 26930 18656 26936
rect 18420 26784 18472 26790
rect 18420 26726 18472 26732
rect 18144 26376 18196 26382
rect 18144 26318 18196 26324
rect 18144 25900 18196 25906
rect 18144 25842 18196 25848
rect 18156 24138 18184 25842
rect 18236 24608 18288 24614
rect 18236 24550 18288 24556
rect 18248 24206 18276 24550
rect 18328 24268 18380 24274
rect 18328 24210 18380 24216
rect 18236 24200 18288 24206
rect 18236 24142 18288 24148
rect 18144 24132 18196 24138
rect 18144 24074 18196 24080
rect 18156 23730 18184 24074
rect 18248 23769 18276 24142
rect 18340 23798 18368 24210
rect 18328 23792 18380 23798
rect 18234 23760 18290 23769
rect 18144 23724 18196 23730
rect 18328 23734 18380 23740
rect 18234 23695 18290 23704
rect 18144 23666 18196 23672
rect 18052 22092 18104 22098
rect 18156 22094 18184 23666
rect 18156 22066 18368 22094
rect 18052 22034 18104 22040
rect 17960 21956 18012 21962
rect 17960 21898 18012 21904
rect 18064 21690 18092 22034
rect 18340 22030 18368 22066
rect 18328 22024 18380 22030
rect 18328 21966 18380 21972
rect 18052 21684 18104 21690
rect 18052 21626 18104 21632
rect 18236 21072 18288 21078
rect 18236 21014 18288 21020
rect 18248 20466 18276 21014
rect 18328 20868 18380 20874
rect 18328 20810 18380 20816
rect 18340 20534 18368 20810
rect 18328 20528 18380 20534
rect 18328 20470 18380 20476
rect 18052 20460 18104 20466
rect 18052 20402 18104 20408
rect 18236 20460 18288 20466
rect 18236 20402 18288 20408
rect 18064 20346 18092 20402
rect 18064 20318 18184 20346
rect 18156 19718 18184 20318
rect 18144 19712 18196 19718
rect 18144 19654 18196 19660
rect 18052 19304 18104 19310
rect 18052 19246 18104 19252
rect 18064 18766 18092 19246
rect 18052 18760 18104 18766
rect 18052 18702 18104 18708
rect 18156 17678 18184 19654
rect 18144 17672 18196 17678
rect 18144 17614 18196 17620
rect 18248 16590 18276 20402
rect 18328 18896 18380 18902
rect 18328 18838 18380 18844
rect 18340 18766 18368 18838
rect 18328 18760 18380 18766
rect 18328 18702 18380 18708
rect 18340 17678 18368 18702
rect 18328 17672 18380 17678
rect 18328 17614 18380 17620
rect 18340 17134 18368 17614
rect 18328 17128 18380 17134
rect 18328 17070 18380 17076
rect 18236 16584 18288 16590
rect 18236 16526 18288 16532
rect 18052 16448 18104 16454
rect 18052 16390 18104 16396
rect 17960 16108 18012 16114
rect 17960 16050 18012 16056
rect 17972 15434 18000 16050
rect 18064 15502 18092 16390
rect 18248 16250 18276 16526
rect 18236 16244 18288 16250
rect 18236 16186 18288 16192
rect 18052 15496 18104 15502
rect 18052 15438 18104 15444
rect 17960 15428 18012 15434
rect 17960 15370 18012 15376
rect 17972 15162 18000 15370
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 18144 13932 18196 13938
rect 18144 13874 18196 13880
rect 18156 12986 18184 13874
rect 17960 12980 18012 12986
rect 17960 12922 18012 12928
rect 18144 12980 18196 12986
rect 18144 12922 18196 12928
rect 17868 12640 17920 12646
rect 17868 12582 17920 12588
rect 17972 12434 18000 12922
rect 17972 12406 18092 12434
rect 17868 12232 17920 12238
rect 17920 12192 18000 12220
rect 17868 12174 17920 12180
rect 17868 11824 17920 11830
rect 17868 11766 17920 11772
rect 17880 11354 17908 11766
rect 17868 11348 17920 11354
rect 17868 11290 17920 11296
rect 17972 10146 18000 12192
rect 18064 11642 18092 12406
rect 18144 12164 18196 12170
rect 18144 12106 18196 12112
rect 18156 11762 18184 12106
rect 18248 11937 18276 16186
rect 18234 11928 18290 11937
rect 18234 11863 18290 11872
rect 18144 11756 18196 11762
rect 18144 11698 18196 11704
rect 18064 11614 18184 11642
rect 18052 11076 18104 11082
rect 18052 11018 18104 11024
rect 18064 10266 18092 11018
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 17972 10118 18092 10146
rect 18064 9654 18092 10118
rect 18052 9648 18104 9654
rect 17958 9616 18014 9625
rect 17880 9586 17958 9602
rect 17868 9580 17958 9586
rect 17920 9574 17958 9580
rect 18052 9590 18104 9596
rect 17958 9551 18014 9560
rect 17868 9522 17920 9528
rect 18064 9466 18092 9590
rect 17972 9438 18092 9466
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 17684 9172 17736 9178
rect 17684 9114 17736 9120
rect 17774 9072 17830 9081
rect 17774 9007 17830 9016
rect 17788 8974 17816 9007
rect 17776 8968 17828 8974
rect 17776 8910 17828 8916
rect 17972 8906 18000 9438
rect 18156 8974 18184 11614
rect 18432 11354 18460 26726
rect 19076 26246 19104 27066
rect 18696 26240 18748 26246
rect 18696 26182 18748 26188
rect 19064 26240 19116 26246
rect 19064 26182 19116 26188
rect 18708 25906 18736 26182
rect 18696 25900 18748 25906
rect 18696 25842 18748 25848
rect 18880 25900 18932 25906
rect 18880 25842 18932 25848
rect 18892 25498 18920 25842
rect 18880 25492 18932 25498
rect 18880 25434 18932 25440
rect 18604 25288 18656 25294
rect 18604 25230 18656 25236
rect 18616 24886 18644 25230
rect 18604 24880 18656 24886
rect 18604 24822 18656 24828
rect 18616 23866 18644 24822
rect 18604 23860 18656 23866
rect 18604 23802 18656 23808
rect 18880 22636 18932 22642
rect 18880 22578 18932 22584
rect 19064 22636 19116 22642
rect 19064 22578 19116 22584
rect 18512 22432 18564 22438
rect 18512 22374 18564 22380
rect 18524 22030 18552 22374
rect 18512 22024 18564 22030
rect 18512 21966 18564 21972
rect 18892 21894 18920 22578
rect 19076 22234 19104 22578
rect 19064 22228 19116 22234
rect 19064 22170 19116 22176
rect 19168 22094 19196 29446
rect 19260 29306 19288 29582
rect 19614 29543 19616 29552
rect 19668 29543 19670 29552
rect 19616 29514 19668 29520
rect 19432 29504 19484 29510
rect 19432 29446 19484 29452
rect 19248 29300 19300 29306
rect 19248 29242 19300 29248
rect 19444 29170 19472 29446
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19432 29164 19484 29170
rect 19432 29106 19484 29112
rect 19340 28552 19392 28558
rect 19340 28494 19392 28500
rect 19352 28014 19380 28494
rect 19432 28416 19484 28422
rect 19432 28358 19484 28364
rect 19444 28082 19472 28358
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19432 28076 19484 28082
rect 19432 28018 19484 28024
rect 19340 28008 19392 28014
rect 19340 27950 19392 27956
rect 19892 27872 19944 27878
rect 19892 27814 19944 27820
rect 19904 27674 19932 27814
rect 19892 27668 19944 27674
rect 19892 27610 19944 27616
rect 19340 27532 19392 27538
rect 19340 27474 19392 27480
rect 19352 26994 19380 27474
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19996 26994 20024 30110
rect 20996 30048 21048 30054
rect 20996 29990 21048 29996
rect 20260 29504 20312 29510
rect 20260 29446 20312 29452
rect 20168 29028 20220 29034
rect 20168 28970 20220 28976
rect 20076 28076 20128 28082
rect 20076 28018 20128 28024
rect 20088 27946 20116 28018
rect 20076 27940 20128 27946
rect 20076 27882 20128 27888
rect 19340 26988 19392 26994
rect 19340 26930 19392 26936
rect 19984 26988 20036 26994
rect 19984 26930 20036 26936
rect 19248 26852 19300 26858
rect 19248 26794 19300 26800
rect 19260 26382 19288 26794
rect 19352 26450 19380 26930
rect 19340 26444 19392 26450
rect 19340 26386 19392 26392
rect 19248 26376 19300 26382
rect 19248 26318 19300 26324
rect 19260 25430 19288 26318
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19708 25696 19760 25702
rect 19708 25638 19760 25644
rect 19248 25424 19300 25430
rect 19248 25366 19300 25372
rect 19720 25294 19748 25638
rect 19432 25288 19484 25294
rect 19432 25230 19484 25236
rect 19708 25288 19760 25294
rect 19708 25230 19760 25236
rect 19340 24200 19392 24206
rect 19340 24142 19392 24148
rect 19352 23662 19380 24142
rect 19340 23656 19392 23662
rect 19340 23598 19392 23604
rect 19248 23588 19300 23594
rect 19248 23530 19300 23536
rect 19076 22066 19196 22094
rect 18880 21888 18932 21894
rect 18880 21830 18932 21836
rect 18880 21344 18932 21350
rect 18880 21286 18932 21292
rect 18892 20874 18920 21286
rect 18880 20868 18932 20874
rect 18880 20810 18932 20816
rect 18696 18828 18748 18834
rect 18696 18770 18748 18776
rect 18708 18290 18736 18770
rect 18696 18284 18748 18290
rect 18696 18226 18748 18232
rect 18708 17678 18736 18226
rect 18696 17672 18748 17678
rect 18748 17620 18828 17626
rect 18696 17614 18828 17620
rect 18708 17598 18828 17614
rect 18696 17536 18748 17542
rect 18696 17478 18748 17484
rect 18708 16114 18736 17478
rect 18800 17270 18828 17598
rect 18788 17264 18840 17270
rect 18788 17206 18840 17212
rect 18892 17202 18920 20810
rect 18972 20256 19024 20262
rect 18970 20224 18972 20233
rect 19024 20224 19026 20233
rect 18970 20159 19026 20168
rect 18970 19408 19026 19417
rect 18970 19343 18972 19352
rect 19024 19343 19026 19352
rect 18972 19314 19024 19320
rect 18972 17536 19024 17542
rect 18972 17478 19024 17484
rect 18880 17196 18932 17202
rect 18880 17138 18932 17144
rect 18696 16108 18748 16114
rect 18696 16050 18748 16056
rect 18984 15094 19012 17478
rect 19076 15745 19104 22066
rect 19156 20936 19208 20942
rect 19156 20878 19208 20884
rect 19168 20398 19196 20878
rect 19156 20392 19208 20398
rect 19156 20334 19208 20340
rect 19168 19922 19196 20334
rect 19156 19916 19208 19922
rect 19156 19858 19208 19864
rect 19156 19780 19208 19786
rect 19156 19722 19208 19728
rect 19168 19378 19196 19722
rect 19156 19372 19208 19378
rect 19156 19314 19208 19320
rect 19168 18902 19196 19314
rect 19156 18896 19208 18902
rect 19156 18838 19208 18844
rect 19260 17796 19288 23530
rect 19352 23361 19380 23598
rect 19338 23352 19394 23361
rect 19338 23287 19394 23296
rect 19340 23180 19392 23186
rect 19340 23122 19392 23128
rect 19352 22710 19380 23122
rect 19444 23118 19472 25230
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19708 24812 19760 24818
rect 19708 24754 19760 24760
rect 19720 24410 19748 24754
rect 19708 24404 19760 24410
rect 19708 24346 19760 24352
rect 19996 24206 20024 26930
rect 19984 24200 20036 24206
rect 19984 24142 20036 24148
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19616 23656 19668 23662
rect 19616 23598 19668 23604
rect 19628 23118 19656 23598
rect 19432 23112 19484 23118
rect 19432 23054 19484 23060
rect 19616 23112 19668 23118
rect 19616 23054 19668 23060
rect 19340 22704 19392 22710
rect 19340 22646 19392 22652
rect 19444 22642 19472 23054
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19432 22636 19484 22642
rect 19432 22578 19484 22584
rect 19996 22506 20024 24142
rect 20076 23112 20128 23118
rect 20076 23054 20128 23060
rect 19984 22500 20036 22506
rect 19984 22442 20036 22448
rect 20088 22438 20116 23054
rect 20076 22432 20128 22438
rect 20076 22374 20128 22380
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 20088 21554 20116 22374
rect 19800 21548 19852 21554
rect 19800 21490 19852 21496
rect 20076 21548 20128 21554
rect 20076 21490 20128 21496
rect 19812 21146 19840 21490
rect 20076 21412 20128 21418
rect 20076 21354 20128 21360
rect 19800 21140 19852 21146
rect 19800 21082 19852 21088
rect 19984 21072 20036 21078
rect 19984 21014 20036 21020
rect 19616 20936 19668 20942
rect 19444 20896 19616 20924
rect 19340 20392 19392 20398
rect 19340 20334 19392 20340
rect 19352 18766 19380 20334
rect 19444 20262 19472 20896
rect 19616 20878 19668 20884
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19798 20360 19854 20369
rect 19798 20295 19854 20304
rect 19432 20256 19484 20262
rect 19432 20198 19484 20204
rect 19522 20088 19578 20097
rect 19522 20023 19578 20032
rect 19536 19854 19564 20023
rect 19812 19854 19840 20295
rect 19892 20256 19944 20262
rect 19892 20198 19944 20204
rect 19904 19990 19932 20198
rect 19892 19984 19944 19990
rect 19892 19926 19944 19932
rect 19432 19848 19484 19854
rect 19432 19790 19484 19796
rect 19524 19848 19576 19854
rect 19524 19790 19576 19796
rect 19800 19848 19852 19854
rect 19800 19790 19852 19796
rect 19444 19378 19472 19790
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 19444 18834 19472 19314
rect 19432 18828 19484 18834
rect 19432 18770 19484 18776
rect 19996 18766 20024 21014
rect 20088 21010 20116 21354
rect 20076 21004 20128 21010
rect 20076 20946 20128 20952
rect 20088 20602 20116 20946
rect 20076 20596 20128 20602
rect 20076 20538 20128 20544
rect 20088 19786 20116 20538
rect 20076 19780 20128 19786
rect 20076 19722 20128 19728
rect 19340 18760 19392 18766
rect 19340 18702 19392 18708
rect 19984 18760 20036 18766
rect 19984 18702 20036 18708
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 20076 18284 20128 18290
rect 20076 18226 20128 18232
rect 19432 18148 19484 18154
rect 19432 18090 19484 18096
rect 19260 17768 19380 17796
rect 19062 15736 19118 15745
rect 19062 15671 19118 15680
rect 18972 15088 19024 15094
rect 18972 15030 19024 15036
rect 18788 14272 18840 14278
rect 18788 14214 18840 14220
rect 18696 13252 18748 13258
rect 18696 13194 18748 13200
rect 18708 12850 18736 13194
rect 18512 12844 18564 12850
rect 18512 12786 18564 12792
rect 18696 12844 18748 12850
rect 18696 12786 18748 12792
rect 18524 12442 18552 12786
rect 18512 12436 18564 12442
rect 18512 12378 18564 12384
rect 18512 11552 18564 11558
rect 18512 11494 18564 11500
rect 18420 11348 18472 11354
rect 18420 11290 18472 11296
rect 18236 11008 18288 11014
rect 18236 10950 18288 10956
rect 18248 10198 18276 10950
rect 18432 10810 18460 11290
rect 18420 10804 18472 10810
rect 18420 10746 18472 10752
rect 18326 10296 18382 10305
rect 18326 10231 18382 10240
rect 18236 10192 18288 10198
rect 18236 10134 18288 10140
rect 18340 10062 18368 10231
rect 18524 10062 18552 11494
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18512 10056 18564 10062
rect 18512 9998 18564 10004
rect 18340 9450 18368 9998
rect 18800 9722 18828 14214
rect 19352 13530 19380 17768
rect 19444 17610 19472 18090
rect 19984 18080 20036 18086
rect 19984 18022 20036 18028
rect 19432 17604 19484 17610
rect 19432 17546 19484 17552
rect 19444 16726 19472 17546
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19432 16720 19484 16726
rect 19432 16662 19484 16668
rect 19616 16720 19668 16726
rect 19616 16662 19668 16668
rect 19628 16590 19656 16662
rect 19616 16584 19668 16590
rect 19616 16526 19668 16532
rect 19432 16516 19484 16522
rect 19432 16458 19484 16464
rect 19444 16182 19472 16458
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19432 16176 19484 16182
rect 19432 16118 19484 16124
rect 19800 16176 19852 16182
rect 19800 16118 19852 16124
rect 19708 16108 19760 16114
rect 19708 16050 19760 16056
rect 19432 15972 19484 15978
rect 19432 15914 19484 15920
rect 19444 15502 19472 15914
rect 19720 15706 19748 16050
rect 19812 15706 19840 16118
rect 19708 15700 19760 15706
rect 19708 15642 19760 15648
rect 19800 15700 19852 15706
rect 19800 15642 19852 15648
rect 19812 15570 19840 15642
rect 19800 15564 19852 15570
rect 19800 15506 19852 15512
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19996 14056 20024 18022
rect 20088 17678 20116 18226
rect 20076 17672 20128 17678
rect 20076 17614 20128 17620
rect 20088 17202 20116 17614
rect 20076 17196 20128 17202
rect 20076 17138 20128 17144
rect 20088 16114 20116 17138
rect 20076 16108 20128 16114
rect 20076 16050 20128 16056
rect 20088 15502 20116 16050
rect 20076 15496 20128 15502
rect 20076 15438 20128 15444
rect 20076 15360 20128 15366
rect 20076 15302 20128 15308
rect 19904 14028 20024 14056
rect 19432 13728 19484 13734
rect 19432 13670 19484 13676
rect 19340 13524 19392 13530
rect 19340 13466 19392 13472
rect 19340 13388 19392 13394
rect 19340 13330 19392 13336
rect 19156 13184 19208 13190
rect 19352 13138 19380 13330
rect 19156 13126 19208 13132
rect 19064 12776 19116 12782
rect 19064 12718 19116 12724
rect 19076 12434 19104 12718
rect 18984 12406 19104 12434
rect 18984 12102 19012 12406
rect 18972 12096 19024 12102
rect 18972 12038 19024 12044
rect 18984 11694 19012 12038
rect 18880 11688 18932 11694
rect 18880 11630 18932 11636
rect 18972 11688 19024 11694
rect 18972 11630 19024 11636
rect 18788 9716 18840 9722
rect 18788 9658 18840 9664
rect 18420 9580 18472 9586
rect 18420 9522 18472 9528
rect 18432 9489 18460 9522
rect 18418 9480 18474 9489
rect 18328 9444 18380 9450
rect 18418 9415 18474 9424
rect 18328 9386 18380 9392
rect 18144 8968 18196 8974
rect 18144 8910 18196 8916
rect 18420 8968 18472 8974
rect 18420 8910 18472 8916
rect 17960 8900 18012 8906
rect 17960 8842 18012 8848
rect 17500 8832 17552 8838
rect 17500 8774 17552 8780
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17420 7886 17448 8230
rect 17512 8090 17540 8774
rect 17500 8084 17552 8090
rect 17500 8026 17552 8032
rect 17868 8016 17920 8022
rect 17868 7958 17920 7964
rect 17408 7880 17460 7886
rect 17408 7822 17460 7828
rect 17316 5704 17368 5710
rect 17316 5646 17368 5652
rect 17316 5568 17368 5574
rect 17316 5510 17368 5516
rect 17328 5234 17356 5510
rect 17316 5228 17368 5234
rect 17316 5170 17368 5176
rect 17144 5086 17264 5114
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 17144 2961 17172 5086
rect 17222 4992 17278 5001
rect 17222 4927 17278 4936
rect 17130 2952 17186 2961
rect 17130 2887 17186 2896
rect 16776 2746 16988 2774
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 16776 2145 16804 2246
rect 16762 2136 16818 2145
rect 16762 2071 16818 2080
rect 16776 2038 16804 2071
rect 16764 2032 16816 2038
rect 16764 1974 16816 1980
rect 16672 1896 16724 1902
rect 16672 1838 16724 1844
rect 16684 800 16712 1838
rect 16960 800 16988 2746
rect 17236 800 17264 4927
rect 17420 3534 17448 7822
rect 17500 7200 17552 7206
rect 17500 7142 17552 7148
rect 17408 3528 17460 3534
rect 17408 3470 17460 3476
rect 17512 800 17540 7142
rect 17684 6248 17736 6254
rect 17684 6190 17736 6196
rect 17592 5772 17644 5778
rect 17592 5714 17644 5720
rect 17604 5234 17632 5714
rect 17696 5710 17724 6190
rect 17880 5914 17908 7958
rect 17868 5908 17920 5914
rect 17868 5850 17920 5856
rect 17776 5840 17828 5846
rect 17776 5782 17828 5788
rect 17684 5704 17736 5710
rect 17684 5646 17736 5652
rect 17592 5228 17644 5234
rect 17592 5170 17644 5176
rect 17682 4856 17738 4865
rect 17682 4791 17738 4800
rect 17592 3052 17644 3058
rect 17592 2994 17644 3000
rect 17604 2825 17632 2994
rect 17590 2816 17646 2825
rect 17590 2751 17646 2760
rect 17604 2582 17632 2751
rect 17592 2576 17644 2582
rect 17592 2518 17644 2524
rect 17592 2372 17644 2378
rect 17592 2314 17644 2320
rect 17604 1426 17632 2314
rect 17592 1420 17644 1426
rect 17592 1362 17644 1368
rect 17696 898 17724 4791
rect 17788 4146 17816 5782
rect 17868 5024 17920 5030
rect 17868 4966 17920 4972
rect 17776 4140 17828 4146
rect 17776 4082 17828 4088
rect 17880 3890 17908 4966
rect 17972 4826 18000 8842
rect 18052 8492 18104 8498
rect 18052 8434 18104 8440
rect 18064 8090 18092 8434
rect 18432 8242 18460 8910
rect 18432 8214 18644 8242
rect 18052 8084 18104 8090
rect 18052 8026 18104 8032
rect 18328 7880 18380 7886
rect 18328 7822 18380 7828
rect 18052 6452 18104 6458
rect 18052 6394 18104 6400
rect 17960 4820 18012 4826
rect 17960 4762 18012 4768
rect 17960 4684 18012 4690
rect 17960 4626 18012 4632
rect 17972 4214 18000 4626
rect 18064 4554 18092 6394
rect 18236 5364 18288 5370
rect 18236 5306 18288 5312
rect 18144 5092 18196 5098
rect 18144 5034 18196 5040
rect 18156 4758 18184 5034
rect 18248 4826 18276 5306
rect 18236 4820 18288 4826
rect 18236 4762 18288 4768
rect 18144 4752 18196 4758
rect 18144 4694 18196 4700
rect 18052 4548 18104 4554
rect 18052 4490 18104 4496
rect 17960 4208 18012 4214
rect 17960 4150 18012 4156
rect 18064 4146 18092 4490
rect 18236 4480 18288 4486
rect 18236 4422 18288 4428
rect 18248 4282 18276 4422
rect 18144 4276 18196 4282
rect 18144 4218 18196 4224
rect 18236 4276 18288 4282
rect 18236 4218 18288 4224
rect 18052 4140 18104 4146
rect 18052 4082 18104 4088
rect 17880 3862 18092 3890
rect 17960 3664 18012 3670
rect 17960 3606 18012 3612
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 17880 3126 17908 3470
rect 17868 3120 17920 3126
rect 17868 3062 17920 3068
rect 17774 2952 17830 2961
rect 17774 2887 17830 2896
rect 17788 2854 17816 2887
rect 17776 2848 17828 2854
rect 17776 2790 17828 2796
rect 17972 2650 18000 3606
rect 17960 2644 18012 2650
rect 17960 2586 18012 2592
rect 17696 870 17816 898
rect 17788 800 17816 870
rect 18064 800 18092 3862
rect 18156 2446 18184 4218
rect 18144 2440 18196 2446
rect 18144 2382 18196 2388
rect 18340 800 18368 7822
rect 18512 7744 18564 7750
rect 18512 7686 18564 7692
rect 18524 7410 18552 7686
rect 18512 7404 18564 7410
rect 18512 7346 18564 7352
rect 18420 7336 18472 7342
rect 18420 7278 18472 7284
rect 18432 3466 18460 7278
rect 18512 6792 18564 6798
rect 18616 6780 18644 8214
rect 18564 6752 18644 6780
rect 18512 6734 18564 6740
rect 18512 5160 18564 5166
rect 18512 5102 18564 5108
rect 18524 4078 18552 5102
rect 18616 4282 18644 6752
rect 18892 5914 18920 11630
rect 18880 5908 18932 5914
rect 18880 5850 18932 5856
rect 18788 5228 18840 5234
rect 18788 5170 18840 5176
rect 18696 4752 18748 4758
rect 18696 4694 18748 4700
rect 18604 4276 18656 4282
rect 18604 4218 18656 4224
rect 18708 4146 18736 4694
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 18512 4072 18564 4078
rect 18512 4014 18564 4020
rect 18604 4072 18656 4078
rect 18604 4014 18656 4020
rect 18420 3460 18472 3466
rect 18420 3402 18472 3408
rect 18616 800 18644 4014
rect 18696 4004 18748 4010
rect 18696 3946 18748 3952
rect 18708 2990 18736 3946
rect 18696 2984 18748 2990
rect 18696 2926 18748 2932
rect 18800 2310 18828 5170
rect 18892 4486 18920 5850
rect 18880 4480 18932 4486
rect 18880 4422 18932 4428
rect 18892 3754 18920 4422
rect 18984 4010 19012 11630
rect 19168 6322 19196 13126
rect 19260 13110 19380 13138
rect 19260 12986 19288 13110
rect 19444 13002 19472 13670
rect 19904 13394 19932 14028
rect 19984 13932 20036 13938
rect 19984 13874 20036 13880
rect 19892 13388 19944 13394
rect 19892 13330 19944 13336
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19248 12980 19300 12986
rect 19248 12922 19300 12928
rect 19352 12974 19472 13002
rect 19352 12238 19380 12974
rect 19524 12912 19576 12918
rect 19892 12912 19944 12918
rect 19524 12854 19576 12860
rect 19798 12880 19854 12889
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 19340 12232 19392 12238
rect 19340 12174 19392 12180
rect 19340 12096 19392 12102
rect 19340 12038 19392 12044
rect 19248 11076 19300 11082
rect 19248 11018 19300 11024
rect 19260 10810 19288 11018
rect 19248 10804 19300 10810
rect 19248 10746 19300 10752
rect 19352 9994 19380 12038
rect 19444 11150 19472 12786
rect 19536 12102 19564 12854
rect 19892 12854 19944 12860
rect 19798 12815 19800 12824
rect 19852 12815 19854 12824
rect 19800 12786 19852 12792
rect 19800 12436 19852 12442
rect 19904 12434 19932 12854
rect 19852 12406 19932 12434
rect 19800 12378 19852 12384
rect 19812 12238 19840 12378
rect 19800 12232 19852 12238
rect 19800 12174 19852 12180
rect 19524 12096 19576 12102
rect 19524 12038 19576 12044
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19708 11824 19760 11830
rect 19706 11792 19708 11801
rect 19800 11824 19852 11830
rect 19760 11792 19762 11801
rect 19800 11766 19852 11772
rect 19706 11727 19762 11736
rect 19706 11384 19762 11393
rect 19812 11354 19840 11766
rect 19892 11756 19944 11762
rect 19996 11744 20024 13874
rect 20088 13326 20116 15302
rect 20180 14618 20208 28970
rect 20272 22094 20300 29446
rect 20628 28552 20680 28558
rect 20628 28494 20680 28500
rect 20352 28212 20404 28218
rect 20352 28154 20404 28160
rect 20364 27538 20392 28154
rect 20536 27940 20588 27946
rect 20536 27882 20588 27888
rect 20352 27532 20404 27538
rect 20352 27474 20404 27480
rect 20352 26988 20404 26994
rect 20352 26930 20404 26936
rect 20364 26518 20392 26930
rect 20352 26512 20404 26518
rect 20352 26454 20404 26460
rect 20352 26376 20404 26382
rect 20352 26318 20404 26324
rect 20364 25974 20392 26318
rect 20352 25968 20404 25974
rect 20352 25910 20404 25916
rect 20364 25362 20392 25910
rect 20548 25906 20576 27882
rect 20640 26042 20668 28494
rect 20720 28484 20772 28490
rect 20720 28426 20772 28432
rect 20732 28218 20760 28426
rect 20720 28212 20772 28218
rect 20720 28154 20772 28160
rect 21008 28150 21036 29990
rect 21376 29714 21404 30534
rect 21836 30326 21864 31962
rect 22376 31816 22428 31822
rect 22376 31758 22428 31764
rect 22192 31748 22244 31754
rect 22192 31690 22244 31696
rect 22204 31210 22232 31690
rect 22388 31346 22416 31758
rect 22284 31340 22336 31346
rect 22284 31282 22336 31288
rect 22376 31340 22428 31346
rect 22376 31282 22428 31288
rect 22192 31204 22244 31210
rect 22192 31146 22244 31152
rect 21824 30320 21876 30326
rect 21824 30262 21876 30268
rect 21456 30184 21508 30190
rect 21456 30126 21508 30132
rect 21364 29708 21416 29714
rect 21364 29650 21416 29656
rect 21468 28626 21496 30126
rect 21456 28620 21508 28626
rect 21456 28562 21508 28568
rect 20996 28144 21048 28150
rect 20996 28086 21048 28092
rect 21008 27674 21036 28086
rect 21836 28082 21864 30262
rect 22008 30116 22060 30122
rect 22008 30058 22060 30064
rect 22020 29238 22048 30058
rect 22100 30048 22152 30054
rect 22100 29990 22152 29996
rect 22112 29782 22140 29990
rect 22204 29782 22232 31146
rect 22100 29776 22152 29782
rect 22100 29718 22152 29724
rect 22192 29776 22244 29782
rect 22192 29718 22244 29724
rect 22008 29232 22060 29238
rect 22008 29174 22060 29180
rect 22008 28416 22060 28422
rect 22008 28358 22060 28364
rect 21824 28076 21876 28082
rect 21824 28018 21876 28024
rect 21272 28008 21324 28014
rect 21272 27950 21324 27956
rect 21284 27878 21312 27950
rect 21272 27872 21324 27878
rect 21272 27814 21324 27820
rect 20996 27668 21048 27674
rect 20996 27610 21048 27616
rect 21836 27470 21864 28018
rect 22020 27606 22048 28358
rect 22204 28150 22232 29718
rect 22296 29628 22324 31282
rect 22480 30734 22508 32166
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 65654 32124 65962 32133
rect 65654 32122 65660 32124
rect 65716 32122 65740 32124
rect 65796 32122 65820 32124
rect 65876 32122 65900 32124
rect 65956 32122 65962 32124
rect 65716 32070 65718 32122
rect 65898 32070 65900 32122
rect 65654 32068 65660 32070
rect 65716 32068 65740 32070
rect 65796 32068 65820 32070
rect 65876 32068 65900 32070
rect 65956 32068 65962 32070
rect 65654 32059 65962 32068
rect 67652 32065 67680 32166
rect 67638 32056 67694 32065
rect 67638 31991 67694 32000
rect 23296 31816 23348 31822
rect 23296 31758 23348 31764
rect 22468 30728 22520 30734
rect 22468 30670 22520 30676
rect 23308 30394 23336 31758
rect 23572 31748 23624 31754
rect 23572 31690 23624 31696
rect 23388 31680 23440 31686
rect 23388 31622 23440 31628
rect 23400 31278 23428 31622
rect 23480 31340 23532 31346
rect 23480 31282 23532 31288
rect 23388 31272 23440 31278
rect 23388 31214 23440 31220
rect 23296 30388 23348 30394
rect 23296 30330 23348 30336
rect 22560 30252 22612 30258
rect 22560 30194 22612 30200
rect 22572 29850 22600 30194
rect 22560 29844 22612 29850
rect 22560 29786 22612 29792
rect 22376 29640 22428 29646
rect 22296 29600 22376 29628
rect 22192 28144 22244 28150
rect 22192 28086 22244 28092
rect 22008 27600 22060 27606
rect 22008 27542 22060 27548
rect 22204 27538 22232 28086
rect 22192 27532 22244 27538
rect 22192 27474 22244 27480
rect 21824 27464 21876 27470
rect 21824 27406 21876 27412
rect 21836 27130 21864 27406
rect 21824 27124 21876 27130
rect 21824 27066 21876 27072
rect 22008 26852 22060 26858
rect 22008 26794 22060 26800
rect 20628 26036 20680 26042
rect 20628 25978 20680 25984
rect 20536 25900 20588 25906
rect 20536 25842 20588 25848
rect 20548 25430 20576 25842
rect 20536 25424 20588 25430
rect 20536 25366 20588 25372
rect 20352 25356 20404 25362
rect 20352 25298 20404 25304
rect 20364 24138 20392 25298
rect 20536 25288 20588 25294
rect 20536 25230 20588 25236
rect 20548 24614 20576 25230
rect 20640 24818 20668 25978
rect 22020 25906 22048 26794
rect 22008 25900 22060 25906
rect 22008 25842 22060 25848
rect 22192 25900 22244 25906
rect 22192 25842 22244 25848
rect 21732 25696 21784 25702
rect 21732 25638 21784 25644
rect 20628 24812 20680 24818
rect 20628 24754 20680 24760
rect 20536 24608 20588 24614
rect 20536 24550 20588 24556
rect 20352 24132 20404 24138
rect 20352 24074 20404 24080
rect 20364 23186 20392 24074
rect 20444 23860 20496 23866
rect 20444 23802 20496 23808
rect 20352 23180 20404 23186
rect 20352 23122 20404 23128
rect 20272 22066 20392 22094
rect 20260 22024 20312 22030
rect 20260 21966 20312 21972
rect 20272 20806 20300 21966
rect 20260 20800 20312 20806
rect 20260 20742 20312 20748
rect 20260 19848 20312 19854
rect 20260 19790 20312 19796
rect 20272 19514 20300 19790
rect 20260 19508 20312 19514
rect 20260 19450 20312 19456
rect 20260 18828 20312 18834
rect 20260 18770 20312 18776
rect 20272 16046 20300 18770
rect 20260 16040 20312 16046
rect 20260 15982 20312 15988
rect 20272 15484 20300 15982
rect 20364 15978 20392 22066
rect 20456 21078 20484 23802
rect 20548 22094 20576 24550
rect 20640 23118 20668 24754
rect 20628 23112 20680 23118
rect 20628 23054 20680 23060
rect 21640 22568 21692 22574
rect 21640 22510 21692 22516
rect 21652 22098 21680 22510
rect 20548 22066 20668 22094
rect 20444 21072 20496 21078
rect 20444 21014 20496 21020
rect 20640 21010 20668 22066
rect 21640 22092 21692 22098
rect 21640 22034 21692 22040
rect 21088 21548 21140 21554
rect 21088 21490 21140 21496
rect 20720 21480 20772 21486
rect 20720 21422 20772 21428
rect 20628 21004 20680 21010
rect 20628 20946 20680 20952
rect 20628 20868 20680 20874
rect 20628 20810 20680 20816
rect 20444 19848 20496 19854
rect 20444 19790 20496 19796
rect 20456 19310 20484 19790
rect 20536 19712 20588 19718
rect 20536 19654 20588 19660
rect 20548 19378 20576 19654
rect 20640 19446 20668 20810
rect 20732 20806 20760 21422
rect 21100 21078 21128 21490
rect 21744 21146 21772 25638
rect 22204 24954 22232 25842
rect 22192 24948 22244 24954
rect 22192 24890 22244 24896
rect 22296 24818 22324 29600
rect 22376 29582 22428 29588
rect 23492 29510 23520 31282
rect 23584 31260 23612 31690
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 23584 31232 23704 31260
rect 23480 29504 23532 29510
rect 23480 29446 23532 29452
rect 22560 28484 22612 28490
rect 22560 28426 22612 28432
rect 22572 28218 22600 28426
rect 22560 28212 22612 28218
rect 22560 28154 22612 28160
rect 22468 28076 22520 28082
rect 22468 28018 22520 28024
rect 22480 27538 22508 28018
rect 22560 28008 22612 28014
rect 22560 27950 22612 27956
rect 22572 27878 22600 27950
rect 22560 27872 22612 27878
rect 22560 27814 22612 27820
rect 23572 27872 23624 27878
rect 23572 27814 23624 27820
rect 22468 27532 22520 27538
rect 22468 27474 22520 27480
rect 23584 27470 23612 27814
rect 23204 27464 23256 27470
rect 23202 27432 23204 27441
rect 23572 27464 23624 27470
rect 23256 27432 23258 27441
rect 23572 27406 23624 27412
rect 23202 27367 23258 27376
rect 23480 27328 23532 27334
rect 23480 27270 23532 27276
rect 23492 27130 23520 27270
rect 23480 27124 23532 27130
rect 23480 27066 23532 27072
rect 22560 27056 22612 27062
rect 22560 26998 22612 27004
rect 22468 26308 22520 26314
rect 22468 26250 22520 26256
rect 22480 26042 22508 26250
rect 22468 26036 22520 26042
rect 22468 25978 22520 25984
rect 22284 24812 22336 24818
rect 22284 24754 22336 24760
rect 21824 24608 21876 24614
rect 21824 24550 21876 24556
rect 21836 24070 21864 24550
rect 22296 24342 22324 24754
rect 22284 24336 22336 24342
rect 22284 24278 22336 24284
rect 22376 24200 22428 24206
rect 21928 24138 22232 24154
rect 22376 24142 22428 24148
rect 21916 24132 22232 24138
rect 21968 24126 22232 24132
rect 21916 24074 21968 24080
rect 21824 24064 21876 24070
rect 21824 24006 21876 24012
rect 21836 23730 21864 24006
rect 21916 23792 21968 23798
rect 21916 23734 21968 23740
rect 21824 23724 21876 23730
rect 21824 23666 21876 23672
rect 21928 23322 21956 23734
rect 22100 23520 22152 23526
rect 22100 23462 22152 23468
rect 21916 23316 21968 23322
rect 21916 23258 21968 23264
rect 21916 22024 21968 22030
rect 21914 21992 21916 22001
rect 21968 21992 21970 22001
rect 21914 21927 21970 21936
rect 21732 21140 21784 21146
rect 21732 21082 21784 21088
rect 21088 21072 21140 21078
rect 21088 21014 21140 21020
rect 20720 20800 20772 20806
rect 20720 20742 20772 20748
rect 20732 20602 20760 20742
rect 20720 20596 20772 20602
rect 20720 20538 20772 20544
rect 21100 20466 21128 21014
rect 21548 20868 21600 20874
rect 21548 20810 21600 20816
rect 21088 20460 21140 20466
rect 21088 20402 21140 20408
rect 21272 20392 21324 20398
rect 21272 20334 21324 20340
rect 20720 20324 20772 20330
rect 20720 20266 20772 20272
rect 20628 19440 20680 19446
rect 20628 19382 20680 19388
rect 20536 19372 20588 19378
rect 20536 19314 20588 19320
rect 20444 19304 20496 19310
rect 20444 19246 20496 19252
rect 20628 19168 20680 19174
rect 20628 19110 20680 19116
rect 20444 18760 20496 18766
rect 20444 18702 20496 18708
rect 20456 16726 20484 18702
rect 20640 18290 20668 19110
rect 20732 18970 20760 20266
rect 21284 19854 21312 20334
rect 21560 20262 21588 20810
rect 21548 20256 21600 20262
rect 21548 20198 21600 20204
rect 21822 20224 21878 20233
rect 21180 19848 21232 19854
rect 21180 19790 21232 19796
rect 21272 19848 21324 19854
rect 21272 19790 21324 19796
rect 21192 19310 21220 19790
rect 21180 19304 21232 19310
rect 21178 19272 21180 19281
rect 21364 19304 21416 19310
rect 21232 19272 21234 19281
rect 21364 19246 21416 19252
rect 21178 19207 21234 19216
rect 20720 18964 20772 18970
rect 20720 18906 20772 18912
rect 21192 18766 21220 19207
rect 21272 18964 21324 18970
rect 21272 18906 21324 18912
rect 21180 18760 21232 18766
rect 21180 18702 21232 18708
rect 20812 18624 20864 18630
rect 20812 18566 20864 18572
rect 20904 18624 20956 18630
rect 20904 18566 20956 18572
rect 20536 18284 20588 18290
rect 20536 18226 20588 18232
rect 20628 18284 20680 18290
rect 20628 18226 20680 18232
rect 20548 18057 20576 18226
rect 20720 18148 20772 18154
rect 20720 18090 20772 18096
rect 20534 18048 20590 18057
rect 20534 17983 20590 17992
rect 20536 17876 20588 17882
rect 20536 17818 20588 17824
rect 20444 16720 20496 16726
rect 20444 16662 20496 16668
rect 20352 15972 20404 15978
rect 20352 15914 20404 15920
rect 20444 15904 20496 15910
rect 20444 15846 20496 15852
rect 20352 15496 20404 15502
rect 20272 15456 20352 15484
rect 20352 15438 20404 15444
rect 20168 14612 20220 14618
rect 20168 14554 20220 14560
rect 20168 14408 20220 14414
rect 20168 14350 20220 14356
rect 20180 14074 20208 14350
rect 20168 14068 20220 14074
rect 20168 14010 20220 14016
rect 20168 13932 20220 13938
rect 20168 13874 20220 13880
rect 20076 13320 20128 13326
rect 20076 13262 20128 13268
rect 20180 12986 20208 13874
rect 20260 13728 20312 13734
rect 20260 13670 20312 13676
rect 20168 12980 20220 12986
rect 20168 12922 20220 12928
rect 20272 12918 20300 13670
rect 20260 12912 20312 12918
rect 20166 12880 20222 12889
rect 20260 12854 20312 12860
rect 20166 12815 20222 12824
rect 20076 12096 20128 12102
rect 20076 12038 20128 12044
rect 19944 11716 20024 11744
rect 19892 11698 19944 11704
rect 19706 11319 19762 11328
rect 19800 11348 19852 11354
rect 19614 11248 19670 11257
rect 19614 11183 19616 11192
rect 19668 11183 19670 11192
rect 19720 11200 19748 11319
rect 19800 11290 19852 11296
rect 19904 11286 19932 11698
rect 20088 11393 20116 12038
rect 20180 11558 20208 12815
rect 20260 12436 20312 12442
rect 20260 12378 20312 12384
rect 20272 12322 20300 12378
rect 20272 12294 20392 12322
rect 20260 12232 20312 12238
rect 20260 12174 20312 12180
rect 20272 11801 20300 12174
rect 20258 11792 20314 11801
rect 20258 11727 20314 11736
rect 20168 11552 20220 11558
rect 20220 11512 20300 11540
rect 20168 11494 20220 11500
rect 20074 11384 20130 11393
rect 20074 11319 20130 11328
rect 19892 11280 19944 11286
rect 20076 11280 20128 11286
rect 19944 11240 20024 11268
rect 19892 11222 19944 11228
rect 19800 11212 19852 11218
rect 19720 11172 19800 11200
rect 19616 11154 19668 11160
rect 19800 11154 19852 11160
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19444 10062 19472 11086
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19800 10736 19852 10742
rect 19800 10678 19852 10684
rect 19524 10192 19576 10198
rect 19524 10134 19576 10140
rect 19706 10160 19762 10169
rect 19432 10056 19484 10062
rect 19432 9998 19484 10004
rect 19340 9988 19392 9994
rect 19340 9930 19392 9936
rect 19536 9908 19564 10134
rect 19706 10095 19708 10104
rect 19760 10095 19762 10104
rect 19708 10066 19760 10072
rect 19812 9926 19840 10678
rect 19996 10674 20024 11240
rect 20076 11222 20128 11228
rect 20168 11280 20220 11286
rect 20168 11222 20220 11228
rect 19984 10668 20036 10674
rect 19984 10610 20036 10616
rect 19444 9880 19564 9908
rect 19800 9920 19852 9926
rect 19340 9716 19392 9722
rect 19444 9704 19472 9880
rect 19800 9862 19852 9868
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19996 9761 20024 10610
rect 20088 9926 20116 11222
rect 20180 10266 20208 11222
rect 20168 10260 20220 10266
rect 20168 10202 20220 10208
rect 20180 10062 20208 10202
rect 20168 10056 20220 10062
rect 20168 9998 20220 10004
rect 20076 9920 20128 9926
rect 20180 9897 20208 9998
rect 20076 9862 20128 9868
rect 20166 9888 20222 9897
rect 19982 9752 20038 9761
rect 19524 9716 19576 9722
rect 19444 9676 19524 9704
rect 19340 9658 19392 9664
rect 20088 9722 20116 9862
rect 20166 9823 20222 9832
rect 19982 9687 20038 9696
rect 20076 9716 20128 9722
rect 19524 9658 19576 9664
rect 19352 8537 19380 9658
rect 19524 9580 19576 9586
rect 19524 9522 19576 9528
rect 19536 9110 19564 9522
rect 19524 9104 19576 9110
rect 19524 9046 19576 9052
rect 19996 9042 20024 9687
rect 20076 9658 20128 9664
rect 20076 9512 20128 9518
rect 20076 9454 20128 9460
rect 20088 9382 20116 9454
rect 20076 9376 20128 9382
rect 20076 9318 20128 9324
rect 19984 9036 20036 9042
rect 19984 8978 20036 8984
rect 19892 8968 19944 8974
rect 19430 8936 19486 8945
rect 19892 8910 19944 8916
rect 19430 8871 19486 8880
rect 19444 8566 19472 8871
rect 19904 8838 19932 8910
rect 19892 8832 19944 8838
rect 19892 8774 19944 8780
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19524 8628 19576 8634
rect 19524 8570 19576 8576
rect 19432 8560 19484 8566
rect 19338 8528 19394 8537
rect 19432 8502 19484 8508
rect 19338 8463 19394 8472
rect 19536 8480 19564 8570
rect 19616 8492 19668 8498
rect 19352 8294 19380 8463
rect 19536 8452 19616 8480
rect 19536 8412 19564 8452
rect 19616 8434 19668 8440
rect 19444 8384 19564 8412
rect 19340 8288 19392 8294
rect 19340 8230 19392 8236
rect 19156 6316 19208 6322
rect 19156 6258 19208 6264
rect 19156 5568 19208 5574
rect 19156 5510 19208 5516
rect 19168 5234 19196 5510
rect 19156 5228 19208 5234
rect 19156 5170 19208 5176
rect 19352 5114 19380 8230
rect 19444 6798 19472 8384
rect 19996 8362 20024 8978
rect 20088 8634 20116 9318
rect 20272 8922 20300 11512
rect 20364 9110 20392 12294
rect 20456 9518 20484 15846
rect 20548 10538 20576 17818
rect 20628 17604 20680 17610
rect 20732 17592 20760 18090
rect 20824 17678 20852 18566
rect 20916 18426 20944 18566
rect 20994 18456 21050 18465
rect 20904 18420 20956 18426
rect 20994 18391 21050 18400
rect 20904 18362 20956 18368
rect 20904 17808 20956 17814
rect 20904 17750 20956 17756
rect 20812 17672 20864 17678
rect 20812 17614 20864 17620
rect 20680 17564 20760 17592
rect 20628 17546 20680 17552
rect 20640 17184 20668 17546
rect 20916 17202 20944 17750
rect 20812 17196 20864 17202
rect 20640 17156 20812 17184
rect 20812 17138 20864 17144
rect 20904 17196 20956 17202
rect 20904 17138 20956 17144
rect 20628 16992 20680 16998
rect 20628 16934 20680 16940
rect 20536 10532 20588 10538
rect 20536 10474 20588 10480
rect 20640 10418 20668 16934
rect 20824 15706 20852 17138
rect 20916 17066 20944 17138
rect 20904 17060 20956 17066
rect 20904 17002 20956 17008
rect 20904 15904 20956 15910
rect 20904 15846 20956 15852
rect 20812 15700 20864 15706
rect 20812 15642 20864 15648
rect 20720 15564 20772 15570
rect 20720 15506 20772 15512
rect 20732 15026 20760 15506
rect 20720 15020 20772 15026
rect 20720 14962 20772 14968
rect 20720 14408 20772 14414
rect 20720 14350 20772 14356
rect 20732 14278 20760 14350
rect 20720 14272 20772 14278
rect 20720 14214 20772 14220
rect 20718 13560 20774 13569
rect 20718 13495 20774 13504
rect 20732 13326 20760 13495
rect 20720 13320 20772 13326
rect 20720 13262 20772 13268
rect 20732 13190 20760 13262
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 20732 11286 20760 13126
rect 20720 11280 20772 11286
rect 20720 11222 20772 11228
rect 20812 11008 20864 11014
rect 20812 10950 20864 10956
rect 20824 10606 20852 10950
rect 20812 10600 20864 10606
rect 20812 10542 20864 10548
rect 20548 10390 20668 10418
rect 20444 9512 20496 9518
rect 20444 9454 20496 9460
rect 20352 9104 20404 9110
rect 20352 9046 20404 9052
rect 20548 9042 20576 10390
rect 20628 10260 20680 10266
rect 20628 10202 20680 10208
rect 20640 9654 20668 10202
rect 20812 10124 20864 10130
rect 20812 10066 20864 10072
rect 20720 9920 20772 9926
rect 20720 9862 20772 9868
rect 20628 9648 20680 9654
rect 20628 9590 20680 9596
rect 20536 9036 20588 9042
rect 20536 8978 20588 8984
rect 20272 8894 20392 8922
rect 20732 8906 20760 9862
rect 20824 9761 20852 10066
rect 20810 9752 20866 9761
rect 20810 9687 20866 9696
rect 20076 8628 20128 8634
rect 20076 8570 20128 8576
rect 20260 8628 20312 8634
rect 20260 8570 20312 8576
rect 19984 8356 20036 8362
rect 20088 8344 20116 8570
rect 20272 8537 20300 8570
rect 20258 8528 20314 8537
rect 20258 8463 20314 8472
rect 20088 8316 20208 8344
rect 19984 8298 20036 8304
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19984 7472 20036 7478
rect 19984 7414 20036 7420
rect 19708 7268 19760 7274
rect 19708 7210 19760 7216
rect 19432 6792 19484 6798
rect 19720 6780 19748 7210
rect 19800 6792 19852 6798
rect 19720 6752 19800 6780
rect 19432 6734 19484 6740
rect 19800 6734 19852 6740
rect 19996 6662 20024 7414
rect 20180 6798 20208 8316
rect 20260 7200 20312 7206
rect 20260 7142 20312 7148
rect 20168 6792 20220 6798
rect 20168 6734 20220 6740
rect 19432 6656 19484 6662
rect 19432 6598 19484 6604
rect 19984 6656 20036 6662
rect 19984 6598 20036 6604
rect 19444 6458 19472 6598
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19432 6452 19484 6458
rect 19432 6394 19484 6400
rect 19996 6322 20024 6598
rect 19984 6316 20036 6322
rect 19984 6258 20036 6264
rect 19982 6216 20038 6225
rect 19982 6151 20038 6160
rect 19432 5772 19484 5778
rect 19432 5714 19484 5720
rect 19260 5086 19380 5114
rect 19444 5098 19472 5714
rect 19616 5704 19668 5710
rect 19614 5672 19616 5681
rect 19668 5672 19670 5681
rect 19614 5607 19670 5616
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19996 5166 20024 6151
rect 20076 6112 20128 6118
rect 20076 6054 20128 6060
rect 19984 5160 20036 5166
rect 19984 5102 20036 5108
rect 20088 5114 20116 6054
rect 20180 5710 20208 6734
rect 20272 5778 20300 7142
rect 20260 5772 20312 5778
rect 20260 5714 20312 5720
rect 20168 5704 20220 5710
rect 20168 5646 20220 5652
rect 20260 5568 20312 5574
rect 20260 5510 20312 5516
rect 19432 5092 19484 5098
rect 19156 4616 19208 4622
rect 19156 4558 19208 4564
rect 19064 4208 19116 4214
rect 19064 4150 19116 4156
rect 18972 4004 19024 4010
rect 18972 3946 19024 3952
rect 18892 3726 19012 3754
rect 18984 3670 19012 3726
rect 18972 3664 19024 3670
rect 18972 3606 19024 3612
rect 18880 3596 18932 3602
rect 18880 3538 18932 3544
rect 18788 2304 18840 2310
rect 18788 2246 18840 2252
rect 18892 800 18920 3538
rect 19076 2774 19104 4150
rect 19168 3074 19196 4558
rect 19260 3641 19288 5086
rect 20088 5086 20208 5114
rect 19432 5034 19484 5040
rect 19340 5024 19392 5030
rect 19340 4966 19392 4972
rect 19984 5024 20036 5030
rect 19984 4966 20036 4972
rect 20076 5024 20128 5030
rect 20076 4966 20128 4972
rect 19352 3754 19380 4966
rect 19996 4622 20024 4966
rect 19984 4616 20036 4622
rect 19984 4558 20036 4564
rect 19432 4480 19484 4486
rect 19432 4422 19484 4428
rect 19444 4282 19472 4422
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19432 4276 19484 4282
rect 19432 4218 19484 4224
rect 19352 3726 19472 3754
rect 19340 3664 19392 3670
rect 19246 3632 19302 3641
rect 19340 3606 19392 3612
rect 19246 3567 19302 3576
rect 19352 3194 19380 3606
rect 19444 3466 19472 3726
rect 20088 3602 20116 4966
rect 20180 4078 20208 5086
rect 20272 4758 20300 5510
rect 20260 4752 20312 4758
rect 20260 4694 20312 4700
rect 20168 4072 20220 4078
rect 20168 4014 20220 4020
rect 20260 4004 20312 4010
rect 20260 3946 20312 3952
rect 20076 3596 20128 3602
rect 20076 3538 20128 3544
rect 19984 3528 20036 3534
rect 19984 3470 20036 3476
rect 20074 3496 20130 3505
rect 19432 3460 19484 3466
rect 19432 3402 19484 3408
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 19432 3188 19484 3194
rect 19432 3130 19484 3136
rect 19168 3046 19380 3074
rect 19076 2746 19196 2774
rect 19168 800 19196 2746
rect 19248 2304 19300 2310
rect 19248 2246 19300 2252
rect 19260 800 19288 2246
rect 19352 898 19380 3046
rect 19444 1442 19472 3130
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19800 1760 19852 1766
rect 19800 1702 19852 1708
rect 19444 1414 19748 1442
rect 19524 1352 19576 1358
rect 19524 1294 19576 1300
rect 19352 870 19472 898
rect 19444 800 19472 870
rect 19536 800 19564 1294
rect 19720 800 19748 1414
rect 19812 800 19840 1702
rect 19996 800 20024 3470
rect 20074 3431 20076 3440
rect 20128 3431 20130 3440
rect 20076 3402 20128 3408
rect 20168 3392 20220 3398
rect 20168 3334 20220 3340
rect 20180 3074 20208 3334
rect 20272 3194 20300 3946
rect 20260 3188 20312 3194
rect 20260 3130 20312 3136
rect 20088 3058 20208 3074
rect 20076 3052 20208 3058
rect 20128 3046 20208 3052
rect 20076 2994 20128 3000
rect 20088 800 20116 2994
rect 20260 2916 20312 2922
rect 20260 2858 20312 2864
rect 20168 2848 20220 2854
rect 20168 2790 20220 2796
rect 20180 1358 20208 2790
rect 20168 1352 20220 1358
rect 20168 1294 20220 1300
rect 20272 800 20300 2858
rect 20364 2106 20392 8894
rect 20720 8900 20772 8906
rect 20720 8842 20772 8848
rect 20444 8832 20496 8838
rect 20444 8774 20496 8780
rect 20456 8430 20484 8774
rect 20444 8424 20496 8430
rect 20444 8366 20496 8372
rect 20536 8356 20588 8362
rect 20536 8298 20588 8304
rect 20548 7886 20576 8298
rect 20536 7880 20588 7886
rect 20536 7822 20588 7828
rect 20444 7744 20496 7750
rect 20444 7686 20496 7692
rect 20456 5250 20484 7686
rect 20548 6866 20576 7822
rect 20536 6860 20588 6866
rect 20536 6802 20588 6808
rect 20732 6322 20760 8842
rect 20812 8560 20864 8566
rect 20812 8502 20864 8508
rect 20824 7886 20852 8502
rect 20916 8294 20944 15846
rect 21008 15094 21036 18391
rect 21088 18352 21140 18358
rect 21086 18320 21088 18329
rect 21180 18352 21232 18358
rect 21140 18320 21142 18329
rect 21180 18294 21232 18300
rect 21086 18255 21142 18264
rect 21192 17610 21220 18294
rect 21284 18290 21312 18906
rect 21376 18834 21404 19246
rect 21364 18828 21416 18834
rect 21364 18770 21416 18776
rect 21272 18284 21324 18290
rect 21272 18226 21324 18232
rect 21362 17640 21418 17649
rect 21180 17604 21232 17610
rect 21362 17575 21364 17584
rect 21180 17546 21232 17552
rect 21416 17575 21418 17584
rect 21364 17546 21416 17552
rect 21272 17536 21324 17542
rect 21272 17478 21324 17484
rect 21088 16720 21140 16726
rect 21088 16662 21140 16668
rect 20996 15088 21048 15094
rect 20996 15030 21048 15036
rect 21100 11014 21128 16662
rect 21284 16522 21312 17478
rect 21364 16720 21416 16726
rect 21364 16662 21416 16668
rect 21272 16516 21324 16522
rect 21272 16458 21324 16464
rect 21272 13728 21324 13734
rect 21272 13670 21324 13676
rect 21284 12850 21312 13670
rect 21272 12844 21324 12850
rect 21272 12786 21324 12792
rect 21272 12164 21324 12170
rect 21272 12106 21324 12112
rect 21284 11898 21312 12106
rect 21272 11892 21324 11898
rect 21272 11834 21324 11840
rect 21284 11558 21312 11834
rect 21272 11552 21324 11558
rect 21272 11494 21324 11500
rect 21376 11150 21404 16662
rect 21560 12434 21588 20198
rect 21822 20159 21878 20168
rect 21640 18828 21692 18834
rect 21640 18770 21692 18776
rect 21652 16454 21680 18770
rect 21836 16590 21864 20159
rect 22112 18766 22140 23462
rect 22008 18760 22060 18766
rect 22008 18702 22060 18708
rect 22100 18760 22152 18766
rect 22100 18702 22152 18708
rect 21916 18420 21968 18426
rect 22020 18408 22048 18702
rect 21968 18380 22048 18408
rect 21916 18362 21968 18368
rect 22100 17196 22152 17202
rect 22100 17138 22152 17144
rect 22112 16794 22140 17138
rect 22100 16788 22152 16794
rect 22100 16730 22152 16736
rect 21824 16584 21876 16590
rect 21824 16526 21876 16532
rect 21640 16448 21692 16454
rect 21836 16425 21864 16526
rect 21640 16390 21692 16396
rect 21822 16416 21878 16425
rect 21822 16351 21878 16360
rect 21836 16250 21864 16351
rect 21824 16244 21876 16250
rect 21824 16186 21876 16192
rect 21824 16040 21876 16046
rect 21824 15982 21876 15988
rect 21836 15706 21864 15982
rect 21824 15700 21876 15706
rect 21824 15642 21876 15648
rect 22008 15496 22060 15502
rect 22008 15438 22060 15444
rect 22100 15496 22152 15502
rect 22100 15438 22152 15444
rect 22020 15162 22048 15438
rect 22008 15156 22060 15162
rect 22008 15098 22060 15104
rect 22008 15020 22060 15026
rect 22008 14962 22060 14968
rect 22020 14929 22048 14962
rect 22006 14920 22062 14929
rect 22006 14855 22062 14864
rect 22112 12986 22140 15438
rect 22204 15144 22232 24126
rect 22388 22030 22416 24142
rect 22376 22024 22428 22030
rect 22376 21966 22428 21972
rect 22388 21690 22416 21966
rect 22376 21684 22428 21690
rect 22376 21626 22428 21632
rect 22388 20942 22416 21626
rect 22468 21140 22520 21146
rect 22468 21082 22520 21088
rect 22376 20936 22428 20942
rect 22376 20878 22428 20884
rect 22284 20596 22336 20602
rect 22284 20538 22336 20544
rect 22296 18426 22324 20538
rect 22376 19712 22428 19718
rect 22480 19666 22508 21082
rect 22428 19660 22508 19666
rect 22376 19654 22508 19660
rect 22388 19638 22508 19654
rect 22480 18766 22508 19638
rect 22572 19417 22600 26998
rect 23204 26988 23256 26994
rect 23204 26930 23256 26936
rect 22744 26376 22796 26382
rect 22744 26318 22796 26324
rect 22756 25294 22784 26318
rect 23216 26314 23244 26930
rect 23584 26858 23612 27406
rect 23572 26852 23624 26858
rect 23572 26794 23624 26800
rect 23400 26314 23612 26330
rect 23204 26308 23256 26314
rect 23204 26250 23256 26256
rect 23400 26308 23624 26314
rect 23400 26302 23572 26308
rect 22744 25288 22796 25294
rect 22744 25230 22796 25236
rect 23216 24138 23244 26250
rect 23296 25152 23348 25158
rect 23296 25094 23348 25100
rect 23308 24206 23336 25094
rect 23296 24200 23348 24206
rect 23296 24142 23348 24148
rect 23204 24132 23256 24138
rect 23204 24074 23256 24080
rect 23308 23780 23336 24142
rect 23216 23752 23336 23780
rect 23112 23724 23164 23730
rect 23112 23666 23164 23672
rect 22744 23588 22796 23594
rect 22744 23530 22796 23536
rect 22652 23112 22704 23118
rect 22652 23054 22704 23060
rect 22664 22778 22692 23054
rect 22652 22772 22704 22778
rect 22652 22714 22704 22720
rect 22652 22092 22704 22098
rect 22652 22034 22704 22040
rect 22664 20942 22692 22034
rect 22756 21146 22784 23530
rect 22836 23112 22888 23118
rect 22836 23054 22888 23060
rect 22848 22234 22876 23054
rect 23124 23050 23152 23666
rect 23112 23044 23164 23050
rect 23112 22986 23164 22992
rect 22928 22432 22980 22438
rect 22928 22374 22980 22380
rect 22836 22228 22888 22234
rect 22836 22170 22888 22176
rect 22940 22094 22968 22374
rect 23124 22234 23152 22986
rect 23112 22228 23164 22234
rect 23112 22170 23164 22176
rect 22848 22066 22968 22094
rect 22848 21962 22876 22066
rect 22836 21956 22888 21962
rect 22836 21898 22888 21904
rect 22744 21140 22796 21146
rect 22744 21082 22796 21088
rect 22652 20936 22704 20942
rect 22744 20936 22796 20942
rect 22652 20878 22704 20884
rect 22742 20904 22744 20913
rect 22796 20904 22798 20913
rect 22742 20839 22798 20848
rect 22652 19780 22704 19786
rect 22652 19722 22704 19728
rect 22558 19408 22614 19417
rect 22558 19343 22614 19352
rect 22468 18760 22520 18766
rect 22468 18702 22520 18708
rect 22284 18420 22336 18426
rect 22284 18362 22336 18368
rect 22296 17882 22324 18362
rect 22284 17876 22336 17882
rect 22284 17818 22336 17824
rect 22664 16658 22692 19722
rect 22756 19514 22784 20839
rect 22744 19508 22796 19514
rect 22744 19450 22796 19456
rect 22848 19242 22876 21898
rect 23124 21554 23152 22170
rect 23112 21548 23164 21554
rect 23112 21490 23164 21496
rect 22928 20596 22980 20602
rect 22928 20538 22980 20544
rect 22940 19922 22968 20538
rect 23216 20466 23244 23752
rect 23296 22976 23348 22982
rect 23296 22918 23348 22924
rect 23308 22710 23336 22918
rect 23296 22704 23348 22710
rect 23296 22646 23348 22652
rect 23400 21010 23428 26302
rect 23572 26250 23624 26256
rect 23676 25702 23704 31232
rect 25596 31204 25648 31210
rect 25596 31146 25648 31152
rect 24860 31136 24912 31142
rect 24860 31078 24912 31084
rect 24032 30728 24084 30734
rect 24032 30670 24084 30676
rect 24044 30258 24072 30670
rect 24032 30252 24084 30258
rect 24032 30194 24084 30200
rect 24044 29238 24072 30194
rect 24032 29232 24084 29238
rect 24032 29174 24084 29180
rect 23848 29164 23900 29170
rect 23848 29106 23900 29112
rect 23756 29028 23808 29034
rect 23756 28970 23808 28976
rect 23768 27062 23796 28970
rect 23860 27606 23888 29106
rect 24044 28626 24072 29174
rect 24032 28620 24084 28626
rect 24032 28562 24084 28568
rect 24676 27872 24728 27878
rect 24676 27814 24728 27820
rect 24688 27674 24716 27814
rect 24676 27668 24728 27674
rect 24676 27610 24728 27616
rect 24872 27606 24900 31078
rect 25608 30258 25636 31146
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 65654 31036 65962 31045
rect 65654 31034 65660 31036
rect 65716 31034 65740 31036
rect 65796 31034 65820 31036
rect 65876 31034 65900 31036
rect 65956 31034 65962 31036
rect 65716 30982 65718 31034
rect 65898 30982 65900 31034
rect 65654 30980 65660 30982
rect 65716 30980 65740 30982
rect 65796 30980 65820 30982
rect 65876 30980 65900 30982
rect 65956 30980 65962 30982
rect 65654 30971 65962 30980
rect 68100 30728 68152 30734
rect 68098 30696 68100 30705
rect 68152 30696 68154 30705
rect 68098 30631 68154 30640
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 25596 30252 25648 30258
rect 25596 30194 25648 30200
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 65654 29948 65962 29957
rect 65654 29946 65660 29948
rect 65716 29946 65740 29948
rect 65796 29946 65820 29948
rect 65876 29946 65900 29948
rect 65956 29946 65962 29948
rect 65716 29894 65718 29946
rect 65898 29894 65900 29946
rect 65654 29892 65660 29894
rect 65716 29892 65740 29894
rect 65796 29892 65820 29894
rect 65876 29892 65900 29894
rect 65956 29892 65962 29894
rect 65654 29883 65962 29892
rect 26976 29640 27028 29646
rect 26976 29582 27028 29588
rect 68100 29640 68152 29646
rect 68100 29582 68152 29588
rect 26240 29572 26292 29578
rect 26240 29514 26292 29520
rect 25228 29504 25280 29510
rect 25228 29446 25280 29452
rect 25504 29504 25556 29510
rect 25504 29446 25556 29452
rect 25136 28076 25188 28082
rect 25136 28018 25188 28024
rect 23848 27600 23900 27606
rect 23848 27542 23900 27548
rect 24860 27600 24912 27606
rect 24860 27542 24912 27548
rect 24952 27532 25004 27538
rect 24952 27474 25004 27480
rect 24216 27464 24268 27470
rect 24214 27432 24216 27441
rect 24268 27432 24270 27441
rect 24214 27367 24270 27376
rect 23756 27056 23808 27062
rect 23756 26998 23808 27004
rect 23848 26240 23900 26246
rect 23848 26182 23900 26188
rect 23860 25974 23888 26182
rect 23848 25968 23900 25974
rect 23848 25910 23900 25916
rect 24228 25906 24256 27367
rect 24860 26308 24912 26314
rect 24860 26250 24912 26256
rect 24872 26042 24900 26250
rect 24860 26036 24912 26042
rect 24860 25978 24912 25984
rect 24216 25900 24268 25906
rect 24216 25842 24268 25848
rect 24584 25900 24636 25906
rect 24584 25842 24636 25848
rect 23756 25832 23808 25838
rect 23756 25774 23808 25780
rect 23664 25696 23716 25702
rect 23664 25638 23716 25644
rect 23768 25514 23796 25774
rect 23676 25486 23796 25514
rect 23480 25220 23532 25226
rect 23480 25162 23532 25168
rect 23492 24954 23520 25162
rect 23480 24948 23532 24954
rect 23480 24890 23532 24896
rect 23676 24750 23704 25486
rect 24228 24818 24256 25842
rect 24596 25702 24624 25842
rect 24964 25838 24992 27474
rect 25148 27470 25176 28018
rect 25136 27464 25188 27470
rect 25136 27406 25188 27412
rect 24952 25832 25004 25838
rect 24952 25774 25004 25780
rect 24584 25696 24636 25702
rect 24584 25638 24636 25644
rect 23756 24812 23808 24818
rect 23756 24754 23808 24760
rect 23940 24812 23992 24818
rect 23940 24754 23992 24760
rect 24216 24812 24268 24818
rect 24216 24754 24268 24760
rect 24584 24812 24636 24818
rect 24584 24754 24636 24760
rect 24860 24812 24912 24818
rect 24860 24754 24912 24760
rect 23664 24744 23716 24750
rect 23664 24686 23716 24692
rect 23676 23662 23704 24686
rect 23768 24138 23796 24754
rect 23952 24410 23980 24754
rect 23940 24404 23992 24410
rect 23940 24346 23992 24352
rect 23756 24132 23808 24138
rect 23756 24074 23808 24080
rect 24596 23730 24624 24754
rect 24872 24070 24900 24754
rect 24860 24064 24912 24070
rect 24860 24006 24912 24012
rect 24584 23724 24636 23730
rect 24584 23666 24636 23672
rect 23664 23656 23716 23662
rect 23664 23598 23716 23604
rect 23756 23248 23808 23254
rect 23756 23190 23808 23196
rect 23768 22982 23796 23190
rect 23756 22976 23808 22982
rect 23756 22918 23808 22924
rect 23768 22234 23796 22918
rect 24584 22568 24636 22574
rect 24584 22510 24636 22516
rect 23756 22228 23808 22234
rect 23756 22170 23808 22176
rect 23572 22024 23624 22030
rect 23572 21966 23624 21972
rect 23584 21486 23612 21966
rect 23664 21548 23716 21554
rect 23664 21490 23716 21496
rect 23572 21480 23624 21486
rect 23478 21448 23534 21457
rect 23572 21422 23624 21428
rect 23478 21383 23534 21392
rect 23388 21004 23440 21010
rect 23388 20946 23440 20952
rect 23492 20942 23520 21383
rect 23480 20936 23532 20942
rect 23480 20878 23532 20884
rect 23388 20868 23440 20874
rect 23388 20810 23440 20816
rect 23400 20754 23428 20810
rect 23584 20754 23612 21422
rect 23676 20942 23704 21490
rect 23664 20936 23716 20942
rect 23664 20878 23716 20884
rect 23400 20726 23612 20754
rect 23492 20534 23520 20726
rect 23480 20528 23532 20534
rect 23572 20528 23624 20534
rect 23480 20470 23532 20476
rect 23570 20496 23572 20505
rect 23624 20496 23626 20505
rect 23204 20460 23256 20466
rect 23570 20431 23626 20440
rect 23204 20402 23256 20408
rect 23676 20330 23704 20878
rect 23664 20324 23716 20330
rect 23664 20266 23716 20272
rect 23768 19938 23796 22170
rect 24596 20602 24624 22510
rect 24872 21078 24900 24006
rect 24952 23656 25004 23662
rect 24952 23598 25004 23604
rect 24860 21072 24912 21078
rect 24860 21014 24912 21020
rect 24860 20800 24912 20806
rect 24860 20742 24912 20748
rect 24584 20596 24636 20602
rect 24584 20538 24636 20544
rect 24676 20324 24728 20330
rect 24676 20266 24728 20272
rect 23940 20256 23992 20262
rect 23940 20198 23992 20204
rect 22928 19916 22980 19922
rect 22928 19858 22980 19864
rect 23676 19910 23796 19938
rect 23676 19854 23704 19910
rect 23664 19848 23716 19854
rect 23664 19790 23716 19796
rect 22836 19236 22888 19242
rect 22836 19178 22888 19184
rect 23676 19174 23704 19790
rect 23664 19168 23716 19174
rect 23664 19110 23716 19116
rect 23204 17536 23256 17542
rect 23204 17478 23256 17484
rect 23110 17232 23166 17241
rect 23110 17167 23166 17176
rect 22652 16652 22704 16658
rect 22652 16594 22704 16600
rect 23124 16250 23152 17167
rect 23216 16697 23244 17478
rect 23572 17128 23624 17134
rect 23572 17070 23624 17076
rect 23584 16794 23612 17070
rect 23572 16788 23624 16794
rect 23572 16730 23624 16736
rect 23202 16688 23258 16697
rect 23202 16623 23258 16632
rect 23112 16244 23164 16250
rect 23112 16186 23164 16192
rect 22928 16108 22980 16114
rect 22928 16050 22980 16056
rect 22282 16008 22338 16017
rect 22282 15943 22338 15952
rect 22296 15502 22324 15943
rect 22284 15496 22336 15502
rect 22284 15438 22336 15444
rect 22204 15116 22416 15144
rect 22282 15056 22338 15065
rect 22282 14991 22284 15000
rect 22336 14991 22338 15000
rect 22284 14962 22336 14968
rect 22192 14952 22244 14958
rect 22388 14906 22416 15116
rect 22192 14894 22244 14900
rect 22100 12980 22152 12986
rect 22100 12922 22152 12928
rect 22008 12912 22060 12918
rect 22008 12854 22060 12860
rect 21468 12406 21588 12434
rect 21468 11762 21496 12406
rect 21548 12164 21600 12170
rect 21548 12106 21600 12112
rect 21916 12164 21968 12170
rect 22020 12152 22048 12854
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 21968 12124 22048 12152
rect 21916 12106 21968 12112
rect 21456 11756 21508 11762
rect 21456 11698 21508 11704
rect 21468 11218 21496 11698
rect 21456 11212 21508 11218
rect 21456 11154 21508 11160
rect 21364 11144 21416 11150
rect 21362 11112 21364 11121
rect 21416 11112 21418 11121
rect 21362 11047 21418 11056
rect 21088 11008 21140 11014
rect 21088 10950 21140 10956
rect 21560 10674 21588 12106
rect 22112 11898 22140 12786
rect 22204 12442 22232 14894
rect 22296 14878 22416 14906
rect 22940 14890 22968 16050
rect 23216 15473 23244 16623
rect 23202 15464 23258 15473
rect 23202 15399 23258 15408
rect 22928 14884 22980 14890
rect 22296 13938 22324 14878
rect 22928 14826 22980 14832
rect 22376 14816 22428 14822
rect 22376 14758 22428 14764
rect 22388 14482 22416 14758
rect 22468 14544 22520 14550
rect 22468 14486 22520 14492
rect 22376 14476 22428 14482
rect 22376 14418 22428 14424
rect 22284 13932 22336 13938
rect 22284 13874 22336 13880
rect 22284 13184 22336 13190
rect 22284 13126 22336 13132
rect 22192 12436 22244 12442
rect 22192 12378 22244 12384
rect 22296 12170 22324 13126
rect 22376 12844 22428 12850
rect 22376 12786 22428 12792
rect 22388 12238 22416 12786
rect 22376 12232 22428 12238
rect 22376 12174 22428 12180
rect 22284 12164 22336 12170
rect 22284 12106 22336 12112
rect 22100 11892 22152 11898
rect 22100 11834 22152 11840
rect 22192 11824 22244 11830
rect 22192 11766 22244 11772
rect 22204 11354 22232 11766
rect 22376 11552 22428 11558
rect 22376 11494 22428 11500
rect 22192 11348 22244 11354
rect 22192 11290 22244 11296
rect 22204 10674 22232 11290
rect 22388 11082 22416 11494
rect 22376 11076 22428 11082
rect 22376 11018 22428 11024
rect 21548 10668 21600 10674
rect 21548 10610 21600 10616
rect 22192 10668 22244 10674
rect 22192 10610 22244 10616
rect 21088 10464 21140 10470
rect 21088 10406 21140 10412
rect 21100 9926 21128 10406
rect 21088 9920 21140 9926
rect 21088 9862 21140 9868
rect 21560 9518 21588 10610
rect 22204 9654 22232 10610
rect 22192 9648 22244 9654
rect 22192 9590 22244 9596
rect 21548 9512 21600 9518
rect 21548 9454 21600 9460
rect 20904 8288 20956 8294
rect 20904 8230 20956 8236
rect 20812 7880 20864 7886
rect 20812 7822 20864 7828
rect 21560 7410 21588 9454
rect 21916 8968 21968 8974
rect 22480 8945 22508 14486
rect 23952 14414 23980 20198
rect 24492 19848 24544 19854
rect 24492 19790 24544 19796
rect 24504 18970 24532 19790
rect 24688 19718 24716 20266
rect 24768 19916 24820 19922
rect 24768 19858 24820 19864
rect 24676 19712 24728 19718
rect 24676 19654 24728 19660
rect 24492 18964 24544 18970
rect 24492 18906 24544 18912
rect 24124 18692 24176 18698
rect 24124 18634 24176 18640
rect 24136 18358 24164 18634
rect 24124 18352 24176 18358
rect 24124 18294 24176 18300
rect 24400 18216 24452 18222
rect 24400 18158 24452 18164
rect 24308 17740 24360 17746
rect 24308 17682 24360 17688
rect 24320 17134 24348 17682
rect 24308 17128 24360 17134
rect 24308 17070 24360 17076
rect 24320 16454 24348 17070
rect 24412 16794 24440 18158
rect 24504 17610 24532 18906
rect 24584 18624 24636 18630
rect 24584 18566 24636 18572
rect 24596 17678 24624 18566
rect 24780 17882 24808 19858
rect 24768 17876 24820 17882
rect 24768 17818 24820 17824
rect 24584 17672 24636 17678
rect 24584 17614 24636 17620
rect 24492 17604 24544 17610
rect 24492 17546 24544 17552
rect 24676 17604 24728 17610
rect 24676 17546 24728 17552
rect 24492 17332 24544 17338
rect 24492 17274 24544 17280
rect 24504 17202 24532 17274
rect 24492 17196 24544 17202
rect 24492 17138 24544 17144
rect 24400 16788 24452 16794
rect 24400 16730 24452 16736
rect 24504 16726 24532 17138
rect 24492 16720 24544 16726
rect 24492 16662 24544 16668
rect 24308 16448 24360 16454
rect 24308 16390 24360 16396
rect 24308 14952 24360 14958
rect 24308 14894 24360 14900
rect 23940 14408 23992 14414
rect 23940 14350 23992 14356
rect 22928 14272 22980 14278
rect 22928 14214 22980 14220
rect 22652 13932 22704 13938
rect 22652 13874 22704 13880
rect 22560 13184 22612 13190
rect 22560 13126 22612 13132
rect 22572 12918 22600 13126
rect 22560 12912 22612 12918
rect 22560 12854 22612 12860
rect 22664 10305 22692 13874
rect 22836 10600 22888 10606
rect 22836 10542 22888 10548
rect 22650 10296 22706 10305
rect 22848 10266 22876 10542
rect 22650 10231 22706 10240
rect 22836 10260 22888 10266
rect 22836 10202 22888 10208
rect 22940 9586 22968 14214
rect 23388 14000 23440 14006
rect 23388 13942 23440 13948
rect 23400 12986 23428 13942
rect 23572 13932 23624 13938
rect 23572 13874 23624 13880
rect 23584 13297 23612 13874
rect 23664 13864 23716 13870
rect 23664 13806 23716 13812
rect 23570 13288 23626 13297
rect 23570 13223 23626 13232
rect 23388 12980 23440 12986
rect 23388 12922 23440 12928
rect 23480 12844 23532 12850
rect 23480 12786 23532 12792
rect 23492 12753 23520 12786
rect 23478 12744 23534 12753
rect 23478 12679 23534 12688
rect 23020 12232 23072 12238
rect 23020 12174 23072 12180
rect 23032 10674 23060 12174
rect 23020 10668 23072 10674
rect 23020 10610 23072 10616
rect 23572 10464 23624 10470
rect 23572 10406 23624 10412
rect 23584 10062 23612 10406
rect 23572 10056 23624 10062
rect 23572 9998 23624 10004
rect 22928 9580 22980 9586
rect 22928 9522 22980 9528
rect 23388 8968 23440 8974
rect 21916 8910 21968 8916
rect 22466 8936 22522 8945
rect 21928 8498 21956 8910
rect 23388 8910 23440 8916
rect 22466 8871 22522 8880
rect 23204 8832 23256 8838
rect 23204 8774 23256 8780
rect 23216 8566 23244 8774
rect 23204 8560 23256 8566
rect 23204 8502 23256 8508
rect 21916 8492 21968 8498
rect 21916 8434 21968 8440
rect 23112 8492 23164 8498
rect 23112 8434 23164 8440
rect 21928 8090 21956 8434
rect 21916 8084 21968 8090
rect 21916 8026 21968 8032
rect 23124 7818 23152 8434
rect 22652 7812 22704 7818
rect 22652 7754 22704 7760
rect 23112 7812 23164 7818
rect 23112 7754 23164 7760
rect 22664 7410 22692 7754
rect 21548 7404 21600 7410
rect 21548 7346 21600 7352
rect 22652 7404 22704 7410
rect 22652 7346 22704 7352
rect 21560 6866 21588 7346
rect 22376 7336 22428 7342
rect 22376 7278 22428 7284
rect 21548 6860 21600 6866
rect 21548 6802 21600 6808
rect 22388 6798 22416 7278
rect 22376 6792 22428 6798
rect 22376 6734 22428 6740
rect 23400 6390 23428 8910
rect 23676 8634 23704 13806
rect 24320 13394 24348 14894
rect 24492 13932 24544 13938
rect 24492 13874 24544 13880
rect 23848 13388 23900 13394
rect 23848 13330 23900 13336
rect 24308 13388 24360 13394
rect 24308 13330 24360 13336
rect 23756 12776 23808 12782
rect 23756 12718 23808 12724
rect 23664 8628 23716 8634
rect 23664 8570 23716 8576
rect 23572 8492 23624 8498
rect 23572 8434 23624 8440
rect 23584 8362 23612 8434
rect 23572 8356 23624 8362
rect 23572 8298 23624 8304
rect 23480 7948 23532 7954
rect 23480 7890 23532 7896
rect 23388 6384 23440 6390
rect 23388 6326 23440 6332
rect 20720 6316 20772 6322
rect 20720 6258 20772 6264
rect 22100 6316 22152 6322
rect 22100 6258 22152 6264
rect 22112 5778 22140 6258
rect 23020 6112 23072 6118
rect 23020 6054 23072 6060
rect 22100 5772 22152 5778
rect 22100 5714 22152 5720
rect 21272 5296 21324 5302
rect 20456 5222 20576 5250
rect 21272 5238 21324 5244
rect 20444 5160 20496 5166
rect 20444 5102 20496 5108
rect 20456 4282 20484 5102
rect 20444 4276 20496 4282
rect 20444 4218 20496 4224
rect 20444 3936 20496 3942
rect 20444 3878 20496 3884
rect 20352 2100 20404 2106
rect 20352 2042 20404 2048
rect 20456 800 20484 3878
rect 20548 2378 20576 5222
rect 21284 4554 21312 5238
rect 22008 5228 22060 5234
rect 22008 5170 22060 5176
rect 21272 4548 21324 4554
rect 21272 4490 21324 4496
rect 21180 3936 21232 3942
rect 21180 3878 21232 3884
rect 21192 3738 21220 3878
rect 21180 3732 21232 3738
rect 21180 3674 21232 3680
rect 20996 3528 21048 3534
rect 20996 3470 21048 3476
rect 20628 3120 20680 3126
rect 20628 3062 20680 3068
rect 20536 2372 20588 2378
rect 20536 2314 20588 2320
rect 20640 2310 20668 3062
rect 20720 2984 20772 2990
rect 20720 2926 20772 2932
rect 20628 2304 20680 2310
rect 20628 2246 20680 2252
rect 20640 1766 20668 2246
rect 20628 1760 20680 1766
rect 20628 1702 20680 1708
rect 20732 800 20760 2926
rect 21008 800 21036 3470
rect 22020 3194 22048 5170
rect 22112 4826 22140 5714
rect 23032 5574 23060 6054
rect 23492 5914 23520 7890
rect 23584 7886 23612 8298
rect 23768 8090 23796 12718
rect 23860 11694 23888 13330
rect 23940 12844 23992 12850
rect 23940 12786 23992 12792
rect 24308 12844 24360 12850
rect 24308 12786 24360 12792
rect 23952 12434 23980 12786
rect 23952 12406 24164 12434
rect 23940 12368 23992 12374
rect 23940 12310 23992 12316
rect 23848 11688 23900 11694
rect 23848 11630 23900 11636
rect 23952 11354 23980 12310
rect 23940 11348 23992 11354
rect 23940 11290 23992 11296
rect 23952 10810 23980 11290
rect 24136 11234 24164 12406
rect 24320 12170 24348 12786
rect 24308 12164 24360 12170
rect 24308 12106 24360 12112
rect 24320 11762 24348 12106
rect 24216 11756 24268 11762
rect 24216 11698 24268 11704
rect 24308 11756 24360 11762
rect 24308 11698 24360 11704
rect 24228 11354 24256 11698
rect 24216 11348 24268 11354
rect 24216 11290 24268 11296
rect 24136 11206 24256 11234
rect 23940 10804 23992 10810
rect 23940 10746 23992 10752
rect 23952 10690 23980 10746
rect 23952 10674 24164 10690
rect 23952 10668 24176 10674
rect 23952 10662 24124 10668
rect 24124 10610 24176 10616
rect 24124 9376 24176 9382
rect 24124 9318 24176 9324
rect 24136 8906 24164 9318
rect 24124 8900 24176 8906
rect 24124 8842 24176 8848
rect 24228 8401 24256 11206
rect 24320 10266 24348 11698
rect 24308 10260 24360 10266
rect 24308 10202 24360 10208
rect 24400 10056 24452 10062
rect 24400 9998 24452 10004
rect 24308 9580 24360 9586
rect 24308 9522 24360 9528
rect 24320 8634 24348 9522
rect 24412 8906 24440 9998
rect 24504 9217 24532 13874
rect 24688 12889 24716 17546
rect 24872 16046 24900 20742
rect 24964 19938 24992 23598
rect 25240 22710 25268 29446
rect 25412 28212 25464 28218
rect 25412 28154 25464 28160
rect 25320 27940 25372 27946
rect 25320 27882 25372 27888
rect 25332 27130 25360 27882
rect 25424 27606 25452 28154
rect 25412 27600 25464 27606
rect 25412 27542 25464 27548
rect 25320 27124 25372 27130
rect 25320 27066 25372 27072
rect 25516 26994 25544 29446
rect 25688 28484 25740 28490
rect 25688 28426 25740 28432
rect 25700 27674 25728 28426
rect 26252 28218 26280 29514
rect 26988 29238 27016 29582
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 68112 29345 68140 29582
rect 68098 29336 68154 29345
rect 68098 29271 68154 29280
rect 26976 29232 27028 29238
rect 26976 29174 27028 29180
rect 29092 29164 29144 29170
rect 29092 29106 29144 29112
rect 29000 28552 29052 28558
rect 29000 28494 29052 28500
rect 27712 28484 27764 28490
rect 27712 28426 27764 28432
rect 26424 28416 26476 28422
rect 26424 28358 26476 28364
rect 27620 28416 27672 28422
rect 27620 28358 27672 28364
rect 26240 28212 26292 28218
rect 26240 28154 26292 28160
rect 26332 27872 26384 27878
rect 26332 27814 26384 27820
rect 25688 27668 25740 27674
rect 25688 27610 25740 27616
rect 26056 27464 26108 27470
rect 26056 27406 26108 27412
rect 25504 26988 25556 26994
rect 25504 26930 25556 26936
rect 25412 25900 25464 25906
rect 25412 25842 25464 25848
rect 25424 24818 25452 25842
rect 25412 24812 25464 24818
rect 25412 24754 25464 24760
rect 25424 23526 25452 24754
rect 25412 23520 25464 23526
rect 25412 23462 25464 23468
rect 25228 22704 25280 22710
rect 25228 22646 25280 22652
rect 25240 22506 25268 22646
rect 25228 22500 25280 22506
rect 25228 22442 25280 22448
rect 25516 22094 25544 26930
rect 25964 26308 26016 26314
rect 25964 26250 26016 26256
rect 25688 25152 25740 25158
rect 25688 25094 25740 25100
rect 25700 24818 25728 25094
rect 25688 24812 25740 24818
rect 25688 24754 25740 24760
rect 25596 23792 25648 23798
rect 25596 23734 25648 23740
rect 25608 23322 25636 23734
rect 25596 23316 25648 23322
rect 25648 23276 25820 23304
rect 25596 23258 25648 23264
rect 25516 22066 25728 22094
rect 25320 21888 25372 21894
rect 25320 21830 25372 21836
rect 25136 20800 25188 20806
rect 25136 20742 25188 20748
rect 25148 20448 25176 20742
rect 25228 20460 25280 20466
rect 25148 20420 25228 20448
rect 25228 20402 25280 20408
rect 24964 19922 25176 19938
rect 24964 19916 25188 19922
rect 24964 19910 25136 19916
rect 25136 19858 25188 19864
rect 24952 19780 25004 19786
rect 24952 19722 25004 19728
rect 24964 18766 24992 19722
rect 25044 19712 25096 19718
rect 25044 19654 25096 19660
rect 24952 18760 25004 18766
rect 24952 18702 25004 18708
rect 24860 16040 24912 16046
rect 24860 15982 24912 15988
rect 24858 15736 24914 15745
rect 24858 15671 24914 15680
rect 24872 15570 24900 15671
rect 24860 15564 24912 15570
rect 24860 15506 24912 15512
rect 24872 15094 24900 15506
rect 24860 15088 24912 15094
rect 24860 15030 24912 15036
rect 24952 15020 25004 15026
rect 24952 14962 25004 14968
rect 24964 14618 24992 14962
rect 24952 14612 25004 14618
rect 24952 14554 25004 14560
rect 24952 14272 25004 14278
rect 24952 14214 25004 14220
rect 24964 13977 24992 14214
rect 24950 13968 25006 13977
rect 24950 13903 24952 13912
rect 25004 13903 25006 13912
rect 24952 13874 25004 13880
rect 24768 13728 24820 13734
rect 24768 13670 24820 13676
rect 24780 13326 24808 13670
rect 24952 13388 25004 13394
rect 24952 13330 25004 13336
rect 24768 13320 24820 13326
rect 24768 13262 24820 13268
rect 24674 12880 24730 12889
rect 24674 12815 24730 12824
rect 24964 12442 24992 13330
rect 24952 12436 25004 12442
rect 24952 12378 25004 12384
rect 24768 12096 24820 12102
rect 24964 12050 24992 12378
rect 24768 12038 24820 12044
rect 24780 11150 24808 12038
rect 24872 12022 24992 12050
rect 24872 11354 24900 12022
rect 25056 11914 25084 19654
rect 25148 19310 25176 19858
rect 25240 19854 25268 20402
rect 25228 19848 25280 19854
rect 25228 19790 25280 19796
rect 25136 19304 25188 19310
rect 25136 19246 25188 19252
rect 25240 18222 25268 19790
rect 25228 18216 25280 18222
rect 25228 18158 25280 18164
rect 25136 17672 25188 17678
rect 25136 17614 25188 17620
rect 25148 17202 25176 17614
rect 25332 17338 25360 21830
rect 25412 21548 25464 21554
rect 25412 21490 25464 21496
rect 25424 20942 25452 21490
rect 25504 21480 25556 21486
rect 25504 21422 25556 21428
rect 25412 20936 25464 20942
rect 25410 20904 25412 20913
rect 25464 20904 25466 20913
rect 25410 20839 25466 20848
rect 25424 20448 25452 20839
rect 25516 20602 25544 21422
rect 25700 20641 25728 22066
rect 25686 20632 25742 20641
rect 25504 20596 25556 20602
rect 25686 20567 25742 20576
rect 25504 20538 25556 20544
rect 25792 20466 25820 23276
rect 25872 22024 25924 22030
rect 25872 21966 25924 21972
rect 25884 21554 25912 21966
rect 25872 21548 25924 21554
rect 25872 21490 25924 21496
rect 25872 21072 25924 21078
rect 25872 21014 25924 21020
rect 25688 20460 25740 20466
rect 25424 20420 25688 20448
rect 25424 19854 25452 20420
rect 25688 20402 25740 20408
rect 25780 20460 25832 20466
rect 25780 20402 25832 20408
rect 25504 20256 25556 20262
rect 25504 20198 25556 20204
rect 25516 19922 25544 20198
rect 25688 20052 25740 20058
rect 25688 19994 25740 20000
rect 25504 19916 25556 19922
rect 25504 19858 25556 19864
rect 25700 19854 25728 19994
rect 25412 19848 25464 19854
rect 25412 19790 25464 19796
rect 25688 19848 25740 19854
rect 25688 19790 25740 19796
rect 25884 17610 25912 21014
rect 25976 19786 26004 26250
rect 26068 26042 26096 27406
rect 26148 27396 26200 27402
rect 26148 27338 26200 27344
rect 26160 26926 26188 27338
rect 26344 27130 26372 27814
rect 26436 27402 26464 28358
rect 27436 27532 27488 27538
rect 27436 27474 27488 27480
rect 26792 27464 26844 27470
rect 26792 27406 26844 27412
rect 26424 27396 26476 27402
rect 26424 27338 26476 27344
rect 26332 27124 26384 27130
rect 26332 27066 26384 27072
rect 26148 26920 26200 26926
rect 26148 26862 26200 26868
rect 26332 26852 26384 26858
rect 26332 26794 26384 26800
rect 26240 26376 26292 26382
rect 26240 26318 26292 26324
rect 26056 26036 26108 26042
rect 26056 25978 26108 25984
rect 26068 24954 26096 25978
rect 26148 25220 26200 25226
rect 26148 25162 26200 25168
rect 26056 24948 26108 24954
rect 26056 24890 26108 24896
rect 26056 24676 26108 24682
rect 26056 24618 26108 24624
rect 26068 24324 26096 24618
rect 26160 24614 26188 25162
rect 26148 24608 26200 24614
rect 26148 24550 26200 24556
rect 26252 24410 26280 26318
rect 26344 25158 26372 26794
rect 26332 25152 26384 25158
rect 26332 25094 26384 25100
rect 26344 24886 26372 25094
rect 26332 24880 26384 24886
rect 26332 24822 26384 24828
rect 26240 24404 26292 24410
rect 26240 24346 26292 24352
rect 26148 24336 26200 24342
rect 26068 24296 26148 24324
rect 26148 24278 26200 24284
rect 26160 23662 26188 24278
rect 26148 23656 26200 23662
rect 26148 23598 26200 23604
rect 26344 23526 26372 24822
rect 26332 23520 26384 23526
rect 26332 23462 26384 23468
rect 26146 23352 26202 23361
rect 26146 23287 26202 23296
rect 26056 21344 26108 21350
rect 26056 21286 26108 21292
rect 25964 19780 26016 19786
rect 25964 19722 26016 19728
rect 25872 17604 25924 17610
rect 25872 17546 25924 17552
rect 25320 17332 25372 17338
rect 25320 17274 25372 17280
rect 25136 17196 25188 17202
rect 25136 17138 25188 17144
rect 25148 16182 25176 17138
rect 25688 17060 25740 17066
rect 25688 17002 25740 17008
rect 25136 16176 25188 16182
rect 25136 16118 25188 16124
rect 25320 16176 25372 16182
rect 25320 16118 25372 16124
rect 25148 15434 25176 16118
rect 25136 15428 25188 15434
rect 25136 15370 25188 15376
rect 25228 15360 25280 15366
rect 25228 15302 25280 15308
rect 25240 14958 25268 15302
rect 25332 15026 25360 16118
rect 25504 15904 25556 15910
rect 25504 15846 25556 15852
rect 25596 15904 25648 15910
rect 25596 15846 25648 15852
rect 25412 15632 25464 15638
rect 25412 15574 25464 15580
rect 25320 15020 25372 15026
rect 25320 14962 25372 14968
rect 25228 14952 25280 14958
rect 25228 14894 25280 14900
rect 25332 14550 25360 14962
rect 25320 14544 25372 14550
rect 25320 14486 25372 14492
rect 25320 14408 25372 14414
rect 25320 14350 25372 14356
rect 25332 14006 25360 14350
rect 25320 14000 25372 14006
rect 25320 13942 25372 13948
rect 25228 13932 25280 13938
rect 25228 13874 25280 13880
rect 25240 12986 25268 13874
rect 25320 13864 25372 13870
rect 25320 13806 25372 13812
rect 25332 13326 25360 13806
rect 25320 13320 25372 13326
rect 25320 13262 25372 13268
rect 25228 12980 25280 12986
rect 25228 12922 25280 12928
rect 25332 12850 25360 13262
rect 25320 12844 25372 12850
rect 25320 12786 25372 12792
rect 24964 11886 25084 11914
rect 24860 11348 24912 11354
rect 24860 11290 24912 11296
rect 24964 11257 24992 11886
rect 25044 11824 25096 11830
rect 25044 11766 25096 11772
rect 24950 11248 25006 11257
rect 24950 11183 25006 11192
rect 25056 11150 25084 11766
rect 25332 11762 25360 12786
rect 25320 11756 25372 11762
rect 25320 11698 25372 11704
rect 25136 11552 25188 11558
rect 25136 11494 25188 11500
rect 25148 11150 25176 11494
rect 25332 11150 25360 11698
rect 24768 11144 24820 11150
rect 24768 11086 24820 11092
rect 25044 11144 25096 11150
rect 25044 11086 25096 11092
rect 25136 11144 25188 11150
rect 25136 11086 25188 11092
rect 25320 11144 25372 11150
rect 25320 11086 25372 11092
rect 24780 10810 24808 11086
rect 24950 10840 25006 10849
rect 24768 10804 24820 10810
rect 24950 10775 25006 10784
rect 24768 10746 24820 10752
rect 24860 10532 24912 10538
rect 24860 10474 24912 10480
rect 24872 10130 24900 10474
rect 24964 10441 24992 10775
rect 24950 10432 25006 10441
rect 24950 10367 25006 10376
rect 25056 10130 25084 11086
rect 24860 10124 24912 10130
rect 24860 10066 24912 10072
rect 25044 10124 25096 10130
rect 25044 10066 25096 10072
rect 24872 9654 24900 10066
rect 25332 10062 25360 11086
rect 25424 10849 25452 15574
rect 25516 14414 25544 15846
rect 25608 15706 25636 15846
rect 25596 15700 25648 15706
rect 25596 15642 25648 15648
rect 25504 14408 25556 14414
rect 25504 14350 25556 14356
rect 25504 13796 25556 13802
rect 25504 13738 25556 13744
rect 25516 12918 25544 13738
rect 25504 12912 25556 12918
rect 25504 12854 25556 12860
rect 25516 11898 25544 12854
rect 25596 12844 25648 12850
rect 25596 12786 25648 12792
rect 25608 12442 25636 12786
rect 25596 12436 25648 12442
rect 25596 12378 25648 12384
rect 25504 11892 25556 11898
rect 25504 11834 25556 11840
rect 25700 11762 25728 17002
rect 25780 16516 25832 16522
rect 25780 16458 25832 16464
rect 25792 16250 25820 16458
rect 25780 16244 25832 16250
rect 25780 16186 25832 16192
rect 25964 16108 26016 16114
rect 25964 16050 26016 16056
rect 25780 16040 25832 16046
rect 25780 15982 25832 15988
rect 25792 14890 25820 15982
rect 25872 15496 25924 15502
rect 25872 15438 25924 15444
rect 25884 14890 25912 15438
rect 25780 14884 25832 14890
rect 25780 14826 25832 14832
rect 25872 14884 25924 14890
rect 25872 14826 25924 14832
rect 25792 14482 25820 14826
rect 25976 14498 26004 16050
rect 26068 15502 26096 21286
rect 26160 19786 26188 23287
rect 26240 22636 26292 22642
rect 26240 22578 26292 22584
rect 26252 22098 26280 22578
rect 26240 22092 26292 22098
rect 26240 22034 26292 22040
rect 26436 21418 26464 27338
rect 26804 26994 26832 27406
rect 26884 27328 26936 27334
rect 26884 27270 26936 27276
rect 26792 26988 26844 26994
rect 26792 26930 26844 26936
rect 26804 25906 26832 26930
rect 26792 25900 26844 25906
rect 26792 25842 26844 25848
rect 26896 25702 26924 27270
rect 27344 26988 27396 26994
rect 27344 26930 27396 26936
rect 27068 26852 27120 26858
rect 27068 26794 27120 26800
rect 27080 26586 27108 26794
rect 27068 26580 27120 26586
rect 27068 26522 27120 26528
rect 26976 26308 27028 26314
rect 26976 26250 27028 26256
rect 26884 25696 26936 25702
rect 26884 25638 26936 25644
rect 26896 25430 26924 25638
rect 26884 25424 26936 25430
rect 26884 25366 26936 25372
rect 26700 25288 26752 25294
rect 26700 25230 26752 25236
rect 26608 24608 26660 24614
rect 26608 24550 26660 24556
rect 26516 22024 26568 22030
rect 26516 21966 26568 21972
rect 26424 21412 26476 21418
rect 26424 21354 26476 21360
rect 26528 20890 26556 21966
rect 26436 20862 26556 20890
rect 26436 20058 26464 20862
rect 26424 20052 26476 20058
rect 26424 19994 26476 20000
rect 26436 19854 26464 19994
rect 26620 19938 26648 24550
rect 26712 21690 26740 25230
rect 26988 25226 27016 26250
rect 27252 25900 27304 25906
rect 27252 25842 27304 25848
rect 27160 25696 27212 25702
rect 27160 25638 27212 25644
rect 27172 25294 27200 25638
rect 27264 25498 27292 25842
rect 27252 25492 27304 25498
rect 27252 25434 27304 25440
rect 27160 25288 27212 25294
rect 27160 25230 27212 25236
rect 26976 25220 27028 25226
rect 26976 25162 27028 25168
rect 26988 24698 27016 25162
rect 26896 24670 27016 24698
rect 26896 23730 26924 24670
rect 27068 24608 27120 24614
rect 26988 24568 27068 24596
rect 26988 24410 27016 24568
rect 27068 24550 27120 24556
rect 27356 24410 27384 26930
rect 27448 26926 27476 27474
rect 27528 27396 27580 27402
rect 27528 27338 27580 27344
rect 27540 27130 27568 27338
rect 27528 27124 27580 27130
rect 27528 27066 27580 27072
rect 27528 26988 27580 26994
rect 27528 26930 27580 26936
rect 27436 26920 27488 26926
rect 27436 26862 27488 26868
rect 27448 25770 27476 26862
rect 27540 26314 27568 26930
rect 27632 26382 27660 28358
rect 27724 27130 27752 28426
rect 29012 28150 29040 28494
rect 29000 28144 29052 28150
rect 29000 28086 29052 28092
rect 27712 27124 27764 27130
rect 27712 27066 27764 27072
rect 27620 26376 27672 26382
rect 27620 26318 27672 26324
rect 27528 26308 27580 26314
rect 27528 26250 27580 26256
rect 27528 25900 27580 25906
rect 27528 25842 27580 25848
rect 27436 25764 27488 25770
rect 27436 25706 27488 25712
rect 26976 24404 27028 24410
rect 26976 24346 27028 24352
rect 27344 24404 27396 24410
rect 27344 24346 27396 24352
rect 26884 23724 26936 23730
rect 26884 23666 26936 23672
rect 26792 22568 26844 22574
rect 26792 22510 26844 22516
rect 26700 21684 26752 21690
rect 26700 21626 26752 21632
rect 26804 21010 26832 22510
rect 26792 21004 26844 21010
rect 26792 20946 26844 20952
rect 26896 20330 26924 23666
rect 26988 23594 27016 24346
rect 27252 24132 27304 24138
rect 27252 24074 27304 24080
rect 27264 23798 27292 24074
rect 27252 23792 27304 23798
rect 27252 23734 27304 23740
rect 26976 23588 27028 23594
rect 26976 23530 27028 23536
rect 26988 23186 27016 23530
rect 26976 23180 27028 23186
rect 26976 23122 27028 23128
rect 26988 22574 27016 23122
rect 26976 22568 27028 22574
rect 26976 22510 27028 22516
rect 27356 21962 27384 24346
rect 27448 24342 27476 25706
rect 27540 25498 27568 25842
rect 27528 25492 27580 25498
rect 27528 25434 27580 25440
rect 29000 24812 29052 24818
rect 29000 24754 29052 24760
rect 28816 24608 28868 24614
rect 28816 24550 28868 24556
rect 27436 24336 27488 24342
rect 27436 24278 27488 24284
rect 27804 24200 27856 24206
rect 27804 24142 27856 24148
rect 27816 23866 27844 24142
rect 28356 24064 28408 24070
rect 28356 24006 28408 24012
rect 27804 23860 27856 23866
rect 27804 23802 27856 23808
rect 28368 23118 28396 24006
rect 28828 23798 28856 24550
rect 29012 24206 29040 24754
rect 29000 24200 29052 24206
rect 29000 24142 29052 24148
rect 29104 23866 29132 29106
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 65654 28860 65962 28869
rect 65654 28858 65660 28860
rect 65716 28858 65740 28860
rect 65796 28858 65820 28860
rect 65876 28858 65900 28860
rect 65956 28858 65962 28860
rect 65716 28806 65718 28858
rect 65898 28806 65900 28858
rect 65654 28804 65660 28806
rect 65716 28804 65740 28806
rect 65796 28804 65820 28806
rect 65876 28804 65900 28806
rect 65956 28804 65962 28806
rect 65654 28795 65962 28804
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 30288 28144 30340 28150
rect 30288 28086 30340 28092
rect 29184 28076 29236 28082
rect 29184 28018 29236 28024
rect 29196 27606 29224 28018
rect 29276 27872 29328 27878
rect 29276 27814 29328 27820
rect 29184 27600 29236 27606
rect 29184 27542 29236 27548
rect 29288 27010 29316 27814
rect 29196 26994 29316 27010
rect 29184 26988 29316 26994
rect 29236 26982 29316 26988
rect 29184 26930 29236 26936
rect 29092 23860 29144 23866
rect 29092 23802 29144 23808
rect 28816 23792 28868 23798
rect 28816 23734 28868 23740
rect 28356 23112 28408 23118
rect 28356 23054 28408 23060
rect 28908 23112 28960 23118
rect 28908 23054 28960 23060
rect 28080 23044 28132 23050
rect 28080 22986 28132 22992
rect 28092 22778 28120 22986
rect 28080 22772 28132 22778
rect 28080 22714 28132 22720
rect 28920 22710 28948 23054
rect 29000 22976 29052 22982
rect 29000 22918 29052 22924
rect 29012 22710 29040 22918
rect 28908 22704 28960 22710
rect 28908 22646 28960 22652
rect 29000 22704 29052 22710
rect 29000 22646 29052 22652
rect 27436 22636 27488 22642
rect 27436 22578 27488 22584
rect 27804 22636 27856 22642
rect 27804 22578 27856 22584
rect 27448 22522 27476 22578
rect 27448 22494 27568 22522
rect 27344 21956 27396 21962
rect 27344 21898 27396 21904
rect 27540 21554 27568 22494
rect 27816 22234 27844 22578
rect 27804 22228 27856 22234
rect 27804 22170 27856 22176
rect 28540 22160 28592 22166
rect 28540 22102 28592 22108
rect 28080 21888 28132 21894
rect 28080 21830 28132 21836
rect 27528 21548 27580 21554
rect 27528 21490 27580 21496
rect 27712 21480 27764 21486
rect 27712 21422 27764 21428
rect 27436 21412 27488 21418
rect 27436 21354 27488 21360
rect 27068 21344 27120 21350
rect 27068 21286 27120 21292
rect 27080 20942 27108 21286
rect 27068 20936 27120 20942
rect 27068 20878 27120 20884
rect 27344 20936 27396 20942
rect 27344 20878 27396 20884
rect 26884 20324 26936 20330
rect 26884 20266 26936 20272
rect 26528 19910 26648 19938
rect 26424 19848 26476 19854
rect 26424 19790 26476 19796
rect 26148 19780 26200 19786
rect 26148 19722 26200 19728
rect 26160 19514 26188 19722
rect 26148 19508 26200 19514
rect 26148 19450 26200 19456
rect 26330 18456 26386 18465
rect 26330 18391 26386 18400
rect 26344 18290 26372 18391
rect 26332 18284 26384 18290
rect 26332 18226 26384 18232
rect 26528 18057 26556 19910
rect 26608 19848 26660 19854
rect 26608 19790 26660 19796
rect 26620 18970 26648 19790
rect 27068 19712 27120 19718
rect 27068 19654 27120 19660
rect 27080 19378 27108 19654
rect 26976 19372 27028 19378
rect 26976 19314 27028 19320
rect 27068 19372 27120 19378
rect 27068 19314 27120 19320
rect 26608 18964 26660 18970
rect 26608 18906 26660 18912
rect 26988 18834 27016 19314
rect 26976 18828 27028 18834
rect 26976 18770 27028 18776
rect 26514 18048 26570 18057
rect 26514 17983 26570 17992
rect 26988 17882 27016 18770
rect 26976 17876 27028 17882
rect 26976 17818 27028 17824
rect 27356 17728 27384 20878
rect 27448 19922 27476 21354
rect 27724 20602 27752 21422
rect 28092 20806 28120 21830
rect 28552 21554 28580 22102
rect 28920 21690 28948 22646
rect 29092 22636 29144 22642
rect 29092 22578 29144 22584
rect 29000 22432 29052 22438
rect 29000 22374 29052 22380
rect 28908 21684 28960 21690
rect 28908 21626 28960 21632
rect 28540 21548 28592 21554
rect 28540 21490 28592 21496
rect 28724 21548 28776 21554
rect 28724 21490 28776 21496
rect 28736 21026 28764 21490
rect 28540 21004 28592 21010
rect 28736 20998 28856 21026
rect 28540 20946 28592 20952
rect 28080 20800 28132 20806
rect 28080 20742 28132 20748
rect 28264 20800 28316 20806
rect 28264 20742 28316 20748
rect 27712 20596 27764 20602
rect 27712 20538 27764 20544
rect 28276 20398 28304 20742
rect 28552 20602 28580 20946
rect 28828 20942 28856 20998
rect 28816 20936 28868 20942
rect 28816 20878 28868 20884
rect 28540 20596 28592 20602
rect 28540 20538 28592 20544
rect 28264 20392 28316 20398
rect 28264 20334 28316 20340
rect 27528 20052 27580 20058
rect 27528 19994 27580 20000
rect 27436 19916 27488 19922
rect 27436 19858 27488 19864
rect 27540 19854 27568 19994
rect 27528 19848 27580 19854
rect 27528 19790 27580 19796
rect 28172 18624 28224 18630
rect 28172 18566 28224 18572
rect 28184 18222 28212 18566
rect 27620 18216 27672 18222
rect 27620 18158 27672 18164
rect 28172 18216 28224 18222
rect 28172 18158 28224 18164
rect 27264 17700 27384 17728
rect 27264 17610 27292 17700
rect 27068 17604 27120 17610
rect 27068 17546 27120 17552
rect 27252 17604 27304 17610
rect 27252 17546 27304 17552
rect 27344 17604 27396 17610
rect 27344 17546 27396 17552
rect 26516 17536 26568 17542
rect 26516 17478 26568 17484
rect 26608 17536 26660 17542
rect 26608 17478 26660 17484
rect 26528 17270 26556 17478
rect 26516 17264 26568 17270
rect 26514 17232 26516 17241
rect 26568 17232 26570 17241
rect 26514 17167 26570 17176
rect 26620 17066 26648 17478
rect 26608 17060 26660 17066
rect 26608 17002 26660 17008
rect 26792 17060 26844 17066
rect 26792 17002 26844 17008
rect 26240 16992 26292 16998
rect 26240 16934 26292 16940
rect 26252 16114 26280 16934
rect 26332 16448 26384 16454
rect 26332 16390 26384 16396
rect 26344 16289 26372 16390
rect 26330 16280 26386 16289
rect 26330 16215 26386 16224
rect 26344 16182 26372 16215
rect 26332 16176 26384 16182
rect 26332 16118 26384 16124
rect 26804 16114 26832 17002
rect 26240 16108 26292 16114
rect 26240 16050 26292 16056
rect 26792 16108 26844 16114
rect 26792 16050 26844 16056
rect 26056 15496 26108 15502
rect 26056 15438 26108 15444
rect 26240 15020 26292 15026
rect 26240 14962 26292 14968
rect 25780 14476 25832 14482
rect 25780 14418 25832 14424
rect 25884 14470 26004 14498
rect 25780 13796 25832 13802
rect 25780 13738 25832 13744
rect 25792 12646 25820 13738
rect 25884 12866 25912 14470
rect 26252 14346 26280 14962
rect 26240 14340 26292 14346
rect 26240 14282 26292 14288
rect 27080 13938 27108 17546
rect 27356 17338 27384 17546
rect 27344 17332 27396 17338
rect 27344 17274 27396 17280
rect 27528 17196 27580 17202
rect 27528 17138 27580 17144
rect 27250 16552 27306 16561
rect 27250 16487 27306 16496
rect 27160 15496 27212 15502
rect 27160 15438 27212 15444
rect 27068 13932 27120 13938
rect 26896 13892 27068 13920
rect 26148 13524 26200 13530
rect 26148 13466 26200 13472
rect 26056 13252 26108 13258
rect 26056 13194 26108 13200
rect 26068 12986 26096 13194
rect 26056 12980 26108 12986
rect 26056 12922 26108 12928
rect 25884 12838 26096 12866
rect 25780 12640 25832 12646
rect 25780 12582 25832 12588
rect 25872 12436 25924 12442
rect 25872 12378 25924 12384
rect 25884 12102 25912 12378
rect 25872 12096 25924 12102
rect 25872 12038 25924 12044
rect 25504 11756 25556 11762
rect 25504 11698 25556 11704
rect 25688 11756 25740 11762
rect 25688 11698 25740 11704
rect 25410 10840 25466 10849
rect 25516 10810 25544 11698
rect 25700 11354 25728 11698
rect 25596 11348 25648 11354
rect 25596 11290 25648 11296
rect 25688 11348 25740 11354
rect 25688 11290 25740 11296
rect 25410 10775 25466 10784
rect 25504 10804 25556 10810
rect 25504 10746 25556 10752
rect 25412 10668 25464 10674
rect 25412 10610 25464 10616
rect 25424 10266 25452 10610
rect 25412 10260 25464 10266
rect 25412 10202 25464 10208
rect 25320 10056 25372 10062
rect 25320 9998 25372 10004
rect 25424 9654 25452 10202
rect 24860 9648 24912 9654
rect 24860 9590 24912 9596
rect 25412 9648 25464 9654
rect 25412 9590 25464 9596
rect 24584 9580 24636 9586
rect 24584 9522 24636 9528
rect 24490 9208 24546 9217
rect 24596 9178 24624 9522
rect 24490 9143 24546 9152
rect 24584 9172 24636 9178
rect 24584 9114 24636 9120
rect 24400 8900 24452 8906
rect 24400 8842 24452 8848
rect 24308 8628 24360 8634
rect 24308 8570 24360 8576
rect 24214 8392 24270 8401
rect 24214 8327 24270 8336
rect 23756 8084 23808 8090
rect 23756 8026 23808 8032
rect 24412 7886 24440 8842
rect 24872 8566 24900 9590
rect 25320 9580 25372 9586
rect 25320 9522 25372 9528
rect 25332 9178 25360 9522
rect 25608 9518 25636 11290
rect 25596 9512 25648 9518
rect 25596 9454 25648 9460
rect 25320 9172 25372 9178
rect 25320 9114 25372 9120
rect 25608 8906 25636 9454
rect 25596 8900 25648 8906
rect 25596 8842 25648 8848
rect 24860 8560 24912 8566
rect 24860 8502 24912 8508
rect 25044 8424 25096 8430
rect 25044 8366 25096 8372
rect 24952 7948 25004 7954
rect 24952 7890 25004 7896
rect 23572 7880 23624 7886
rect 23572 7822 23624 7828
rect 24400 7880 24452 7886
rect 24400 7822 24452 7828
rect 23584 7546 23612 7822
rect 23664 7812 23716 7818
rect 23664 7754 23716 7760
rect 23572 7540 23624 7546
rect 23572 7482 23624 7488
rect 23676 7478 23704 7754
rect 24860 7744 24912 7750
rect 24860 7686 24912 7692
rect 23664 7472 23716 7478
rect 23664 7414 23716 7420
rect 23676 6458 23704 7414
rect 24872 7410 24900 7686
rect 24964 7546 24992 7890
rect 24952 7540 25004 7546
rect 24952 7482 25004 7488
rect 24860 7404 24912 7410
rect 24860 7346 24912 7352
rect 25056 7342 25084 8366
rect 25608 8022 25636 8842
rect 26068 8022 26096 12838
rect 26160 11506 26188 13466
rect 26240 13320 26292 13326
rect 26240 13262 26292 13268
rect 26252 12102 26280 13262
rect 26792 13184 26844 13190
rect 26792 13126 26844 13132
rect 26332 12776 26384 12782
rect 26332 12718 26384 12724
rect 26240 12096 26292 12102
rect 26240 12038 26292 12044
rect 26160 11478 26280 11506
rect 26148 11348 26200 11354
rect 26148 11290 26200 11296
rect 26160 10674 26188 11290
rect 26252 10810 26280 11478
rect 26240 10804 26292 10810
rect 26240 10746 26292 10752
rect 26148 10668 26200 10674
rect 26148 10610 26200 10616
rect 26344 10554 26372 12718
rect 26516 12096 26568 12102
rect 26516 12038 26568 12044
rect 26528 11694 26556 12038
rect 26804 11898 26832 13126
rect 26896 12850 26924 13892
rect 27068 13874 27120 13880
rect 27172 12986 27200 15438
rect 27264 15434 27292 16487
rect 27344 16448 27396 16454
rect 27344 16390 27396 16396
rect 27356 15706 27384 16390
rect 27344 15700 27396 15706
rect 27344 15642 27396 15648
rect 27252 15428 27304 15434
rect 27252 15370 27304 15376
rect 27264 14550 27292 15370
rect 27252 14544 27304 14550
rect 27252 14486 27304 14492
rect 27344 14272 27396 14278
rect 27344 14214 27396 14220
rect 27252 13184 27304 13190
rect 27252 13126 27304 13132
rect 27160 12980 27212 12986
rect 27160 12922 27212 12928
rect 27264 12918 27292 13126
rect 27252 12912 27304 12918
rect 27252 12854 27304 12860
rect 26884 12844 26936 12850
rect 26884 12786 26936 12792
rect 26976 12844 27028 12850
rect 26976 12786 27028 12792
rect 26988 12238 27016 12786
rect 26976 12232 27028 12238
rect 26976 12174 27028 12180
rect 26792 11892 26844 11898
rect 26792 11834 26844 11840
rect 26976 11756 27028 11762
rect 26976 11698 27028 11704
rect 26516 11688 26568 11694
rect 26988 11665 27016 11698
rect 27068 11688 27120 11694
rect 26516 11630 26568 11636
rect 26974 11656 27030 11665
rect 26528 11150 26556 11630
rect 27068 11630 27120 11636
rect 26974 11591 27030 11600
rect 26608 11552 26660 11558
rect 26608 11494 26660 11500
rect 26620 11150 26648 11494
rect 26516 11144 26568 11150
rect 26516 11086 26568 11092
rect 26608 11144 26660 11150
rect 26608 11086 26660 11092
rect 26160 10526 26372 10554
rect 26160 10470 26188 10526
rect 26148 10464 26200 10470
rect 26148 10406 26200 10412
rect 26160 8498 26188 10406
rect 26332 10056 26384 10062
rect 26332 9998 26384 10004
rect 26344 9654 26372 9998
rect 26528 9654 26556 11086
rect 26608 10804 26660 10810
rect 26608 10746 26660 10752
rect 26620 10062 26648 10746
rect 26608 10056 26660 10062
rect 26608 9998 26660 10004
rect 26792 9920 26844 9926
rect 26792 9862 26844 9868
rect 26332 9648 26384 9654
rect 26332 9590 26384 9596
rect 26516 9648 26568 9654
rect 26516 9590 26568 9596
rect 26804 8974 26832 9862
rect 26792 8968 26844 8974
rect 26792 8910 26844 8916
rect 26148 8492 26200 8498
rect 26148 8434 26200 8440
rect 26700 8424 26752 8430
rect 26700 8366 26752 8372
rect 25596 8016 25648 8022
rect 25596 7958 25648 7964
rect 26056 8016 26108 8022
rect 26056 7958 26108 7964
rect 26712 7886 26740 8366
rect 27080 8090 27108 11630
rect 27356 11558 27384 14214
rect 27540 11898 27568 17138
rect 27632 12646 27660 18158
rect 27988 17876 28040 17882
rect 27988 17818 28040 17824
rect 28000 17542 28028 17818
rect 27988 17536 28040 17542
rect 27988 17478 28040 17484
rect 27712 17332 27764 17338
rect 27804 17332 27856 17338
rect 27764 17292 27804 17320
rect 27712 17274 27764 17280
rect 27804 17274 27856 17280
rect 27724 16046 27752 17274
rect 27896 17264 27948 17270
rect 27816 17212 27896 17218
rect 27816 17206 27948 17212
rect 27816 17202 27936 17206
rect 27804 17196 27936 17202
rect 27856 17190 27936 17196
rect 27804 17138 27856 17144
rect 28172 16584 28224 16590
rect 28172 16526 28224 16532
rect 27712 16040 27764 16046
rect 27712 15982 27764 15988
rect 28184 15502 28212 16526
rect 28172 15496 28224 15502
rect 28172 15438 28224 15444
rect 28080 15360 28132 15366
rect 28080 15302 28132 15308
rect 27988 14408 28040 14414
rect 27988 14350 28040 14356
rect 27712 14340 27764 14346
rect 27712 14282 27764 14288
rect 27724 14249 27752 14282
rect 27710 14240 27766 14249
rect 27710 14175 27766 14184
rect 28000 13938 28028 14350
rect 27988 13932 28040 13938
rect 27988 13874 28040 13880
rect 27896 13864 27948 13870
rect 27896 13806 27948 13812
rect 27908 13433 27936 13806
rect 27894 13424 27950 13433
rect 27894 13359 27950 13368
rect 27712 12980 27764 12986
rect 27712 12922 27764 12928
rect 27620 12640 27672 12646
rect 27620 12582 27672 12588
rect 27632 12374 27660 12582
rect 27620 12368 27672 12374
rect 27620 12310 27672 12316
rect 27620 12164 27672 12170
rect 27724 12152 27752 12922
rect 27804 12912 27856 12918
rect 27804 12854 27856 12860
rect 27672 12124 27752 12152
rect 27620 12106 27672 12112
rect 27528 11892 27580 11898
rect 27528 11834 27580 11840
rect 27344 11552 27396 11558
rect 27344 11494 27396 11500
rect 27528 10056 27580 10062
rect 27448 10004 27528 10010
rect 27448 9998 27580 10004
rect 27448 9982 27568 9998
rect 27448 9586 27476 9982
rect 27436 9580 27488 9586
rect 27436 9522 27488 9528
rect 27448 9178 27476 9522
rect 27436 9172 27488 9178
rect 27436 9114 27488 9120
rect 27160 8492 27212 8498
rect 27160 8434 27212 8440
rect 27068 8084 27120 8090
rect 27068 8026 27120 8032
rect 25780 7880 25832 7886
rect 25780 7822 25832 7828
rect 25964 7880 26016 7886
rect 25964 7822 26016 7828
rect 26700 7880 26752 7886
rect 26700 7822 26752 7828
rect 25596 7744 25648 7750
rect 25596 7686 25648 7692
rect 25320 7404 25372 7410
rect 25320 7346 25372 7352
rect 25044 7336 25096 7342
rect 25044 7278 25096 7284
rect 23848 7200 23900 7206
rect 23848 7142 23900 7148
rect 23756 6656 23808 6662
rect 23756 6598 23808 6604
rect 23664 6452 23716 6458
rect 23664 6394 23716 6400
rect 23480 5908 23532 5914
rect 23480 5850 23532 5856
rect 23388 5704 23440 5710
rect 23388 5646 23440 5652
rect 23296 5636 23348 5642
rect 23296 5578 23348 5584
rect 23020 5568 23072 5574
rect 23020 5510 23072 5516
rect 22744 5228 22796 5234
rect 22744 5170 22796 5176
rect 22756 5030 22784 5170
rect 22744 5024 22796 5030
rect 22744 4966 22796 4972
rect 22100 4820 22152 4826
rect 22100 4762 22152 4768
rect 22756 4758 22784 4966
rect 22744 4752 22796 4758
rect 22744 4694 22796 4700
rect 22376 3936 22428 3942
rect 22376 3878 22428 3884
rect 22008 3188 22060 3194
rect 22008 3130 22060 3136
rect 21824 2984 21876 2990
rect 21824 2926 21876 2932
rect 21272 2848 21324 2854
rect 21272 2790 21324 2796
rect 21284 800 21312 2790
rect 21548 2576 21600 2582
rect 21548 2518 21600 2524
rect 21560 800 21588 2518
rect 21836 800 21864 2926
rect 22020 2922 22048 3130
rect 22008 2916 22060 2922
rect 22008 2858 22060 2864
rect 22100 2508 22152 2514
rect 22100 2450 22152 2456
rect 22112 800 22140 2450
rect 22388 800 22416 3878
rect 22652 3664 22704 3670
rect 22652 3606 22704 3612
rect 22664 800 22692 3606
rect 22756 2038 22784 4694
rect 23032 4622 23060 5510
rect 23308 5370 23336 5578
rect 23296 5364 23348 5370
rect 23296 5306 23348 5312
rect 23400 5166 23428 5646
rect 23388 5160 23440 5166
rect 23388 5102 23440 5108
rect 23204 5092 23256 5098
rect 23204 5034 23256 5040
rect 23020 4616 23072 4622
rect 23020 4558 23072 4564
rect 23032 3466 23060 4558
rect 23216 4146 23244 5034
rect 23400 4282 23428 5102
rect 23492 4622 23520 5850
rect 23768 5352 23796 6598
rect 23860 6322 23888 7142
rect 25056 6934 25084 7278
rect 25332 7206 25360 7346
rect 25320 7200 25372 7206
rect 25320 7142 25372 7148
rect 25044 6928 25096 6934
rect 25044 6870 25096 6876
rect 25608 6730 25636 7686
rect 25792 7410 25820 7822
rect 25780 7404 25832 7410
rect 25780 7346 25832 7352
rect 25596 6724 25648 6730
rect 25596 6666 25648 6672
rect 25044 6656 25096 6662
rect 25044 6598 25096 6604
rect 25056 6458 25084 6598
rect 25044 6452 25096 6458
rect 25044 6394 25096 6400
rect 23848 6316 23900 6322
rect 23848 6258 23900 6264
rect 24676 5704 24728 5710
rect 24676 5646 24728 5652
rect 23676 5324 23796 5352
rect 23480 4616 23532 4622
rect 23480 4558 23532 4564
rect 23388 4276 23440 4282
rect 23388 4218 23440 4224
rect 23676 4146 23704 5324
rect 24688 5302 24716 5646
rect 25044 5636 25096 5642
rect 25044 5578 25096 5584
rect 25596 5636 25648 5642
rect 25596 5578 25648 5584
rect 24768 5568 24820 5574
rect 24768 5510 24820 5516
rect 24676 5296 24728 5302
rect 24676 5238 24728 5244
rect 24780 5234 24808 5510
rect 25056 5302 25084 5578
rect 25044 5296 25096 5302
rect 25044 5238 25096 5244
rect 23756 5226 23808 5232
rect 23756 5168 23808 5174
rect 24584 5228 24636 5234
rect 24584 5170 24636 5176
rect 24768 5228 24820 5234
rect 24768 5170 24820 5176
rect 24952 5228 25004 5234
rect 24952 5170 25004 5176
rect 23768 4826 23796 5168
rect 23756 4820 23808 4826
rect 23756 4762 23808 4768
rect 24308 4684 24360 4690
rect 24308 4626 24360 4632
rect 24320 4146 24348 4626
rect 23204 4140 23256 4146
rect 23204 4082 23256 4088
rect 23664 4140 23716 4146
rect 23664 4082 23716 4088
rect 24308 4140 24360 4146
rect 24308 4082 24360 4088
rect 23112 4072 23164 4078
rect 23112 4014 23164 4020
rect 23124 3738 23152 4014
rect 23112 3732 23164 3738
rect 23112 3674 23164 3680
rect 24596 3602 24624 5170
rect 24964 4554 24992 5170
rect 25228 5024 25280 5030
rect 25228 4966 25280 4972
rect 25240 4622 25268 4966
rect 25608 4758 25636 5578
rect 25596 4752 25648 4758
rect 25596 4694 25648 4700
rect 25228 4616 25280 4622
rect 25228 4558 25280 4564
rect 24952 4548 25004 4554
rect 24952 4490 25004 4496
rect 25976 4010 26004 7822
rect 26240 7744 26292 7750
rect 26240 7686 26292 7692
rect 26252 6798 26280 7686
rect 26332 7200 26384 7206
rect 26332 7142 26384 7148
rect 26424 7200 26476 7206
rect 26424 7142 26476 7148
rect 26240 6792 26292 6798
rect 26240 6734 26292 6740
rect 26252 6186 26280 6734
rect 26344 6390 26372 7142
rect 26436 6798 26464 7142
rect 26424 6792 26476 6798
rect 26424 6734 26476 6740
rect 26792 6792 26844 6798
rect 26792 6734 26844 6740
rect 26804 6458 26832 6734
rect 27068 6656 27120 6662
rect 27068 6598 27120 6604
rect 26792 6452 26844 6458
rect 26792 6394 26844 6400
rect 27080 6390 27108 6598
rect 26332 6384 26384 6390
rect 26332 6326 26384 6332
rect 27068 6384 27120 6390
rect 27068 6326 27120 6332
rect 26240 6180 26292 6186
rect 26240 6122 26292 6128
rect 26344 5914 26372 6326
rect 26332 5908 26384 5914
rect 26332 5850 26384 5856
rect 26424 5840 26476 5846
rect 26424 5782 26476 5788
rect 26436 5642 26464 5782
rect 27172 5642 27200 8434
rect 27528 7948 27580 7954
rect 27528 7890 27580 7896
rect 27540 7478 27568 7890
rect 27528 7472 27580 7478
rect 27528 7414 27580 7420
rect 27344 7404 27396 7410
rect 27344 7346 27396 7352
rect 26424 5636 26476 5642
rect 26424 5578 26476 5584
rect 27160 5636 27212 5642
rect 27160 5578 27212 5584
rect 25964 4004 26016 4010
rect 25964 3946 26016 3952
rect 24584 3596 24636 3602
rect 24584 3538 24636 3544
rect 23204 3528 23256 3534
rect 23204 3470 23256 3476
rect 24860 3528 24912 3534
rect 24860 3470 24912 3476
rect 25688 3528 25740 3534
rect 25688 3470 25740 3476
rect 23020 3460 23072 3466
rect 23020 3402 23072 3408
rect 22928 2440 22980 2446
rect 22928 2382 22980 2388
rect 22744 2032 22796 2038
rect 22744 1974 22796 1980
rect 22940 800 22968 2382
rect 23216 800 23244 3470
rect 23480 2916 23532 2922
rect 23480 2858 23532 2864
rect 23492 800 23520 2858
rect 23756 2848 23808 2854
rect 23756 2790 23808 2796
rect 24308 2848 24360 2854
rect 24308 2790 24360 2796
rect 23768 800 23796 2790
rect 24032 2576 24084 2582
rect 24032 2518 24084 2524
rect 24044 800 24072 2518
rect 24320 800 24348 2790
rect 24584 2508 24636 2514
rect 24584 2450 24636 2456
rect 24596 800 24624 2450
rect 24872 800 24900 3470
rect 25136 2984 25188 2990
rect 25136 2926 25188 2932
rect 25148 800 25176 2926
rect 25412 2440 25464 2446
rect 25412 2382 25464 2388
rect 25424 800 25452 2382
rect 25700 800 25728 3470
rect 25976 3466 26004 3946
rect 26332 3936 26384 3942
rect 26332 3878 26384 3884
rect 26240 3528 26292 3534
rect 26240 3470 26292 3476
rect 25964 3460 26016 3466
rect 25964 3402 26016 3408
rect 25964 2916 26016 2922
rect 25964 2858 26016 2864
rect 25976 800 26004 2858
rect 26252 800 26280 3470
rect 26344 2961 26372 3878
rect 26436 3194 26464 5578
rect 26792 5160 26844 5166
rect 26792 5102 26844 5108
rect 26700 5024 26752 5030
rect 26700 4966 26752 4972
rect 26712 3534 26740 4966
rect 26804 4214 26832 5102
rect 27172 4826 27200 5578
rect 27252 5228 27304 5234
rect 27356 5216 27384 7346
rect 27632 6322 27660 12106
rect 27816 11558 27844 12854
rect 28000 12850 28028 13874
rect 28092 13734 28120 15302
rect 28184 14550 28212 15438
rect 28172 14544 28224 14550
rect 28172 14486 28224 14492
rect 28276 13938 28304 20334
rect 28540 19848 28592 19854
rect 28540 19790 28592 19796
rect 28552 19514 28580 19790
rect 28540 19508 28592 19514
rect 28540 19450 28592 19456
rect 28356 19168 28408 19174
rect 28356 19110 28408 19116
rect 28368 18766 28396 19110
rect 28828 18850 28856 20878
rect 29012 20874 29040 22374
rect 29104 21146 29132 22578
rect 29196 22438 29224 26930
rect 30300 26450 30328 28086
rect 67638 27976 67694 27985
rect 67638 27911 67640 27920
rect 67692 27911 67694 27920
rect 67640 27882 67692 27888
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 65654 27772 65962 27781
rect 65654 27770 65660 27772
rect 65716 27770 65740 27772
rect 65796 27770 65820 27772
rect 65876 27770 65900 27772
rect 65956 27770 65962 27772
rect 65716 27718 65718 27770
rect 65898 27718 65900 27770
rect 65654 27716 65660 27718
rect 65716 27716 65740 27718
rect 65796 27716 65820 27718
rect 65876 27716 65900 27718
rect 65956 27716 65962 27718
rect 65654 27707 65962 27716
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 67640 26784 67692 26790
rect 67640 26726 67692 26732
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 65654 26684 65962 26693
rect 65654 26682 65660 26684
rect 65716 26682 65740 26684
rect 65796 26682 65820 26684
rect 65876 26682 65900 26684
rect 65956 26682 65962 26684
rect 65716 26630 65718 26682
rect 65898 26630 65900 26682
rect 65654 26628 65660 26630
rect 65716 26628 65740 26630
rect 65796 26628 65820 26630
rect 65876 26628 65900 26630
rect 65956 26628 65962 26630
rect 65654 26619 65962 26628
rect 67652 26625 67680 26726
rect 67638 26616 67694 26625
rect 67638 26551 67694 26560
rect 30288 26444 30340 26450
rect 30288 26386 30340 26392
rect 30300 26042 30328 26386
rect 30748 26308 30800 26314
rect 30748 26250 30800 26256
rect 30760 26042 30788 26250
rect 31576 26240 31628 26246
rect 31576 26182 31628 26188
rect 30288 26036 30340 26042
rect 30288 25978 30340 25984
rect 30748 26036 30800 26042
rect 30748 25978 30800 25984
rect 31588 25974 31616 26182
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 31576 25968 31628 25974
rect 31576 25910 31628 25916
rect 30104 25900 30156 25906
rect 30104 25842 30156 25848
rect 30288 25900 30340 25906
rect 30288 25842 30340 25848
rect 30564 25900 30616 25906
rect 30564 25842 30616 25848
rect 31024 25900 31076 25906
rect 31024 25842 31076 25848
rect 29828 25764 29880 25770
rect 29828 25706 29880 25712
rect 29460 25288 29512 25294
rect 29460 25230 29512 25236
rect 29472 24818 29500 25230
rect 29840 24886 29868 25706
rect 30116 25294 30144 25842
rect 30300 25702 30328 25842
rect 30288 25696 30340 25702
rect 30288 25638 30340 25644
rect 30576 25498 30604 25842
rect 30564 25492 30616 25498
rect 30564 25434 30616 25440
rect 30104 25288 30156 25294
rect 30104 25230 30156 25236
rect 31036 24886 31064 25842
rect 31392 25220 31444 25226
rect 31392 25162 31444 25168
rect 31116 25152 31168 25158
rect 31116 25094 31168 25100
rect 31128 24954 31156 25094
rect 31116 24948 31168 24954
rect 31116 24890 31168 24896
rect 29828 24880 29880 24886
rect 29828 24822 29880 24828
rect 31024 24880 31076 24886
rect 31024 24822 31076 24828
rect 29460 24812 29512 24818
rect 29460 24754 29512 24760
rect 29472 24206 29500 24754
rect 29460 24200 29512 24206
rect 29460 24142 29512 24148
rect 29276 23860 29328 23866
rect 29276 23802 29328 23808
rect 29184 22432 29236 22438
rect 29184 22374 29236 22380
rect 29092 21140 29144 21146
rect 29092 21082 29144 21088
rect 29000 20868 29052 20874
rect 29000 20810 29052 20816
rect 29000 20460 29052 20466
rect 29000 20402 29052 20408
rect 29012 19990 29040 20402
rect 29000 19984 29052 19990
rect 29000 19926 29052 19932
rect 28828 18822 28948 18850
rect 28356 18760 28408 18766
rect 28356 18702 28408 18708
rect 28816 18760 28868 18766
rect 28816 18702 28868 18708
rect 28368 14414 28396 18702
rect 28828 18630 28856 18702
rect 28816 18624 28868 18630
rect 28816 18566 28868 18572
rect 28828 18426 28856 18566
rect 28724 18420 28776 18426
rect 28724 18362 28776 18368
rect 28816 18420 28868 18426
rect 28816 18362 28868 18368
rect 28448 18352 28500 18358
rect 28448 18294 28500 18300
rect 28460 18154 28488 18294
rect 28736 18222 28764 18362
rect 28724 18216 28776 18222
rect 28724 18158 28776 18164
rect 28448 18148 28500 18154
rect 28448 18090 28500 18096
rect 28632 17264 28684 17270
rect 28630 17232 28632 17241
rect 28684 17232 28686 17241
rect 28630 17167 28686 17176
rect 28920 17134 28948 18822
rect 29012 18630 29040 19926
rect 29104 19854 29132 21082
rect 29288 20466 29316 23802
rect 29472 22506 29500 24142
rect 29840 23186 29868 24822
rect 30012 24812 30064 24818
rect 30012 24754 30064 24760
rect 30024 23526 30052 24754
rect 31036 23730 31064 24822
rect 31404 24206 31432 25162
rect 31392 24200 31444 24206
rect 31392 24142 31444 24148
rect 31208 24064 31260 24070
rect 31208 24006 31260 24012
rect 31220 23866 31248 24006
rect 31208 23860 31260 23866
rect 31208 23802 31260 23808
rect 31024 23724 31076 23730
rect 31024 23666 31076 23672
rect 31300 23724 31352 23730
rect 31300 23666 31352 23672
rect 30012 23520 30064 23526
rect 30012 23462 30064 23468
rect 30656 23520 30708 23526
rect 30656 23462 30708 23468
rect 29828 23180 29880 23186
rect 29828 23122 29880 23128
rect 29920 23112 29972 23118
rect 29920 23054 29972 23060
rect 29552 22704 29604 22710
rect 29552 22646 29604 22652
rect 29460 22500 29512 22506
rect 29460 22442 29512 22448
rect 29276 20460 29328 20466
rect 29276 20402 29328 20408
rect 29092 19848 29144 19854
rect 29092 19790 29144 19796
rect 29184 19712 29236 19718
rect 29184 19654 29236 19660
rect 29196 19378 29224 19654
rect 29460 19508 29512 19514
rect 29460 19450 29512 19456
rect 29184 19372 29236 19378
rect 29184 19314 29236 19320
rect 29472 18970 29500 19450
rect 29460 18964 29512 18970
rect 29460 18906 29512 18912
rect 29564 18850 29592 22646
rect 29932 22642 29960 23054
rect 29920 22636 29972 22642
rect 29920 22578 29972 22584
rect 29828 21956 29880 21962
rect 29828 21898 29880 21904
rect 29472 18822 29592 18850
rect 29000 18624 29052 18630
rect 29000 18566 29052 18572
rect 29184 18148 29236 18154
rect 29184 18090 29236 18096
rect 29196 17678 29224 18090
rect 29184 17672 29236 17678
rect 29184 17614 29236 17620
rect 29276 17672 29328 17678
rect 29276 17614 29328 17620
rect 29092 17536 29144 17542
rect 29092 17478 29144 17484
rect 29104 17202 29132 17478
rect 29288 17338 29316 17614
rect 29276 17332 29328 17338
rect 29276 17274 29328 17280
rect 29092 17196 29144 17202
rect 29092 17138 29144 17144
rect 28908 17128 28960 17134
rect 28908 17070 28960 17076
rect 28920 16674 28948 17070
rect 28828 16646 28948 16674
rect 29000 16652 29052 16658
rect 28630 16552 28686 16561
rect 28630 16487 28686 16496
rect 28644 16182 28672 16487
rect 28632 16176 28684 16182
rect 28632 16118 28684 16124
rect 28540 16040 28592 16046
rect 28540 15982 28592 15988
rect 28552 15586 28580 15982
rect 28644 15706 28672 16118
rect 28828 16114 28856 16646
rect 29000 16594 29052 16600
rect 28908 16516 28960 16522
rect 28908 16458 28960 16464
rect 28920 16250 28948 16458
rect 28908 16244 28960 16250
rect 28908 16186 28960 16192
rect 28816 16108 28868 16114
rect 28816 16050 28868 16056
rect 28632 15700 28684 15706
rect 28632 15642 28684 15648
rect 28552 15558 28672 15586
rect 28644 15366 28672 15558
rect 28632 15360 28684 15366
rect 28632 15302 28684 15308
rect 28356 14408 28408 14414
rect 28356 14350 28408 14356
rect 28644 14346 28672 15302
rect 28920 15162 28948 16186
rect 29012 15502 29040 16594
rect 29000 15496 29052 15502
rect 29000 15438 29052 15444
rect 28908 15156 28960 15162
rect 28908 15098 28960 15104
rect 28920 14618 28948 15098
rect 29012 15026 29040 15438
rect 29000 15020 29052 15026
rect 29000 14962 29052 14968
rect 28908 14612 28960 14618
rect 28908 14554 28960 14560
rect 28632 14340 28684 14346
rect 28632 14282 28684 14288
rect 28264 13932 28316 13938
rect 28264 13874 28316 13880
rect 28644 13870 28672 14282
rect 28632 13864 28684 13870
rect 28632 13806 28684 13812
rect 28080 13728 28132 13734
rect 28080 13670 28132 13676
rect 28722 13424 28778 13433
rect 28722 13359 28778 13368
rect 28736 13326 28764 13359
rect 28724 13320 28776 13326
rect 28724 13262 28776 13268
rect 28264 13184 28316 13190
rect 28264 13126 28316 13132
rect 27988 12844 28040 12850
rect 27988 12786 28040 12792
rect 28000 12434 28028 12786
rect 28276 12442 28304 13126
rect 28920 12986 28948 14554
rect 29104 14346 29132 17138
rect 29288 15094 29316 17274
rect 29368 16992 29420 16998
rect 29368 16934 29420 16940
rect 29276 15088 29328 15094
rect 29276 15030 29328 15036
rect 29380 14822 29408 16934
rect 29472 15434 29500 18822
rect 29552 18760 29604 18766
rect 29552 18702 29604 18708
rect 29564 17202 29592 18702
rect 29736 18216 29788 18222
rect 29736 18158 29788 18164
rect 29748 17746 29776 18158
rect 29736 17740 29788 17746
rect 29736 17682 29788 17688
rect 29642 17504 29698 17513
rect 29642 17439 29698 17448
rect 29656 17270 29684 17439
rect 29644 17264 29696 17270
rect 29644 17206 29696 17212
rect 29552 17196 29604 17202
rect 29552 17138 29604 17144
rect 29564 16726 29592 17138
rect 29736 17060 29788 17066
rect 29736 17002 29788 17008
rect 29552 16720 29604 16726
rect 29552 16662 29604 16668
rect 29748 15570 29776 17002
rect 29736 15564 29788 15570
rect 29736 15506 29788 15512
rect 29460 15428 29512 15434
rect 29460 15370 29512 15376
rect 29552 15428 29604 15434
rect 29552 15370 29604 15376
rect 29564 15162 29592 15370
rect 29552 15156 29604 15162
rect 29552 15098 29604 15104
rect 29644 15020 29696 15026
rect 29644 14962 29696 14968
rect 29368 14816 29420 14822
rect 29368 14758 29420 14764
rect 29092 14340 29144 14346
rect 29092 14282 29144 14288
rect 29656 14278 29684 14962
rect 29736 14544 29788 14550
rect 29736 14486 29788 14492
rect 29748 14346 29776 14486
rect 29736 14340 29788 14346
rect 29736 14282 29788 14288
rect 29644 14272 29696 14278
rect 29644 14214 29696 14220
rect 29656 13870 29684 14214
rect 29184 13864 29236 13870
rect 29184 13806 29236 13812
rect 29644 13864 29696 13870
rect 29644 13806 29696 13812
rect 29000 13728 29052 13734
rect 29000 13670 29052 13676
rect 29012 13326 29040 13670
rect 29000 13320 29052 13326
rect 29000 13262 29052 13268
rect 29092 13320 29144 13326
rect 29092 13262 29144 13268
rect 28908 12980 28960 12986
rect 28908 12922 28960 12928
rect 29104 12850 29132 13262
rect 29196 13258 29224 13806
rect 29184 13252 29236 13258
rect 29184 13194 29236 13200
rect 29552 13184 29604 13190
rect 29552 13126 29604 13132
rect 29460 12912 29512 12918
rect 29460 12854 29512 12860
rect 29092 12844 29144 12850
rect 29092 12786 29144 12792
rect 27908 12406 28028 12434
rect 28264 12436 28316 12442
rect 27908 12306 27936 12406
rect 28264 12378 28316 12384
rect 27986 12336 28042 12345
rect 27896 12300 27948 12306
rect 27986 12271 28042 12280
rect 28080 12300 28132 12306
rect 27896 12242 27948 12248
rect 28000 12238 28028 12271
rect 28080 12242 28132 12248
rect 28172 12300 28224 12306
rect 28172 12242 28224 12248
rect 27988 12232 28040 12238
rect 27988 12174 28040 12180
rect 27896 11756 27948 11762
rect 27896 11698 27948 11704
rect 27804 11552 27856 11558
rect 27804 11494 27856 11500
rect 27816 9994 27844 11494
rect 27804 9988 27856 9994
rect 27804 9930 27856 9936
rect 27816 8566 27844 9930
rect 27804 8560 27856 8566
rect 27804 8502 27856 8508
rect 27712 8424 27764 8430
rect 27712 8366 27764 8372
rect 27724 7410 27752 8366
rect 27816 7954 27844 8502
rect 27804 7948 27856 7954
rect 27804 7890 27856 7896
rect 27712 7404 27764 7410
rect 27712 7346 27764 7352
rect 27804 7404 27856 7410
rect 27804 7346 27856 7352
rect 27620 6316 27672 6322
rect 27620 6258 27672 6264
rect 27632 5574 27660 6258
rect 27620 5568 27672 5574
rect 27620 5510 27672 5516
rect 27816 5234 27844 7346
rect 27304 5188 27384 5216
rect 27252 5170 27304 5176
rect 27356 4826 27384 5188
rect 27804 5228 27856 5234
rect 27804 5170 27856 5176
rect 27620 5024 27672 5030
rect 27620 4966 27672 4972
rect 27160 4820 27212 4826
rect 27160 4762 27212 4768
rect 27344 4820 27396 4826
rect 27344 4762 27396 4768
rect 26792 4208 26844 4214
rect 27632 4162 27660 4966
rect 27712 4548 27764 4554
rect 27712 4490 27764 4496
rect 26792 4150 26844 4156
rect 26804 3534 26832 4150
rect 27540 4146 27660 4162
rect 27344 4140 27396 4146
rect 27344 4082 27396 4088
rect 27528 4140 27660 4146
rect 27580 4134 27660 4140
rect 27528 4082 27580 4088
rect 27356 3602 27384 4082
rect 27724 3738 27752 4490
rect 27816 4010 27844 5170
rect 27908 4146 27936 11698
rect 28092 10266 28120 12242
rect 28184 11898 28212 12242
rect 29104 12238 29132 12786
rect 28264 12232 28316 12238
rect 29092 12232 29144 12238
rect 28264 12174 28316 12180
rect 28446 12200 28502 12209
rect 28172 11892 28224 11898
rect 28172 11834 28224 11840
rect 28184 11626 28212 11834
rect 28276 11626 28304 12174
rect 29092 12174 29144 12180
rect 28446 12135 28502 12144
rect 28460 12102 28488 12135
rect 28448 12096 28500 12102
rect 28448 12038 28500 12044
rect 29104 11762 29132 12174
rect 29184 12096 29236 12102
rect 29184 12038 29236 12044
rect 29092 11756 29144 11762
rect 29092 11698 29144 11704
rect 28172 11620 28224 11626
rect 28172 11562 28224 11568
rect 28264 11620 28316 11626
rect 28264 11562 28316 11568
rect 28184 11200 28212 11562
rect 28540 11552 28592 11558
rect 28540 11494 28592 11500
rect 29092 11552 29144 11558
rect 29092 11494 29144 11500
rect 28184 11172 28304 11200
rect 28080 10260 28132 10266
rect 28080 10202 28132 10208
rect 27988 9580 28040 9586
rect 27988 9522 28040 9528
rect 28000 9353 28028 9522
rect 28080 9512 28132 9518
rect 28080 9454 28132 9460
rect 27986 9344 28042 9353
rect 27986 9279 28042 9288
rect 28092 7546 28120 9454
rect 28172 9444 28224 9450
rect 28172 9386 28224 9392
rect 28184 8362 28212 9386
rect 28172 8356 28224 8362
rect 28172 8298 28224 8304
rect 28080 7540 28132 7546
rect 28080 7482 28132 7488
rect 28276 6118 28304 11172
rect 28552 11150 28580 11494
rect 28540 11144 28592 11150
rect 28540 11086 28592 11092
rect 28448 11076 28500 11082
rect 28448 11018 28500 11024
rect 28460 10062 28488 11018
rect 28814 10704 28870 10713
rect 28814 10639 28816 10648
rect 28868 10639 28870 10648
rect 28816 10610 28868 10616
rect 28998 10568 29054 10577
rect 28724 10532 28776 10538
rect 28998 10503 29054 10512
rect 28724 10474 28776 10480
rect 28540 10192 28592 10198
rect 28538 10160 28540 10169
rect 28592 10160 28594 10169
rect 28538 10095 28594 10104
rect 28736 10062 28764 10474
rect 29012 10062 29040 10503
rect 28448 10056 28500 10062
rect 28448 9998 28500 10004
rect 28724 10056 28776 10062
rect 28724 9998 28776 10004
rect 28816 10056 28868 10062
rect 29000 10056 29052 10062
rect 28816 9998 28868 10004
rect 28906 10024 28962 10033
rect 28460 9738 28488 9998
rect 28460 9710 28580 9738
rect 28446 9616 28502 9625
rect 28446 9551 28502 9560
rect 28460 9450 28488 9551
rect 28448 9444 28500 9450
rect 28448 9386 28500 9392
rect 28552 8514 28580 9710
rect 28828 8634 28856 9998
rect 29000 9998 29052 10004
rect 28906 9959 28962 9968
rect 28920 9586 28948 9959
rect 28908 9580 28960 9586
rect 28908 9522 28960 9528
rect 29000 9580 29052 9586
rect 29000 9522 29052 9528
rect 28920 9178 28948 9522
rect 28908 9172 28960 9178
rect 28908 9114 28960 9120
rect 28632 8628 28684 8634
rect 28816 8628 28868 8634
rect 28684 8588 28764 8616
rect 28632 8570 28684 8576
rect 28552 8498 28672 8514
rect 28552 8492 28684 8498
rect 28552 8486 28632 8492
rect 28632 8434 28684 8440
rect 28736 8430 28764 8588
rect 28816 8570 28868 8576
rect 28724 8424 28776 8430
rect 28724 8366 28776 8372
rect 28540 7948 28592 7954
rect 28540 7890 28592 7896
rect 28448 7472 28500 7478
rect 28448 7414 28500 7420
rect 28264 6112 28316 6118
rect 28264 6054 28316 6060
rect 28460 5710 28488 7414
rect 28552 7410 28580 7890
rect 29012 7546 29040 9522
rect 29104 9382 29132 11494
rect 29196 10266 29224 12038
rect 29472 11830 29500 12854
rect 29460 11824 29512 11830
rect 29460 11766 29512 11772
rect 29368 11756 29420 11762
rect 29368 11698 29420 11704
rect 29276 11348 29328 11354
rect 29276 11290 29328 11296
rect 29184 10260 29236 10266
rect 29184 10202 29236 10208
rect 29288 9450 29316 11290
rect 29380 11150 29408 11698
rect 29460 11280 29512 11286
rect 29460 11222 29512 11228
rect 29368 11144 29420 11150
rect 29368 11086 29420 11092
rect 29472 10606 29500 11222
rect 29460 10600 29512 10606
rect 29460 10542 29512 10548
rect 29564 10470 29592 13126
rect 29552 10464 29604 10470
rect 29552 10406 29604 10412
rect 29552 9512 29604 9518
rect 29552 9454 29604 9460
rect 29276 9444 29328 9450
rect 29276 9386 29328 9392
rect 29092 9376 29144 9382
rect 29092 9318 29144 9324
rect 29368 9376 29420 9382
rect 29368 9318 29420 9324
rect 29380 9081 29408 9318
rect 29366 9072 29422 9081
rect 29366 9007 29422 9016
rect 29276 8492 29328 8498
rect 29276 8434 29328 8440
rect 29460 8492 29512 8498
rect 29460 8434 29512 8440
rect 29092 7880 29144 7886
rect 29092 7822 29144 7828
rect 29000 7540 29052 7546
rect 29000 7482 29052 7488
rect 28540 7404 28592 7410
rect 28540 7346 28592 7352
rect 29104 7206 29132 7822
rect 29092 7200 29144 7206
rect 29092 7142 29144 7148
rect 28908 6656 28960 6662
rect 28908 6598 28960 6604
rect 28920 5914 28948 6598
rect 29104 6322 29132 7142
rect 29288 6798 29316 8434
rect 29472 7546 29500 8434
rect 29460 7540 29512 7546
rect 29460 7482 29512 7488
rect 29564 7410 29592 9454
rect 29656 7562 29684 13806
rect 29840 13734 29868 21898
rect 29920 20460 29972 20466
rect 29920 20402 29972 20408
rect 29932 16250 29960 20402
rect 30024 17202 30052 23462
rect 30472 23180 30524 23186
rect 30472 23122 30524 23128
rect 30484 22642 30512 23122
rect 30668 22642 30696 23462
rect 30932 23112 30984 23118
rect 30932 23054 30984 23060
rect 30196 22636 30248 22642
rect 30196 22578 30248 22584
rect 30380 22636 30432 22642
rect 30380 22578 30432 22584
rect 30472 22636 30524 22642
rect 30472 22578 30524 22584
rect 30656 22636 30708 22642
rect 30656 22578 30708 22584
rect 30208 21554 30236 22578
rect 30392 22234 30420 22578
rect 30380 22228 30432 22234
rect 30380 22170 30432 22176
rect 30944 22098 30972 23054
rect 31036 22982 31064 23666
rect 31116 23044 31168 23050
rect 31116 22986 31168 22992
rect 31024 22976 31076 22982
rect 31024 22918 31076 22924
rect 30932 22092 30984 22098
rect 30932 22034 30984 22040
rect 30562 21992 30618 22001
rect 30562 21927 30618 21936
rect 30196 21548 30248 21554
rect 30196 21490 30248 21496
rect 30104 20868 30156 20874
rect 30104 20810 30156 20816
rect 30012 17196 30064 17202
rect 30012 17138 30064 17144
rect 29920 16244 29972 16250
rect 29920 16186 29972 16192
rect 30012 15020 30064 15026
rect 30012 14962 30064 14968
rect 30024 14550 30052 14962
rect 30012 14544 30064 14550
rect 30012 14486 30064 14492
rect 29828 13728 29880 13734
rect 29828 13670 29880 13676
rect 29920 13252 29972 13258
rect 29920 13194 29972 13200
rect 29932 12238 29960 13194
rect 30116 12238 30144 20810
rect 30208 20058 30236 21490
rect 30288 20936 30340 20942
rect 30288 20878 30340 20884
rect 30196 20052 30248 20058
rect 30196 19994 30248 20000
rect 30208 19786 30236 19994
rect 30300 19990 30328 20878
rect 30472 20256 30524 20262
rect 30472 20198 30524 20204
rect 30288 19984 30340 19990
rect 30288 19926 30340 19932
rect 30300 19854 30328 19926
rect 30288 19848 30340 19854
rect 30288 19790 30340 19796
rect 30484 19786 30512 20198
rect 30196 19780 30248 19786
rect 30196 19722 30248 19728
rect 30472 19780 30524 19786
rect 30472 19722 30524 19728
rect 30380 19712 30432 19718
rect 30380 19654 30432 19660
rect 30196 19508 30248 19514
rect 30196 19450 30248 19456
rect 30208 18766 30236 19450
rect 30196 18760 30248 18766
rect 30196 18702 30248 18708
rect 29920 12232 29972 12238
rect 29920 12174 29972 12180
rect 30104 12232 30156 12238
rect 30104 12174 30156 12180
rect 29932 11830 29960 12174
rect 29920 11824 29972 11830
rect 29920 11766 29972 11772
rect 29932 11150 29960 11766
rect 30208 11150 30236 18702
rect 30288 18352 30340 18358
rect 30288 18294 30340 18300
rect 30300 18154 30328 18294
rect 30288 18148 30340 18154
rect 30288 18090 30340 18096
rect 30392 16425 30420 19654
rect 30378 16416 30434 16425
rect 30378 16351 30434 16360
rect 30484 11762 30512 19722
rect 30576 14550 30604 21927
rect 30656 21548 30708 21554
rect 30656 21490 30708 21496
rect 30840 21548 30892 21554
rect 30840 21490 30892 21496
rect 30668 21146 30696 21490
rect 30656 21140 30708 21146
rect 30656 21082 30708 21088
rect 30852 20806 30880 21490
rect 30840 20800 30892 20806
rect 30840 20742 30892 20748
rect 30852 19281 30880 20742
rect 30944 20534 30972 22034
rect 31036 22030 31064 22918
rect 31128 22778 31156 22986
rect 31116 22772 31168 22778
rect 31116 22714 31168 22720
rect 31116 22500 31168 22506
rect 31116 22442 31168 22448
rect 31024 22024 31076 22030
rect 31024 21966 31076 21972
rect 30932 20528 30984 20534
rect 30932 20470 30984 20476
rect 30944 19446 30972 20470
rect 31128 20330 31156 22442
rect 31208 21956 31260 21962
rect 31208 21898 31260 21904
rect 31220 21690 31248 21898
rect 31208 21684 31260 21690
rect 31208 21626 31260 21632
rect 31116 20324 31168 20330
rect 31116 20266 31168 20272
rect 31128 19446 31156 20266
rect 30932 19440 30984 19446
rect 30932 19382 30984 19388
rect 31116 19440 31168 19446
rect 31116 19382 31168 19388
rect 30838 19272 30894 19281
rect 30838 19207 30894 19216
rect 31024 18624 31076 18630
rect 31024 18566 31076 18572
rect 31036 18290 31064 18566
rect 31024 18284 31076 18290
rect 31024 18226 31076 18232
rect 31036 18193 31064 18226
rect 31116 18216 31168 18222
rect 31022 18184 31078 18193
rect 31116 18158 31168 18164
rect 31022 18119 31078 18128
rect 31024 18080 31076 18086
rect 31024 18022 31076 18028
rect 30840 17672 30892 17678
rect 30840 17614 30892 17620
rect 30852 16658 30880 17614
rect 31036 17202 31064 18022
rect 31128 17202 31156 18158
rect 31024 17196 31076 17202
rect 31024 17138 31076 17144
rect 31116 17196 31168 17202
rect 31116 17138 31168 17144
rect 30932 17128 30984 17134
rect 30932 17070 30984 17076
rect 30840 16652 30892 16658
rect 30840 16594 30892 16600
rect 30852 16114 30880 16594
rect 30840 16108 30892 16114
rect 30840 16050 30892 16056
rect 30944 14958 30972 17070
rect 31024 16992 31076 16998
rect 31024 16934 31076 16940
rect 31036 16794 31064 16934
rect 31024 16788 31076 16794
rect 31024 16730 31076 16736
rect 31036 15450 31064 16730
rect 31114 16552 31170 16561
rect 31114 16487 31116 16496
rect 31168 16487 31170 16496
rect 31208 16516 31260 16522
rect 31116 16458 31168 16464
rect 31208 16458 31260 16464
rect 31220 16114 31248 16458
rect 31208 16108 31260 16114
rect 31208 16050 31260 16056
rect 31036 15422 31156 15450
rect 31024 15360 31076 15366
rect 31024 15302 31076 15308
rect 30932 14952 30984 14958
rect 30932 14894 30984 14900
rect 30944 14550 30972 14894
rect 30564 14544 30616 14550
rect 30564 14486 30616 14492
rect 30932 14544 30984 14550
rect 30932 14486 30984 14492
rect 30576 14414 30604 14486
rect 30564 14408 30616 14414
rect 30564 14350 30616 14356
rect 31036 14346 31064 15302
rect 31128 15094 31156 15422
rect 31116 15088 31168 15094
rect 31116 15030 31168 15036
rect 31024 14340 31076 14346
rect 31024 14282 31076 14288
rect 30564 14000 30616 14006
rect 30564 13942 30616 13948
rect 30576 13462 30604 13942
rect 30564 13456 30616 13462
rect 30564 13398 30616 13404
rect 31312 13326 31340 23666
rect 31404 23186 31432 24142
rect 31392 23180 31444 23186
rect 31392 23122 31444 23128
rect 31484 22636 31536 22642
rect 31484 22578 31536 22584
rect 31496 22001 31524 22578
rect 31482 21992 31538 22001
rect 31482 21927 31538 21936
rect 31392 21480 31444 21486
rect 31392 21422 31444 21428
rect 31404 19854 31432 21422
rect 31392 19848 31444 19854
rect 31392 19790 31444 19796
rect 31484 18692 31536 18698
rect 31484 18634 31536 18640
rect 31392 18148 31444 18154
rect 31392 18090 31444 18096
rect 31404 17678 31432 18090
rect 31392 17672 31444 17678
rect 31392 17614 31444 17620
rect 31404 17542 31432 17614
rect 31392 17536 31444 17542
rect 31392 17478 31444 17484
rect 31392 17264 31444 17270
rect 31392 17206 31444 17212
rect 31404 15910 31432 17206
rect 31496 17202 31524 18634
rect 31484 17196 31536 17202
rect 31484 17138 31536 17144
rect 31496 16454 31524 17138
rect 31588 16590 31616 25910
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 65654 25596 65962 25605
rect 65654 25594 65660 25596
rect 65716 25594 65740 25596
rect 65796 25594 65820 25596
rect 65876 25594 65900 25596
rect 65956 25594 65962 25596
rect 65716 25542 65718 25594
rect 65898 25542 65900 25594
rect 65654 25540 65660 25542
rect 65716 25540 65740 25542
rect 65796 25540 65820 25542
rect 65876 25540 65900 25542
rect 65956 25540 65962 25542
rect 65654 25531 65962 25540
rect 33968 25288 34020 25294
rect 68100 25288 68152 25294
rect 33968 25230 34020 25236
rect 68098 25256 68100 25265
rect 68152 25256 68154 25265
rect 31668 25152 31720 25158
rect 31668 25094 31720 25100
rect 31680 24818 31708 25094
rect 31668 24812 31720 24818
rect 31668 24754 31720 24760
rect 31576 16584 31628 16590
rect 31576 16526 31628 16532
rect 31484 16448 31536 16454
rect 31484 16390 31536 16396
rect 31680 16114 31708 24754
rect 33980 24206 34008 25230
rect 68098 25191 68154 25200
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 65654 24508 65962 24517
rect 65654 24506 65660 24508
rect 65716 24506 65740 24508
rect 65796 24506 65820 24508
rect 65876 24506 65900 24508
rect 65956 24506 65962 24508
rect 65716 24454 65718 24506
rect 65898 24454 65900 24506
rect 65654 24452 65660 24454
rect 65716 24452 65740 24454
rect 65796 24452 65820 24454
rect 65876 24452 65900 24454
rect 65956 24452 65962 24454
rect 65654 24443 65962 24452
rect 33968 24200 34020 24206
rect 33968 24142 34020 24148
rect 68100 24200 68152 24206
rect 68100 24142 68152 24148
rect 32588 24064 32640 24070
rect 32588 24006 32640 24012
rect 32600 23730 32628 24006
rect 32588 23724 32640 23730
rect 32588 23666 32640 23672
rect 32956 22976 33008 22982
rect 32956 22918 33008 22924
rect 32968 22030 32996 22918
rect 32956 22024 33008 22030
rect 32956 21966 33008 21972
rect 33600 21956 33652 21962
rect 33600 21898 33652 21904
rect 32128 21888 32180 21894
rect 32128 21830 32180 21836
rect 32312 21888 32364 21894
rect 32312 21830 32364 21836
rect 32772 21888 32824 21894
rect 32772 21830 32824 21836
rect 32140 21486 32168 21830
rect 32128 21480 32180 21486
rect 32128 21422 32180 21428
rect 32324 20874 32352 21830
rect 32784 21622 32812 21830
rect 32772 21616 32824 21622
rect 32772 21558 32824 21564
rect 33416 21548 33468 21554
rect 33416 21490 33468 21496
rect 33140 21344 33192 21350
rect 33140 21286 33192 21292
rect 33152 20942 33180 21286
rect 33140 20936 33192 20942
rect 33140 20878 33192 20884
rect 32312 20868 32364 20874
rect 32312 20810 32364 20816
rect 33428 20466 33456 21490
rect 33612 21146 33640 21898
rect 33980 21622 34008 24142
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 68112 23905 68140 24142
rect 68098 23896 68154 23905
rect 68098 23831 68154 23840
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 65654 23420 65962 23429
rect 65654 23418 65660 23420
rect 65716 23418 65740 23420
rect 65796 23418 65820 23420
rect 65876 23418 65900 23420
rect 65956 23418 65962 23420
rect 65716 23366 65718 23418
rect 65898 23366 65900 23418
rect 65654 23364 65660 23366
rect 65716 23364 65740 23366
rect 65796 23364 65820 23366
rect 65876 23364 65900 23366
rect 65956 23364 65962 23366
rect 65654 23355 65962 23364
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 67638 22536 67694 22545
rect 67638 22471 67640 22480
rect 67692 22471 67694 22480
rect 67640 22442 67692 22448
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 65654 22332 65962 22341
rect 65654 22330 65660 22332
rect 65716 22330 65740 22332
rect 65796 22330 65820 22332
rect 65876 22330 65900 22332
rect 65956 22330 65962 22332
rect 65716 22278 65718 22330
rect 65898 22278 65900 22330
rect 65654 22276 65660 22278
rect 65716 22276 65740 22278
rect 65796 22276 65820 22278
rect 65876 22276 65900 22278
rect 65956 22276 65962 22278
rect 65654 22267 65962 22276
rect 34152 22024 34204 22030
rect 34152 21966 34204 21972
rect 33968 21616 34020 21622
rect 33968 21558 34020 21564
rect 33600 21140 33652 21146
rect 33600 21082 33652 21088
rect 33508 20868 33560 20874
rect 33508 20810 33560 20816
rect 31760 20460 31812 20466
rect 31760 20402 31812 20408
rect 33416 20460 33468 20466
rect 33416 20402 33468 20408
rect 31772 20058 31800 20402
rect 31760 20052 31812 20058
rect 31760 19994 31812 20000
rect 33520 19446 33548 20810
rect 34164 20330 34192 21966
rect 35900 21888 35952 21894
rect 35900 21830 35952 21836
rect 37648 21888 37700 21894
rect 37648 21830 37700 21836
rect 35624 21548 35676 21554
rect 35624 21490 35676 21496
rect 34796 21344 34848 21350
rect 34796 21286 34848 21292
rect 34808 21010 34836 21286
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 35636 21146 35664 21490
rect 35624 21140 35676 21146
rect 35624 21082 35676 21088
rect 34520 21004 34572 21010
rect 34520 20946 34572 20952
rect 34796 21004 34848 21010
rect 34796 20946 34848 20952
rect 34152 20324 34204 20330
rect 34152 20266 34204 20272
rect 33508 19440 33560 19446
rect 33508 19382 33560 19388
rect 33140 19304 33192 19310
rect 33140 19246 33192 19252
rect 33152 18766 33180 19246
rect 33324 19168 33376 19174
rect 33324 19110 33376 19116
rect 32956 18760 33008 18766
rect 32956 18702 33008 18708
rect 33140 18760 33192 18766
rect 33140 18702 33192 18708
rect 31944 18692 31996 18698
rect 31944 18634 31996 18640
rect 31760 17740 31812 17746
rect 31760 17682 31812 17688
rect 31772 17270 31800 17682
rect 31956 17338 31984 18634
rect 32312 17672 32364 17678
rect 32312 17614 32364 17620
rect 31944 17332 31996 17338
rect 31944 17274 31996 17280
rect 31760 17264 31812 17270
rect 31760 17206 31812 17212
rect 32128 16516 32180 16522
rect 32128 16458 32180 16464
rect 31668 16108 31720 16114
rect 31668 16050 31720 16056
rect 31392 15904 31444 15910
rect 31392 15846 31444 15852
rect 31404 15026 31432 15846
rect 32140 15094 32168 16458
rect 32324 16114 32352 17614
rect 32968 17270 32996 18702
rect 33152 17746 33180 18702
rect 33336 18358 33364 19110
rect 33324 18352 33376 18358
rect 33322 18320 33324 18329
rect 33376 18320 33378 18329
rect 33322 18255 33378 18264
rect 33336 18229 33364 18255
rect 33520 18222 33548 19382
rect 33876 19372 33928 19378
rect 33876 19314 33928 19320
rect 33692 19236 33744 19242
rect 33692 19178 33744 19184
rect 33600 18760 33652 18766
rect 33600 18702 33652 18708
rect 33508 18216 33560 18222
rect 33508 18158 33560 18164
rect 33416 18080 33468 18086
rect 33416 18022 33468 18028
rect 33140 17740 33192 17746
rect 33140 17682 33192 17688
rect 33428 17678 33456 18022
rect 33520 17678 33548 18158
rect 33232 17672 33284 17678
rect 33232 17614 33284 17620
rect 33416 17672 33468 17678
rect 33416 17614 33468 17620
rect 33508 17672 33560 17678
rect 33508 17614 33560 17620
rect 32956 17264 33008 17270
rect 32956 17206 33008 17212
rect 32496 16992 32548 16998
rect 32496 16934 32548 16940
rect 32508 16114 32536 16934
rect 32968 16658 32996 17206
rect 33140 17196 33192 17202
rect 33140 17138 33192 17144
rect 32956 16652 33008 16658
rect 32956 16594 33008 16600
rect 32864 16584 32916 16590
rect 32864 16526 32916 16532
rect 32588 16448 32640 16454
rect 32588 16390 32640 16396
rect 32312 16108 32364 16114
rect 32312 16050 32364 16056
rect 32496 16108 32548 16114
rect 32496 16050 32548 16056
rect 32600 16096 32628 16390
rect 32876 16182 32904 16526
rect 32864 16176 32916 16182
rect 32864 16118 32916 16124
rect 32680 16108 32732 16114
rect 32600 16068 32680 16096
rect 32324 15502 32352 16050
rect 32496 15564 32548 15570
rect 32496 15506 32548 15512
rect 32312 15496 32364 15502
rect 32312 15438 32364 15444
rect 32508 15162 32536 15506
rect 32600 15366 32628 16068
rect 32680 16050 32732 16056
rect 32876 15638 32904 16118
rect 32968 16046 32996 16594
rect 33152 16250 33180 17138
rect 33244 16794 33272 17614
rect 33232 16788 33284 16794
rect 33232 16730 33284 16736
rect 33416 16584 33468 16590
rect 33416 16526 33468 16532
rect 33140 16244 33192 16250
rect 33140 16186 33192 16192
rect 32956 16040 33008 16046
rect 32956 15982 33008 15988
rect 32864 15632 32916 15638
rect 32864 15574 32916 15580
rect 32588 15360 32640 15366
rect 32588 15302 32640 15308
rect 32772 15360 32824 15366
rect 32772 15302 32824 15308
rect 32496 15156 32548 15162
rect 32496 15098 32548 15104
rect 32128 15088 32180 15094
rect 32128 15030 32180 15036
rect 32312 15088 32364 15094
rect 32312 15030 32364 15036
rect 31392 15020 31444 15026
rect 31392 14962 31444 14968
rect 31484 15020 31536 15026
rect 31484 14962 31536 14968
rect 31496 14278 31524 14962
rect 31576 14408 31628 14414
rect 31668 14408 31720 14414
rect 31628 14368 31668 14396
rect 31576 14350 31628 14356
rect 31668 14350 31720 14356
rect 31484 14272 31536 14278
rect 31484 14214 31536 14220
rect 32140 13938 32168 15030
rect 32324 14550 32352 15030
rect 32312 14544 32364 14550
rect 32312 14486 32364 14492
rect 32496 14068 32548 14074
rect 32496 14010 32548 14016
rect 32128 13932 32180 13938
rect 32128 13874 32180 13880
rect 31300 13320 31352 13326
rect 31300 13262 31352 13268
rect 31944 13320 31996 13326
rect 31944 13262 31996 13268
rect 31852 12844 31904 12850
rect 31852 12786 31904 12792
rect 30656 12640 30708 12646
rect 30656 12582 30708 12588
rect 30668 12434 30696 12582
rect 30668 12406 30788 12434
rect 30472 11756 30524 11762
rect 30472 11698 30524 11704
rect 30288 11552 30340 11558
rect 30288 11494 30340 11500
rect 30300 11218 30328 11494
rect 30656 11280 30708 11286
rect 30656 11222 30708 11228
rect 30288 11212 30340 11218
rect 30288 11154 30340 11160
rect 29920 11144 29972 11150
rect 29920 11086 29972 11092
rect 30196 11144 30248 11150
rect 30196 11086 30248 11092
rect 30668 10674 30696 11222
rect 30760 10742 30788 12406
rect 31864 11150 31892 12786
rect 31956 11762 31984 13262
rect 32140 12850 32168 13874
rect 32404 13728 32456 13734
rect 32404 13670 32456 13676
rect 32312 13388 32364 13394
rect 32312 13330 32364 13336
rect 32128 12844 32180 12850
rect 32128 12786 32180 12792
rect 32324 12238 32352 13330
rect 32416 13258 32444 13670
rect 32404 13252 32456 13258
rect 32404 13194 32456 13200
rect 32312 12232 32364 12238
rect 32312 12174 32364 12180
rect 32324 11898 32352 12174
rect 32128 11892 32180 11898
rect 32128 11834 32180 11840
rect 32312 11892 32364 11898
rect 32312 11834 32364 11840
rect 31944 11756 31996 11762
rect 31944 11698 31996 11704
rect 31852 11144 31904 11150
rect 31852 11086 31904 11092
rect 30748 10736 30800 10742
rect 30748 10678 30800 10684
rect 30656 10668 30708 10674
rect 30656 10610 30708 10616
rect 31392 10260 31444 10266
rect 31392 10202 31444 10208
rect 31404 9926 31432 10202
rect 31392 9920 31444 9926
rect 31392 9862 31444 9868
rect 29736 9580 29788 9586
rect 29736 9522 29788 9528
rect 29748 9110 29776 9522
rect 31116 9376 31168 9382
rect 31116 9318 31168 9324
rect 30838 9208 30894 9217
rect 30838 9143 30840 9152
rect 30892 9143 30894 9152
rect 30840 9114 30892 9120
rect 29736 9104 29788 9110
rect 29736 9046 29788 9052
rect 31128 8974 31156 9318
rect 31404 8974 31432 9862
rect 31024 8968 31076 8974
rect 31024 8910 31076 8916
rect 31116 8968 31168 8974
rect 31116 8910 31168 8916
rect 31392 8968 31444 8974
rect 31392 8910 31444 8916
rect 31036 8566 31064 8910
rect 31208 8900 31260 8906
rect 31208 8842 31260 8848
rect 31024 8560 31076 8566
rect 31024 8502 31076 8508
rect 31220 8362 31248 8842
rect 32140 8634 32168 11834
rect 32508 11762 32536 14010
rect 32496 11756 32548 11762
rect 32496 11698 32548 11704
rect 32508 11218 32536 11698
rect 32600 11234 32628 15302
rect 32784 14074 32812 15302
rect 32772 14068 32824 14074
rect 32772 14010 32824 14016
rect 32784 13394 32812 14010
rect 32876 13802 32904 15574
rect 32956 15360 33008 15366
rect 32956 15302 33008 15308
rect 33232 15360 33284 15366
rect 33232 15302 33284 15308
rect 33324 15360 33376 15366
rect 33324 15302 33376 15308
rect 32968 14278 32996 15302
rect 33244 15094 33272 15302
rect 33232 15088 33284 15094
rect 33232 15030 33284 15036
rect 33140 14408 33192 14414
rect 33140 14350 33192 14356
rect 32956 14272 33008 14278
rect 32954 14240 32956 14249
rect 33008 14240 33010 14249
rect 32954 14175 33010 14184
rect 32864 13796 32916 13802
rect 32864 13738 32916 13744
rect 32772 13388 32824 13394
rect 32772 13330 32824 13336
rect 32772 13184 32824 13190
rect 32772 13126 32824 13132
rect 32784 12918 32812 13126
rect 32772 12912 32824 12918
rect 32772 12854 32824 12860
rect 32876 12764 32904 13738
rect 32784 12736 32904 12764
rect 32680 12640 32732 12646
rect 32680 12582 32732 12588
rect 32692 12374 32720 12582
rect 32784 12374 32812 12736
rect 32680 12368 32732 12374
rect 32680 12310 32732 12316
rect 32772 12368 32824 12374
rect 32772 12310 32824 12316
rect 32784 11830 32812 12310
rect 32772 11824 32824 11830
rect 32772 11766 32824 11772
rect 32680 11756 32732 11762
rect 32680 11698 32732 11704
rect 32692 11354 32720 11698
rect 32680 11348 32732 11354
rect 32680 11290 32732 11296
rect 32220 11212 32272 11218
rect 32220 11154 32272 11160
rect 32496 11212 32548 11218
rect 32600 11206 32720 11234
rect 32496 11154 32548 11160
rect 32128 8628 32180 8634
rect 32128 8570 32180 8576
rect 31208 8356 31260 8362
rect 31208 8298 31260 8304
rect 32232 8294 32260 11154
rect 32588 11076 32640 11082
rect 32588 11018 32640 11024
rect 32600 10266 32628 11018
rect 32692 10810 32720 11206
rect 32680 10804 32732 10810
rect 32680 10746 32732 10752
rect 32692 10674 32720 10746
rect 32680 10668 32732 10674
rect 32680 10610 32732 10616
rect 32588 10260 32640 10266
rect 32588 10202 32640 10208
rect 32692 9722 32720 10610
rect 32680 9716 32732 9722
rect 32680 9658 32732 9664
rect 32496 8832 32548 8838
rect 32496 8774 32548 8780
rect 32508 8566 32536 8774
rect 32496 8560 32548 8566
rect 32496 8502 32548 8508
rect 32404 8492 32456 8498
rect 32404 8434 32456 8440
rect 32588 8492 32640 8498
rect 32588 8434 32640 8440
rect 29736 8288 29788 8294
rect 29736 8230 29788 8236
rect 32140 8266 32260 8294
rect 29748 8022 29776 8230
rect 29736 8016 29788 8022
rect 29736 7958 29788 7964
rect 29828 8016 29880 8022
rect 29828 7958 29880 7964
rect 29656 7534 29776 7562
rect 29644 7472 29696 7478
rect 29644 7414 29696 7420
rect 29552 7404 29604 7410
rect 29552 7346 29604 7352
rect 29656 6798 29684 7414
rect 29276 6792 29328 6798
rect 29276 6734 29328 6740
rect 29644 6792 29696 6798
rect 29644 6734 29696 6740
rect 29288 6474 29316 6734
rect 29552 6656 29604 6662
rect 29552 6598 29604 6604
rect 29196 6446 29316 6474
rect 29092 6316 29144 6322
rect 29092 6258 29144 6264
rect 29000 6248 29052 6254
rect 29000 6190 29052 6196
rect 28908 5908 28960 5914
rect 28908 5850 28960 5856
rect 28448 5704 28500 5710
rect 28448 5646 28500 5652
rect 28460 5370 28488 5646
rect 28448 5364 28500 5370
rect 28448 5306 28500 5312
rect 29012 5302 29040 6190
rect 29104 5710 29132 6258
rect 29092 5704 29144 5710
rect 29092 5646 29144 5652
rect 29196 5642 29224 6446
rect 29564 6322 29592 6598
rect 29656 6458 29684 6734
rect 29644 6452 29696 6458
rect 29644 6394 29696 6400
rect 29748 6390 29776 7534
rect 29840 6934 29868 7958
rect 31208 7880 31260 7886
rect 31208 7822 31260 7828
rect 30196 7744 30248 7750
rect 30196 7686 30248 7692
rect 30208 7478 30236 7686
rect 30196 7472 30248 7478
rect 30196 7414 30248 7420
rect 31220 7342 31248 7822
rect 31208 7336 31260 7342
rect 31208 7278 31260 7284
rect 31576 7336 31628 7342
rect 31576 7278 31628 7284
rect 29828 6928 29880 6934
rect 29828 6870 29880 6876
rect 30196 6928 30248 6934
rect 30196 6870 30248 6876
rect 29920 6656 29972 6662
rect 29920 6598 29972 6604
rect 29736 6384 29788 6390
rect 29736 6326 29788 6332
rect 29552 6316 29604 6322
rect 29552 6258 29604 6264
rect 29276 6180 29328 6186
rect 29276 6122 29328 6128
rect 29288 5914 29316 6122
rect 29276 5908 29328 5914
rect 29276 5850 29328 5856
rect 29932 5710 29960 6598
rect 30208 6254 30236 6870
rect 31588 6866 31616 7278
rect 31576 6860 31628 6866
rect 31576 6802 31628 6808
rect 30472 6316 30524 6322
rect 30472 6258 30524 6264
rect 30196 6248 30248 6254
rect 30196 6190 30248 6196
rect 29920 5704 29972 5710
rect 29920 5646 29972 5652
rect 30104 5704 30156 5710
rect 30208 5692 30236 6190
rect 30288 6112 30340 6118
rect 30288 6054 30340 6060
rect 30300 5710 30328 6054
rect 30484 5914 30512 6258
rect 31588 6254 31616 6802
rect 32140 6730 32168 8266
rect 32128 6724 32180 6730
rect 32128 6666 32180 6672
rect 31576 6248 31628 6254
rect 31576 6190 31628 6196
rect 30564 6180 30616 6186
rect 30564 6122 30616 6128
rect 30472 5908 30524 5914
rect 30472 5850 30524 5856
rect 30156 5664 30236 5692
rect 30288 5704 30340 5710
rect 30104 5646 30156 5652
rect 30288 5646 30340 5652
rect 29184 5636 29236 5642
rect 29184 5578 29236 5584
rect 29000 5296 29052 5302
rect 29000 5238 29052 5244
rect 29012 4690 29040 5238
rect 30576 5234 30604 6122
rect 30932 6112 30984 6118
rect 30932 6054 30984 6060
rect 30944 5846 30972 6054
rect 30932 5840 30984 5846
rect 30932 5782 30984 5788
rect 31588 5642 31616 6190
rect 31576 5636 31628 5642
rect 31576 5578 31628 5584
rect 31588 5302 31616 5578
rect 30840 5296 30892 5302
rect 30840 5238 30892 5244
rect 31576 5296 31628 5302
rect 31576 5238 31628 5244
rect 30564 5228 30616 5234
rect 30564 5170 30616 5176
rect 29000 4684 29052 4690
rect 29000 4626 29052 4632
rect 30852 4146 30880 5238
rect 32416 4622 32444 8434
rect 32600 7750 32628 8434
rect 32692 8362 32720 9658
rect 32680 8356 32732 8362
rect 32680 8298 32732 8304
rect 32968 7886 32996 14175
rect 33152 14006 33180 14350
rect 33140 14000 33192 14006
rect 33140 13942 33192 13948
rect 33048 13728 33100 13734
rect 33048 13670 33100 13676
rect 33060 13433 33088 13670
rect 33046 13424 33102 13433
rect 33046 13359 33102 13368
rect 33140 13252 33192 13258
rect 33140 13194 33192 13200
rect 33152 12442 33180 13194
rect 33140 12436 33192 12442
rect 33140 12378 33192 12384
rect 33232 10464 33284 10470
rect 33232 10406 33284 10412
rect 33244 10062 33272 10406
rect 33232 10056 33284 10062
rect 33232 9998 33284 10004
rect 33336 9042 33364 15302
rect 33428 12102 33456 16526
rect 33612 16114 33640 18702
rect 33704 17954 33732 19178
rect 33704 17926 33824 17954
rect 33796 17814 33824 17926
rect 33888 17882 33916 19314
rect 34532 18970 34560 20946
rect 34980 20936 35032 20942
rect 34980 20878 35032 20884
rect 34992 20806 35020 20878
rect 35440 20868 35492 20874
rect 35440 20810 35492 20816
rect 35716 20868 35768 20874
rect 35716 20810 35768 20816
rect 34796 20800 34848 20806
rect 34796 20742 34848 20748
rect 34980 20800 35032 20806
rect 34980 20742 35032 20748
rect 34808 20466 34836 20742
rect 34704 20460 34756 20466
rect 34704 20402 34756 20408
rect 34796 20460 34848 20466
rect 34796 20402 34848 20408
rect 34716 19786 34744 20402
rect 34704 19780 34756 19786
rect 34704 19722 34756 19728
rect 34520 18964 34572 18970
rect 34520 18906 34572 18912
rect 34612 18896 34664 18902
rect 34612 18838 34664 18844
rect 33876 17876 33928 17882
rect 33876 17818 33928 17824
rect 33784 17808 33836 17814
rect 33784 17750 33836 17756
rect 33690 16280 33746 16289
rect 33690 16215 33746 16224
rect 33600 16108 33652 16114
rect 33600 16050 33652 16056
rect 33704 16046 33732 16215
rect 33692 16040 33744 16046
rect 33692 15982 33744 15988
rect 33704 15638 33732 15982
rect 33692 15632 33744 15638
rect 33692 15574 33744 15580
rect 33416 12096 33468 12102
rect 33416 12038 33468 12044
rect 33692 11008 33744 11014
rect 33692 10950 33744 10956
rect 33704 10674 33732 10950
rect 33692 10668 33744 10674
rect 33692 10610 33744 10616
rect 33796 10656 33824 17750
rect 34624 17746 34652 18838
rect 34716 18290 34744 19722
rect 34808 19718 34836 20402
rect 35452 20330 35480 20810
rect 35728 20602 35756 20810
rect 35716 20596 35768 20602
rect 35716 20538 35768 20544
rect 35532 20460 35584 20466
rect 35532 20402 35584 20408
rect 35348 20324 35400 20330
rect 35348 20266 35400 20272
rect 35440 20324 35492 20330
rect 35440 20266 35492 20272
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35360 19854 35388 20266
rect 35348 19848 35400 19854
rect 35348 19790 35400 19796
rect 34796 19712 34848 19718
rect 34796 19654 34848 19660
rect 35256 19712 35308 19718
rect 35256 19654 35308 19660
rect 34808 19378 34836 19654
rect 35268 19378 35296 19654
rect 34796 19372 34848 19378
rect 34796 19314 34848 19320
rect 35164 19372 35216 19378
rect 35164 19314 35216 19320
rect 35256 19372 35308 19378
rect 35256 19314 35308 19320
rect 35176 19174 35204 19314
rect 35360 19242 35388 19790
rect 35348 19236 35400 19242
rect 35348 19178 35400 19184
rect 35164 19168 35216 19174
rect 35164 19110 35216 19116
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35360 18834 35388 19178
rect 35348 18828 35400 18834
rect 35348 18770 35400 18776
rect 35360 18290 35388 18770
rect 34704 18284 34756 18290
rect 34704 18226 34756 18232
rect 35348 18284 35400 18290
rect 35348 18226 35400 18232
rect 35440 18284 35492 18290
rect 35440 18226 35492 18232
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34612 17740 34664 17746
rect 34612 17682 34664 17688
rect 34796 17672 34848 17678
rect 34796 17614 34848 17620
rect 33968 17536 34020 17542
rect 33968 17478 34020 17484
rect 34704 17536 34756 17542
rect 34704 17478 34756 17484
rect 33980 11354 34008 17478
rect 34520 16516 34572 16522
rect 34520 16458 34572 16464
rect 34060 16448 34112 16454
rect 34060 16390 34112 16396
rect 34072 16114 34100 16390
rect 34532 16250 34560 16458
rect 34520 16244 34572 16250
rect 34520 16186 34572 16192
rect 34060 16108 34112 16114
rect 34060 16050 34112 16056
rect 34428 14952 34480 14958
rect 34428 14894 34480 14900
rect 34244 14408 34296 14414
rect 34244 14350 34296 14356
rect 34256 14006 34284 14350
rect 34440 14278 34468 14894
rect 34428 14272 34480 14278
rect 34428 14214 34480 14220
rect 34244 14000 34296 14006
rect 34244 13942 34296 13948
rect 34440 13394 34468 14214
rect 34520 14068 34572 14074
rect 34520 14010 34572 14016
rect 34428 13388 34480 13394
rect 34428 13330 34480 13336
rect 34532 12442 34560 14010
rect 34716 13977 34744 17478
rect 34808 16794 34836 17614
rect 35360 17202 35388 18226
rect 35452 17882 35480 18226
rect 35440 17876 35492 17882
rect 35440 17818 35492 17824
rect 35544 17610 35572 20402
rect 35808 19780 35860 19786
rect 35808 19722 35860 19728
rect 35820 19514 35848 19722
rect 35808 19508 35860 19514
rect 35808 19450 35860 19456
rect 35716 19372 35768 19378
rect 35716 19314 35768 19320
rect 35624 19168 35676 19174
rect 35624 19110 35676 19116
rect 35636 18714 35664 19110
rect 35728 18902 35756 19314
rect 35716 18896 35768 18902
rect 35716 18838 35768 18844
rect 35636 18686 35756 18714
rect 35532 17604 35584 17610
rect 35532 17546 35584 17552
rect 35624 17536 35676 17542
rect 35624 17478 35676 17484
rect 35636 17202 35664 17478
rect 35348 17196 35400 17202
rect 35348 17138 35400 17144
rect 35624 17196 35676 17202
rect 35624 17138 35676 17144
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34796 16788 34848 16794
rect 34796 16730 34848 16736
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 35348 15428 35400 15434
rect 35348 15370 35400 15376
rect 35256 15020 35308 15026
rect 35360 15008 35388 15370
rect 35728 15366 35756 18686
rect 35912 18630 35940 21830
rect 37660 21622 37688 21830
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 37648 21616 37700 21622
rect 37648 21558 37700 21564
rect 37660 21146 37688 21558
rect 67640 21344 67692 21350
rect 67640 21286 67692 21292
rect 65654 21244 65962 21253
rect 65654 21242 65660 21244
rect 65716 21242 65740 21244
rect 65796 21242 65820 21244
rect 65876 21242 65900 21244
rect 65956 21242 65962 21244
rect 65716 21190 65718 21242
rect 65898 21190 65900 21242
rect 65654 21188 65660 21190
rect 65716 21188 65740 21190
rect 65796 21188 65820 21190
rect 65876 21188 65900 21190
rect 65956 21188 65962 21190
rect 65654 21179 65962 21188
rect 67652 21185 67680 21286
rect 67638 21176 67694 21185
rect 37648 21140 37700 21146
rect 67638 21111 67694 21120
rect 37648 21082 37700 21088
rect 38200 21004 38252 21010
rect 38200 20946 38252 20952
rect 37464 20936 37516 20942
rect 37464 20878 37516 20884
rect 36636 20800 36688 20806
rect 36636 20742 36688 20748
rect 36648 20534 36676 20742
rect 36636 20528 36688 20534
rect 36636 20470 36688 20476
rect 37476 20330 37504 20878
rect 38212 20466 38240 20946
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 38200 20460 38252 20466
rect 38200 20402 38252 20408
rect 38292 20460 38344 20466
rect 38292 20402 38344 20408
rect 37464 20324 37516 20330
rect 37464 20266 37516 20272
rect 38200 20324 38252 20330
rect 38200 20266 38252 20272
rect 37648 20256 37700 20262
rect 37648 20198 37700 20204
rect 37660 19786 37688 20198
rect 37464 19780 37516 19786
rect 37464 19722 37516 19728
rect 37648 19780 37700 19786
rect 37648 19722 37700 19728
rect 37372 19304 37424 19310
rect 37372 19246 37424 19252
rect 37096 18964 37148 18970
rect 37096 18906 37148 18912
rect 35900 18624 35952 18630
rect 35900 18566 35952 18572
rect 35808 17672 35860 17678
rect 35808 17614 35860 17620
rect 35820 17542 35848 17614
rect 35808 17536 35860 17542
rect 35808 17478 35860 17484
rect 35808 15564 35860 15570
rect 35808 15506 35860 15512
rect 35716 15360 35768 15366
rect 35716 15302 35768 15308
rect 35820 15026 35848 15506
rect 35308 14980 35388 15008
rect 35256 14962 35308 14968
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34702 13968 34758 13977
rect 34702 13903 34758 13912
rect 34716 13462 34744 13903
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 35360 13546 35388 14980
rect 35440 15020 35492 15026
rect 35440 14962 35492 14968
rect 35808 15020 35860 15026
rect 35808 14962 35860 14968
rect 35268 13518 35388 13546
rect 34704 13456 34756 13462
rect 34704 13398 34756 13404
rect 35268 12782 35296 13518
rect 35348 13320 35400 13326
rect 35348 13262 35400 13268
rect 35256 12776 35308 12782
rect 35256 12718 35308 12724
rect 34796 12640 34848 12646
rect 34796 12582 34848 12588
rect 34520 12436 34572 12442
rect 34520 12378 34572 12384
rect 34532 11506 34560 12378
rect 34808 12306 34836 12582
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 35360 12442 35388 13262
rect 35452 12918 35480 14962
rect 35532 13864 35584 13870
rect 35532 13806 35584 13812
rect 35544 13326 35572 13806
rect 35532 13320 35584 13326
rect 35532 13262 35584 13268
rect 35440 12912 35492 12918
rect 35440 12854 35492 12860
rect 35716 12912 35768 12918
rect 35716 12854 35768 12860
rect 35440 12776 35492 12782
rect 35440 12718 35492 12724
rect 35348 12436 35400 12442
rect 35348 12378 35400 12384
rect 34796 12300 34848 12306
rect 34796 12242 34848 12248
rect 35072 12096 35124 12102
rect 35072 12038 35124 12044
rect 35084 11830 35112 12038
rect 35072 11824 35124 11830
rect 35072 11766 35124 11772
rect 34440 11478 34560 11506
rect 33968 11348 34020 11354
rect 33968 11290 34020 11296
rect 33876 10668 33928 10674
rect 33796 10628 33876 10656
rect 33600 9580 33652 9586
rect 33600 9522 33652 9528
rect 33612 9178 33640 9522
rect 33600 9172 33652 9178
rect 33600 9114 33652 9120
rect 33324 9036 33376 9042
rect 33324 8978 33376 8984
rect 33796 8022 33824 10628
rect 33876 10610 33928 10616
rect 34244 9988 34296 9994
rect 34244 9930 34296 9936
rect 34060 9920 34112 9926
rect 34060 9862 34112 9868
rect 34072 8498 34100 9862
rect 34256 9722 34284 9930
rect 34244 9716 34296 9722
rect 34244 9658 34296 9664
rect 34440 9586 34468 11478
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34520 11348 34572 11354
rect 34520 11290 34572 11296
rect 34532 11218 34560 11290
rect 34520 11212 34572 11218
rect 34520 11154 34572 11160
rect 34532 10810 34560 11154
rect 34980 11144 35032 11150
rect 34980 11086 35032 11092
rect 34704 11076 34756 11082
rect 34704 11018 34756 11024
rect 34520 10804 34572 10810
rect 34520 10746 34572 10752
rect 34520 10668 34572 10674
rect 34520 10610 34572 10616
rect 34532 10062 34560 10610
rect 34520 10056 34572 10062
rect 34520 9998 34572 10004
rect 34532 9654 34560 9998
rect 34520 9648 34572 9654
rect 34520 9590 34572 9596
rect 34716 9586 34744 11018
rect 34992 10742 35020 11086
rect 35348 11076 35400 11082
rect 35452 11064 35480 12718
rect 35532 12640 35584 12646
rect 35532 12582 35584 12588
rect 35544 12238 35572 12582
rect 35532 12232 35584 12238
rect 35532 12174 35584 12180
rect 35728 11898 35756 12854
rect 35716 11892 35768 11898
rect 35716 11834 35768 11840
rect 35820 11150 35848 14962
rect 35912 14346 35940 18566
rect 36728 18080 36780 18086
rect 36728 18022 36780 18028
rect 36740 17954 36768 18022
rect 36648 17926 36768 17954
rect 36648 17610 36676 17926
rect 36636 17604 36688 17610
rect 36636 17546 36688 17552
rect 36648 17513 36676 17546
rect 36634 17504 36690 17513
rect 36634 17439 36690 17448
rect 36636 16652 36688 16658
rect 36636 16594 36688 16600
rect 36544 15904 36596 15910
rect 36544 15846 36596 15852
rect 35992 15496 36044 15502
rect 35992 15438 36044 15444
rect 36004 15337 36032 15438
rect 36268 15360 36320 15366
rect 35990 15328 36046 15337
rect 36268 15302 36320 15308
rect 35990 15263 36046 15272
rect 35992 15156 36044 15162
rect 35992 15098 36044 15104
rect 36004 15065 36032 15098
rect 36280 15094 36308 15302
rect 36268 15088 36320 15094
rect 35990 15056 36046 15065
rect 36268 15030 36320 15036
rect 35990 14991 36046 15000
rect 36452 15020 36504 15026
rect 36452 14962 36504 14968
rect 35900 14340 35952 14346
rect 35900 14282 35952 14288
rect 36464 14074 36492 14962
rect 36452 14068 36504 14074
rect 36452 14010 36504 14016
rect 35900 13932 35952 13938
rect 35900 13874 35952 13880
rect 35992 13932 36044 13938
rect 35992 13874 36044 13880
rect 35912 12850 35940 13874
rect 36004 13530 36032 13874
rect 35992 13524 36044 13530
rect 35992 13466 36044 13472
rect 35992 13252 36044 13258
rect 35992 13194 36044 13200
rect 35900 12844 35952 12850
rect 35900 12786 35952 12792
rect 35808 11144 35860 11150
rect 35808 11086 35860 11092
rect 35400 11036 35480 11064
rect 35348 11018 35400 11024
rect 34980 10736 35032 10742
rect 34980 10678 35032 10684
rect 34796 10600 34848 10606
rect 34796 10542 34848 10548
rect 34808 10266 34836 10542
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34796 10260 34848 10266
rect 34796 10202 34848 10208
rect 34428 9580 34480 9586
rect 34428 9522 34480 9528
rect 34612 9580 34664 9586
rect 34612 9522 34664 9528
rect 34704 9580 34756 9586
rect 34704 9522 34756 9528
rect 34520 9512 34572 9518
rect 34520 9454 34572 9460
rect 34532 8838 34560 9454
rect 34624 9178 34652 9522
rect 34612 9172 34664 9178
rect 34612 9114 34664 9120
rect 34612 8968 34664 8974
rect 34612 8910 34664 8916
rect 34520 8832 34572 8838
rect 34520 8774 34572 8780
rect 34060 8492 34112 8498
rect 34060 8434 34112 8440
rect 34428 8492 34480 8498
rect 34428 8434 34480 8440
rect 33874 8392 33930 8401
rect 33874 8327 33876 8336
rect 33928 8327 33930 8336
rect 33876 8298 33928 8304
rect 33784 8016 33836 8022
rect 33784 7958 33836 7964
rect 33692 7948 33744 7954
rect 33692 7890 33744 7896
rect 32956 7880 33008 7886
rect 32956 7822 33008 7828
rect 32588 7744 32640 7750
rect 32588 7686 32640 7692
rect 32600 7478 32628 7686
rect 32588 7472 32640 7478
rect 32588 7414 32640 7420
rect 32968 6882 32996 7822
rect 32876 6854 32996 6882
rect 32876 6798 32904 6854
rect 32864 6792 32916 6798
rect 32864 6734 32916 6740
rect 32876 5370 32904 6734
rect 33600 6724 33652 6730
rect 33600 6666 33652 6672
rect 33612 6458 33640 6666
rect 33704 6458 33732 7890
rect 34244 7880 34296 7886
rect 33968 7874 34020 7880
rect 34244 7822 34296 7828
rect 33968 7816 34020 7822
rect 33980 7546 34008 7816
rect 33968 7540 34020 7546
rect 33968 7482 34020 7488
rect 34060 7200 34112 7206
rect 34060 7142 34112 7148
rect 33600 6452 33652 6458
rect 33600 6394 33652 6400
rect 33692 6452 33744 6458
rect 33692 6394 33744 6400
rect 34072 6322 34100 7142
rect 34256 6322 34284 7822
rect 34440 7410 34468 8434
rect 34532 8430 34560 8774
rect 34520 8424 34572 8430
rect 34520 8366 34572 8372
rect 34532 8090 34560 8366
rect 34520 8084 34572 8090
rect 34520 8026 34572 8032
rect 34428 7404 34480 7410
rect 34428 7346 34480 7352
rect 34440 7002 34468 7346
rect 34428 6996 34480 7002
rect 34428 6938 34480 6944
rect 34624 6798 34652 8910
rect 34716 8498 34744 9522
rect 34808 9042 34836 10202
rect 35360 10062 35388 11018
rect 35532 11008 35584 11014
rect 35532 10950 35584 10956
rect 35440 10736 35492 10742
rect 35440 10678 35492 10684
rect 35348 10056 35400 10062
rect 35348 9998 35400 10004
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 35256 9172 35308 9178
rect 35256 9114 35308 9120
rect 34796 9036 34848 9042
rect 34796 8978 34848 8984
rect 35268 8786 35296 9114
rect 35452 8974 35480 10678
rect 35544 10606 35572 10950
rect 35820 10674 35848 11086
rect 35808 10668 35860 10674
rect 35808 10610 35860 10616
rect 35532 10600 35584 10606
rect 35532 10542 35584 10548
rect 35544 9450 35572 10542
rect 35820 10062 35848 10610
rect 35716 10056 35768 10062
rect 35716 9998 35768 10004
rect 35808 10056 35860 10062
rect 35808 9998 35860 10004
rect 35728 9586 35756 9998
rect 35716 9580 35768 9586
rect 35716 9522 35768 9528
rect 35624 9512 35676 9518
rect 35624 9454 35676 9460
rect 35532 9444 35584 9450
rect 35532 9386 35584 9392
rect 35440 8968 35492 8974
rect 35440 8910 35492 8916
rect 35268 8758 35388 8786
rect 34796 8560 34848 8566
rect 34796 8502 34848 8508
rect 34704 8492 34756 8498
rect 34704 8434 34756 8440
rect 34612 6792 34664 6798
rect 34612 6734 34664 6740
rect 34612 6656 34664 6662
rect 34612 6598 34664 6604
rect 34704 6656 34756 6662
rect 34704 6598 34756 6604
rect 34624 6322 34652 6598
rect 33876 6316 33928 6322
rect 33876 6258 33928 6264
rect 34060 6316 34112 6322
rect 34060 6258 34112 6264
rect 34244 6316 34296 6322
rect 34244 6258 34296 6264
rect 34612 6316 34664 6322
rect 34612 6258 34664 6264
rect 32864 5364 32916 5370
rect 32864 5306 32916 5312
rect 33888 5234 33916 6258
rect 34624 5370 34652 6258
rect 34716 5574 34744 6598
rect 34704 5568 34756 5574
rect 34704 5510 34756 5516
rect 34612 5364 34664 5370
rect 34612 5306 34664 5312
rect 33324 5228 33376 5234
rect 33324 5170 33376 5176
rect 33876 5228 33928 5234
rect 33876 5170 33928 5176
rect 34428 5228 34480 5234
rect 34428 5170 34480 5176
rect 32864 5024 32916 5030
rect 32864 4966 32916 4972
rect 32404 4616 32456 4622
rect 32404 4558 32456 4564
rect 27896 4140 27948 4146
rect 27896 4082 27948 4088
rect 30840 4140 30892 4146
rect 30840 4082 30892 4088
rect 27804 4004 27856 4010
rect 27804 3946 27856 3952
rect 32416 3738 32444 4558
rect 32588 3936 32640 3942
rect 32588 3878 32640 3884
rect 27712 3732 27764 3738
rect 27712 3674 27764 3680
rect 32404 3732 32456 3738
rect 32404 3674 32456 3680
rect 27344 3596 27396 3602
rect 27344 3538 27396 3544
rect 26700 3528 26752 3534
rect 26700 3470 26752 3476
rect 26792 3528 26844 3534
rect 26792 3470 26844 3476
rect 26976 3528 27028 3534
rect 26976 3470 27028 3476
rect 27896 3528 27948 3534
rect 27896 3470 27948 3476
rect 28724 3528 28776 3534
rect 28724 3470 28776 3476
rect 29552 3528 29604 3534
rect 29552 3470 29604 3476
rect 30656 3528 30708 3534
rect 30656 3470 30708 3476
rect 31208 3528 31260 3534
rect 31208 3470 31260 3476
rect 26988 3194 27016 3470
rect 26424 3188 26476 3194
rect 26424 3130 26476 3136
rect 26976 3188 27028 3194
rect 26976 3130 27028 3136
rect 26330 2952 26386 2961
rect 26330 2887 26386 2896
rect 27068 2916 27120 2922
rect 27068 2858 27120 2864
rect 26792 2848 26844 2854
rect 26792 2790 26844 2796
rect 26516 2508 26568 2514
rect 26516 2450 26568 2456
rect 26528 800 26556 2450
rect 26804 800 26832 2790
rect 27080 800 27108 2858
rect 27344 2576 27396 2582
rect 27344 2518 27396 2524
rect 27356 800 27384 2518
rect 27620 2440 27672 2446
rect 27620 2382 27672 2388
rect 27632 800 27660 2382
rect 27908 800 27936 3470
rect 28172 2848 28224 2854
rect 28172 2790 28224 2796
rect 28184 800 28212 2790
rect 28448 2508 28500 2514
rect 28448 2450 28500 2456
rect 28460 800 28488 2450
rect 28736 800 28764 3470
rect 29000 2984 29052 2990
rect 29000 2926 29052 2932
rect 29012 800 29040 2926
rect 29276 2848 29328 2854
rect 29276 2790 29328 2796
rect 29288 800 29316 2790
rect 29564 800 29592 3470
rect 30104 2848 30156 2854
rect 30104 2790 30156 2796
rect 29828 2440 29880 2446
rect 29828 2382 29880 2388
rect 29840 800 29868 2382
rect 30116 800 30144 2790
rect 30380 2508 30432 2514
rect 30380 2450 30432 2456
rect 30392 800 30420 2450
rect 30668 800 30696 3470
rect 30932 2984 30984 2990
rect 30932 2926 30984 2932
rect 30944 800 30972 2926
rect 31220 800 31248 3470
rect 31484 2848 31536 2854
rect 31484 2790 31536 2796
rect 32036 2848 32088 2854
rect 32036 2790 32088 2796
rect 31496 800 31524 2790
rect 31760 2372 31812 2378
rect 31760 2314 31812 2320
rect 31772 800 31800 2314
rect 32048 800 32076 2790
rect 32312 2440 32364 2446
rect 32312 2382 32364 2388
rect 32324 800 32352 2382
rect 32600 800 32628 3878
rect 32876 3534 32904 4966
rect 33336 4826 33364 5170
rect 33784 5024 33836 5030
rect 33784 4966 33836 4972
rect 33324 4820 33376 4826
rect 33324 4762 33376 4768
rect 33796 4146 33824 4966
rect 33888 4826 33916 5170
rect 34440 4826 34468 5170
rect 33876 4820 33928 4826
rect 33876 4762 33928 4768
rect 34428 4820 34480 4826
rect 34428 4762 34480 4768
rect 34716 4554 34744 5510
rect 34808 4622 34836 8502
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 35164 6724 35216 6730
rect 35164 6666 35216 6672
rect 35176 6458 35204 6666
rect 35164 6452 35216 6458
rect 35164 6394 35216 6400
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 35360 5234 35388 8758
rect 35440 6316 35492 6322
rect 35440 6258 35492 6264
rect 35452 5914 35480 6258
rect 35440 5908 35492 5914
rect 35440 5850 35492 5856
rect 35544 5710 35572 9386
rect 35636 8974 35664 9454
rect 35912 9382 35940 12786
rect 36004 12170 36032 13194
rect 36556 12714 36584 15846
rect 36648 14278 36676 16594
rect 37108 15706 37136 18906
rect 37280 18896 37332 18902
rect 37280 18838 37332 18844
rect 37292 17882 37320 18838
rect 37384 18630 37412 19246
rect 37372 18624 37424 18630
rect 37372 18566 37424 18572
rect 37280 17876 37332 17882
rect 37280 17818 37332 17824
rect 37384 17814 37412 18566
rect 37476 18358 37504 19722
rect 37556 19372 37608 19378
rect 37556 19314 37608 19320
rect 37568 18766 37596 19314
rect 37556 18760 37608 18766
rect 37556 18702 37608 18708
rect 37464 18352 37516 18358
rect 37464 18294 37516 18300
rect 37372 17808 37424 17814
rect 37372 17750 37424 17756
rect 37384 17202 37412 17750
rect 37476 17678 37504 18294
rect 37464 17672 37516 17678
rect 37464 17614 37516 17620
rect 37372 17196 37424 17202
rect 37372 17138 37424 17144
rect 37280 16992 37332 16998
rect 37280 16934 37332 16940
rect 37292 16794 37320 16934
rect 37280 16788 37332 16794
rect 37280 16730 37332 16736
rect 37660 16182 37688 19722
rect 37740 19712 37792 19718
rect 37740 19654 37792 19660
rect 37752 19378 37780 19654
rect 38212 19378 38240 20266
rect 38304 19514 38332 20402
rect 65654 20156 65962 20165
rect 65654 20154 65660 20156
rect 65716 20154 65740 20156
rect 65796 20154 65820 20156
rect 65876 20154 65900 20156
rect 65956 20154 65962 20156
rect 65716 20102 65718 20154
rect 65898 20102 65900 20154
rect 65654 20100 65660 20102
rect 65716 20100 65740 20102
rect 65796 20100 65820 20102
rect 65876 20100 65900 20102
rect 65956 20100 65962 20102
rect 65654 20091 65962 20100
rect 39028 19848 39080 19854
rect 68100 19848 68152 19854
rect 39028 19790 39080 19796
rect 68098 19816 68100 19825
rect 68152 19816 68154 19825
rect 38292 19508 38344 19514
rect 38292 19450 38344 19456
rect 37740 19372 37792 19378
rect 37740 19314 37792 19320
rect 38200 19372 38252 19378
rect 38200 19314 38252 19320
rect 37924 19168 37976 19174
rect 37924 19110 37976 19116
rect 37832 18760 37884 18766
rect 37832 18702 37884 18708
rect 37844 17678 37872 18702
rect 37936 18290 37964 19110
rect 38108 18692 38160 18698
rect 38108 18634 38160 18640
rect 38120 18426 38148 18634
rect 38108 18420 38160 18426
rect 38108 18362 38160 18368
rect 37924 18284 37976 18290
rect 37924 18226 37976 18232
rect 37832 17672 37884 17678
rect 37832 17614 37884 17620
rect 37740 17604 37792 17610
rect 37740 17546 37792 17552
rect 37752 17338 37780 17546
rect 37740 17332 37792 17338
rect 37740 17274 37792 17280
rect 37752 16522 37780 17274
rect 37844 17202 37872 17614
rect 37832 17196 37884 17202
rect 37832 17138 37884 17144
rect 37936 16561 37964 18226
rect 38016 17672 38068 17678
rect 38014 17640 38016 17649
rect 38068 17640 38070 17649
rect 38014 17575 38070 17584
rect 38108 17060 38160 17066
rect 38108 17002 38160 17008
rect 38120 16794 38148 17002
rect 38108 16788 38160 16794
rect 38108 16730 38160 16736
rect 37922 16552 37978 16561
rect 37740 16516 37792 16522
rect 37740 16458 37792 16464
rect 37832 16516 37884 16522
rect 37922 16487 37978 16496
rect 37832 16458 37884 16464
rect 37752 16250 37780 16458
rect 37740 16244 37792 16250
rect 37740 16186 37792 16192
rect 37648 16176 37700 16182
rect 37648 16118 37700 16124
rect 37464 16108 37516 16114
rect 37464 16050 37516 16056
rect 37096 15700 37148 15706
rect 37096 15642 37148 15648
rect 37280 15496 37332 15502
rect 37332 15444 37412 15450
rect 37280 15438 37412 15444
rect 37292 15422 37412 15438
rect 37476 15434 37504 16050
rect 37648 16040 37700 16046
rect 37648 15982 37700 15988
rect 37660 15638 37688 15982
rect 37740 15700 37792 15706
rect 37740 15642 37792 15648
rect 37648 15632 37700 15638
rect 37648 15574 37700 15580
rect 37384 15162 37412 15422
rect 37464 15428 37516 15434
rect 37464 15370 37516 15376
rect 37372 15156 37424 15162
rect 37372 15098 37424 15104
rect 36728 14952 36780 14958
rect 36728 14894 36780 14900
rect 36636 14272 36688 14278
rect 36636 14214 36688 14220
rect 36648 13938 36676 14214
rect 36740 14006 36768 14894
rect 36912 14884 36964 14890
rect 36912 14826 36964 14832
rect 36820 14340 36872 14346
rect 36820 14282 36872 14288
rect 36728 14000 36780 14006
rect 36728 13942 36780 13948
rect 36636 13932 36688 13938
rect 36636 13874 36688 13880
rect 36832 13394 36860 14282
rect 36820 13388 36872 13394
rect 36820 13330 36872 13336
rect 36924 13326 36952 14826
rect 37280 14408 37332 14414
rect 37280 14350 37332 14356
rect 36912 13320 36964 13326
rect 36912 13262 36964 13268
rect 37292 12782 37320 14350
rect 37384 13938 37412 15098
rect 37476 14822 37504 15370
rect 37556 15020 37608 15026
rect 37556 14962 37608 14968
rect 37464 14816 37516 14822
rect 37464 14758 37516 14764
rect 37476 14414 37504 14758
rect 37464 14408 37516 14414
rect 37464 14350 37516 14356
rect 37372 13932 37424 13938
rect 37372 13874 37424 13880
rect 37280 12776 37332 12782
rect 37280 12718 37332 12724
rect 36544 12708 36596 12714
rect 36544 12650 36596 12656
rect 37292 12306 37320 12718
rect 37280 12300 37332 12306
rect 37280 12242 37332 12248
rect 35992 12164 36044 12170
rect 35992 12106 36044 12112
rect 37188 12164 37240 12170
rect 37188 12106 37240 12112
rect 36912 11552 36964 11558
rect 36912 11494 36964 11500
rect 36820 10532 36872 10538
rect 36820 10474 36872 10480
rect 35900 9376 35952 9382
rect 35900 9318 35952 9324
rect 35716 9036 35768 9042
rect 35716 8978 35768 8984
rect 35624 8968 35676 8974
rect 35624 8910 35676 8916
rect 35728 8498 35756 8978
rect 35716 8492 35768 8498
rect 35716 8434 35768 8440
rect 35992 8424 36044 8430
rect 35992 8366 36044 8372
rect 35900 8356 35952 8362
rect 35900 8298 35952 8304
rect 35912 7478 35940 8298
rect 36004 7818 36032 8366
rect 36176 7948 36228 7954
rect 36176 7890 36228 7896
rect 35992 7812 36044 7818
rect 35992 7754 36044 7760
rect 35900 7472 35952 7478
rect 35900 7414 35952 7420
rect 35808 6724 35860 6730
rect 35808 6666 35860 6672
rect 35532 5704 35584 5710
rect 35532 5646 35584 5652
rect 35820 5522 35848 6666
rect 36004 6458 36032 7754
rect 36188 7478 36216 7890
rect 36176 7472 36228 7478
rect 36176 7414 36228 7420
rect 36084 7404 36136 7410
rect 36084 7346 36136 7352
rect 36360 7404 36412 7410
rect 36360 7346 36412 7352
rect 35992 6452 36044 6458
rect 35992 6394 36044 6400
rect 35992 5908 36044 5914
rect 35992 5850 36044 5856
rect 35820 5494 35940 5522
rect 35348 5228 35400 5234
rect 35348 5170 35400 5176
rect 35624 5024 35676 5030
rect 35624 4966 35676 4972
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34796 4616 34848 4622
rect 34796 4558 34848 4564
rect 34704 4548 34756 4554
rect 34704 4490 34756 4496
rect 34808 4282 34836 4558
rect 34796 4276 34848 4282
rect 34796 4218 34848 4224
rect 35636 4146 35664 4966
rect 35912 4214 35940 5494
rect 36004 5234 36032 5850
rect 35992 5228 36044 5234
rect 35992 5170 36044 5176
rect 36096 4622 36124 7346
rect 36372 7002 36400 7346
rect 36360 6996 36412 7002
rect 36360 6938 36412 6944
rect 36372 6390 36400 6938
rect 36832 6662 36860 10474
rect 36924 10266 36952 11494
rect 37096 11144 37148 11150
rect 37096 11086 37148 11092
rect 36912 10260 36964 10266
rect 36912 10202 36964 10208
rect 37108 10062 37136 11086
rect 37096 10056 37148 10062
rect 37096 9998 37148 10004
rect 37004 9988 37056 9994
rect 37004 9930 37056 9936
rect 37016 8974 37044 9930
rect 37108 9042 37136 9998
rect 37200 9518 37228 12106
rect 37384 11898 37412 13874
rect 37568 13530 37596 14962
rect 37660 14550 37688 15574
rect 37752 15026 37780 15642
rect 37740 15020 37792 15026
rect 37740 14962 37792 14968
rect 37648 14544 37700 14550
rect 37648 14486 37700 14492
rect 37740 14272 37792 14278
rect 37740 14214 37792 14220
rect 37752 14074 37780 14214
rect 37740 14068 37792 14074
rect 37740 14010 37792 14016
rect 37844 13734 37872 16458
rect 38212 16114 38240 19314
rect 39040 19310 39068 19790
rect 68098 19751 68154 19760
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 39212 19372 39264 19378
rect 39212 19314 39264 19320
rect 39028 19304 39080 19310
rect 39028 19246 39080 19252
rect 38936 18964 38988 18970
rect 38936 18906 38988 18912
rect 38948 18766 38976 18906
rect 39040 18834 39068 19246
rect 39224 18970 39252 19314
rect 65654 19068 65962 19077
rect 65654 19066 65660 19068
rect 65716 19066 65740 19068
rect 65796 19066 65820 19068
rect 65876 19066 65900 19068
rect 65956 19066 65962 19068
rect 65716 19014 65718 19066
rect 65898 19014 65900 19066
rect 65654 19012 65660 19014
rect 65716 19012 65740 19014
rect 65796 19012 65820 19014
rect 65876 19012 65900 19014
rect 65956 19012 65962 19014
rect 65654 19003 65962 19012
rect 39212 18964 39264 18970
rect 39212 18906 39264 18912
rect 39028 18828 39080 18834
rect 39028 18770 39080 18776
rect 38936 18760 38988 18766
rect 38936 18702 38988 18708
rect 38660 18284 38712 18290
rect 38660 18226 38712 18232
rect 38672 17882 38700 18226
rect 39040 18222 39068 18770
rect 68100 18760 68152 18766
rect 68100 18702 68152 18708
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 68112 18465 68140 18702
rect 68098 18456 68154 18465
rect 68098 18391 68154 18400
rect 39028 18216 39080 18222
rect 39028 18158 39080 18164
rect 38292 17876 38344 17882
rect 38292 17818 38344 17824
rect 38660 17876 38712 17882
rect 38660 17818 38712 17824
rect 38200 16108 38252 16114
rect 38200 16050 38252 16056
rect 38304 15994 38332 17818
rect 38752 17672 38804 17678
rect 38752 17614 38804 17620
rect 38384 17196 38436 17202
rect 38384 17138 38436 17144
rect 38396 16726 38424 17138
rect 38384 16720 38436 16726
rect 38384 16662 38436 16668
rect 38212 15966 38332 15994
rect 38016 14884 38068 14890
rect 38016 14826 38068 14832
rect 37924 14544 37976 14550
rect 37924 14486 37976 14492
rect 37832 13728 37884 13734
rect 37832 13670 37884 13676
rect 37556 13524 37608 13530
rect 37556 13466 37608 13472
rect 37556 13320 37608 13326
rect 37556 13262 37608 13268
rect 37568 12850 37596 13262
rect 37556 12844 37608 12850
rect 37556 12786 37608 12792
rect 37568 12238 37596 12786
rect 37832 12640 37884 12646
rect 37832 12582 37884 12588
rect 37844 12238 37872 12582
rect 37464 12232 37516 12238
rect 37464 12174 37516 12180
rect 37556 12232 37608 12238
rect 37556 12174 37608 12180
rect 37832 12232 37884 12238
rect 37832 12174 37884 12180
rect 37372 11892 37424 11898
rect 37372 11834 37424 11840
rect 37280 11552 37332 11558
rect 37280 11494 37332 11500
rect 37292 11150 37320 11494
rect 37280 11144 37332 11150
rect 37280 11086 37332 11092
rect 37280 11008 37332 11014
rect 37280 10950 37332 10956
rect 37292 9994 37320 10950
rect 37384 10470 37412 11834
rect 37476 11762 37504 12174
rect 37464 11756 37516 11762
rect 37464 11698 37516 11704
rect 37476 10674 37504 11698
rect 37464 10668 37516 10674
rect 37464 10610 37516 10616
rect 37372 10464 37424 10470
rect 37372 10406 37424 10412
rect 37280 9988 37332 9994
rect 37280 9930 37332 9936
rect 37372 9920 37424 9926
rect 37372 9862 37424 9868
rect 37188 9512 37240 9518
rect 37188 9454 37240 9460
rect 37188 9376 37240 9382
rect 37188 9318 37240 9324
rect 37096 9036 37148 9042
rect 37096 8978 37148 8984
rect 37004 8968 37056 8974
rect 37004 8910 37056 8916
rect 37016 7954 37044 8910
rect 37108 8498 37136 8978
rect 37200 8956 37228 9318
rect 37280 8968 37332 8974
rect 37200 8928 37280 8956
rect 37280 8910 37332 8916
rect 37384 8786 37412 9862
rect 37568 9586 37596 12174
rect 37936 11694 37964 14486
rect 38028 14414 38056 14826
rect 38016 14408 38068 14414
rect 38016 14350 38068 14356
rect 38016 13728 38068 13734
rect 38016 13670 38068 13676
rect 38028 13326 38056 13670
rect 38016 13320 38068 13326
rect 38016 13262 38068 13268
rect 38108 13184 38160 13190
rect 38108 13126 38160 13132
rect 38016 12232 38068 12238
rect 38016 12174 38068 12180
rect 38028 11762 38056 12174
rect 38120 12170 38148 13126
rect 38212 12238 38240 15966
rect 38292 14272 38344 14278
rect 38292 14214 38344 14220
rect 38304 14006 38332 14214
rect 38292 14000 38344 14006
rect 38292 13942 38344 13948
rect 38292 13524 38344 13530
rect 38292 13466 38344 13472
rect 38304 13326 38332 13466
rect 38292 13320 38344 13326
rect 38292 13262 38344 13268
rect 38200 12232 38252 12238
rect 38200 12174 38252 12180
rect 38108 12164 38160 12170
rect 38108 12106 38160 12112
rect 38016 11756 38068 11762
rect 38016 11698 38068 11704
rect 37924 11688 37976 11694
rect 37924 11630 37976 11636
rect 37936 10606 37964 11630
rect 38028 11354 38056 11698
rect 38016 11348 38068 11354
rect 38016 11290 38068 11296
rect 38396 11014 38424 16662
rect 38660 15904 38712 15910
rect 38660 15846 38712 15852
rect 38672 15434 38700 15846
rect 38476 15428 38528 15434
rect 38476 15370 38528 15376
rect 38660 15428 38712 15434
rect 38660 15370 38712 15376
rect 38488 15162 38516 15370
rect 38476 15156 38528 15162
rect 38476 15098 38528 15104
rect 38672 15094 38700 15370
rect 38660 15088 38712 15094
rect 38660 15030 38712 15036
rect 38764 13462 38792 17614
rect 38844 17604 38896 17610
rect 38844 17546 38896 17552
rect 38856 17338 38884 17546
rect 38844 17332 38896 17338
rect 38844 17274 38896 17280
rect 39040 17202 39068 18158
rect 40408 18080 40460 18086
rect 40408 18022 40460 18028
rect 40420 17678 40448 18022
rect 65654 17980 65962 17989
rect 65654 17978 65660 17980
rect 65716 17978 65740 17980
rect 65796 17978 65820 17980
rect 65876 17978 65900 17980
rect 65956 17978 65962 17980
rect 65716 17926 65718 17978
rect 65898 17926 65900 17978
rect 65654 17924 65660 17926
rect 65716 17924 65740 17926
rect 65796 17924 65820 17926
rect 65876 17924 65900 17926
rect 65956 17924 65962 17926
rect 65654 17915 65962 17924
rect 40408 17672 40460 17678
rect 39302 17640 39358 17649
rect 40408 17614 40460 17620
rect 39302 17575 39304 17584
rect 39356 17575 39358 17584
rect 39304 17546 39356 17552
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 39028 17196 39080 17202
rect 39028 17138 39080 17144
rect 67638 17096 67694 17105
rect 67638 17031 67640 17040
rect 67692 17031 67694 17040
rect 67640 17002 67692 17008
rect 40592 16992 40644 16998
rect 40592 16934 40644 16940
rect 40604 16522 40632 16934
rect 65654 16892 65962 16901
rect 65654 16890 65660 16892
rect 65716 16890 65740 16892
rect 65796 16890 65820 16892
rect 65876 16890 65900 16892
rect 65956 16890 65962 16892
rect 65716 16838 65718 16890
rect 65898 16838 65900 16890
rect 65654 16836 65660 16838
rect 65716 16836 65740 16838
rect 65796 16836 65820 16838
rect 65876 16836 65900 16838
rect 65956 16836 65962 16838
rect 65654 16827 65962 16836
rect 40592 16516 40644 16522
rect 40592 16458 40644 16464
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 38844 16108 38896 16114
rect 38844 16050 38896 16056
rect 38856 15706 38884 16050
rect 41236 16040 41288 16046
rect 41236 15982 41288 15988
rect 38844 15700 38896 15706
rect 38844 15642 38896 15648
rect 41248 15570 41276 15982
rect 67640 15904 67692 15910
rect 67640 15846 67692 15852
rect 65654 15804 65962 15813
rect 65654 15802 65660 15804
rect 65716 15802 65740 15804
rect 65796 15802 65820 15804
rect 65876 15802 65900 15804
rect 65956 15802 65962 15804
rect 65716 15750 65718 15802
rect 65898 15750 65900 15802
rect 65654 15748 65660 15750
rect 65716 15748 65740 15750
rect 65796 15748 65820 15750
rect 65876 15748 65900 15750
rect 65956 15748 65962 15750
rect 65654 15739 65962 15748
rect 67652 15745 67680 15846
rect 67638 15736 67694 15745
rect 67638 15671 67694 15680
rect 41236 15564 41288 15570
rect 41236 15506 41288 15512
rect 38934 15328 38990 15337
rect 38934 15263 38990 15272
rect 38948 14414 38976 15263
rect 38936 14408 38988 14414
rect 38936 14350 38988 14356
rect 38844 14340 38896 14346
rect 38844 14282 38896 14288
rect 38752 13456 38804 13462
rect 38752 13398 38804 13404
rect 38752 13320 38804 13326
rect 38752 13262 38804 13268
rect 38476 13184 38528 13190
rect 38476 13126 38528 13132
rect 38488 12918 38516 13126
rect 38476 12912 38528 12918
rect 38476 12854 38528 12860
rect 38660 12844 38712 12850
rect 38660 12786 38712 12792
rect 38672 12102 38700 12786
rect 38660 12096 38712 12102
rect 38660 12038 38712 12044
rect 38672 11150 38700 12038
rect 38660 11144 38712 11150
rect 38660 11086 38712 11092
rect 38384 11008 38436 11014
rect 38384 10950 38436 10956
rect 38396 10674 38424 10950
rect 38016 10668 38068 10674
rect 38016 10610 38068 10616
rect 38200 10668 38252 10674
rect 38200 10610 38252 10616
rect 38384 10668 38436 10674
rect 38384 10610 38436 10616
rect 37924 10600 37976 10606
rect 37924 10542 37976 10548
rect 37924 10464 37976 10470
rect 37924 10406 37976 10412
rect 37740 10056 37792 10062
rect 37740 9998 37792 10004
rect 37556 9580 37608 9586
rect 37556 9522 37608 9528
rect 37292 8758 37412 8786
rect 37464 8832 37516 8838
rect 37464 8774 37516 8780
rect 37096 8492 37148 8498
rect 37096 8434 37148 8440
rect 37004 7948 37056 7954
rect 37004 7890 37056 7896
rect 37016 6866 37044 7890
rect 37108 7342 37136 8434
rect 37292 8430 37320 8758
rect 37280 8424 37332 8430
rect 37280 8366 37332 8372
rect 37292 8090 37320 8366
rect 37280 8084 37332 8090
rect 37280 8026 37332 8032
rect 37372 7880 37424 7886
rect 37372 7822 37424 7828
rect 37384 7546 37412 7822
rect 37372 7540 37424 7546
rect 37372 7482 37424 7488
rect 37096 7336 37148 7342
rect 37096 7278 37148 7284
rect 37004 6860 37056 6866
rect 37004 6802 37056 6808
rect 37108 6798 37136 7278
rect 37096 6792 37148 6798
rect 37096 6734 37148 6740
rect 36820 6656 36872 6662
rect 36820 6598 36872 6604
rect 36360 6384 36412 6390
rect 36360 6326 36412 6332
rect 37372 6316 37424 6322
rect 37372 6258 37424 6264
rect 37188 6180 37240 6186
rect 37188 6122 37240 6128
rect 37200 5778 37228 6122
rect 37188 5772 37240 5778
rect 37188 5714 37240 5720
rect 36452 5704 36504 5710
rect 36452 5646 36504 5652
rect 36464 5234 36492 5646
rect 37200 5302 37228 5714
rect 37280 5704 37332 5710
rect 37280 5646 37332 5652
rect 37292 5370 37320 5646
rect 37384 5574 37412 6258
rect 37372 5568 37424 5574
rect 37372 5510 37424 5516
rect 37280 5364 37332 5370
rect 37280 5306 37332 5312
rect 37188 5296 37240 5302
rect 37188 5238 37240 5244
rect 37384 5234 37412 5510
rect 37476 5302 37504 8774
rect 37568 7886 37596 9522
rect 37752 9364 37780 9998
rect 37936 9994 37964 10406
rect 37924 9988 37976 9994
rect 37924 9930 37976 9936
rect 38028 9738 38056 10610
rect 38108 10464 38160 10470
rect 38108 10406 38160 10412
rect 38120 10062 38148 10406
rect 38212 10266 38240 10610
rect 38200 10260 38252 10266
rect 38200 10202 38252 10208
rect 38108 10056 38160 10062
rect 38108 9998 38160 10004
rect 38028 9710 38148 9738
rect 38016 9580 38068 9586
rect 38016 9522 38068 9528
rect 37832 9376 37884 9382
rect 37752 9336 37832 9364
rect 37832 9318 37884 9324
rect 37844 8974 37872 9318
rect 38028 9178 38056 9522
rect 38016 9172 38068 9178
rect 38016 9114 38068 9120
rect 38120 9058 38148 9710
rect 38396 9654 38424 10610
rect 38384 9648 38436 9654
rect 38384 9590 38436 9596
rect 38028 9030 38148 9058
rect 37832 8968 37884 8974
rect 37832 8910 37884 8916
rect 37556 7880 37608 7886
rect 37556 7822 37608 7828
rect 37924 7880 37976 7886
rect 37924 7822 37976 7828
rect 37936 7410 37964 7822
rect 37924 7404 37976 7410
rect 37924 7346 37976 7352
rect 38028 6882 38056 9030
rect 38568 8900 38620 8906
rect 38568 8842 38620 8848
rect 38580 8362 38608 8842
rect 38764 8566 38792 13262
rect 38856 12850 38884 14282
rect 38948 12986 38976 14350
rect 39120 14272 39172 14278
rect 39120 14214 39172 14220
rect 39132 13734 39160 14214
rect 41248 13938 41276 15506
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 65654 14716 65962 14725
rect 65654 14714 65660 14716
rect 65716 14714 65740 14716
rect 65796 14714 65820 14716
rect 65876 14714 65900 14716
rect 65956 14714 65962 14716
rect 65716 14662 65718 14714
rect 65898 14662 65900 14714
rect 65654 14660 65660 14662
rect 65716 14660 65740 14662
rect 65796 14660 65820 14662
rect 65876 14660 65900 14662
rect 65956 14660 65962 14662
rect 65654 14651 65962 14660
rect 68100 14408 68152 14414
rect 68098 14376 68100 14385
rect 68152 14376 68154 14385
rect 68098 14311 68154 14320
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 41236 13932 41288 13938
rect 41236 13874 41288 13880
rect 39120 13728 39172 13734
rect 39120 13670 39172 13676
rect 41248 13190 41276 13874
rect 65654 13628 65962 13637
rect 65654 13626 65660 13628
rect 65716 13626 65740 13628
rect 65796 13626 65820 13628
rect 65876 13626 65900 13628
rect 65956 13626 65962 13628
rect 65716 13574 65718 13626
rect 65898 13574 65900 13626
rect 65654 13572 65660 13574
rect 65716 13572 65740 13574
rect 65796 13572 65820 13574
rect 65876 13572 65900 13574
rect 65956 13572 65962 13574
rect 65654 13563 65962 13572
rect 68100 13320 68152 13326
rect 68100 13262 68152 13268
rect 41236 13184 41288 13190
rect 41236 13126 41288 13132
rect 38936 12980 38988 12986
rect 38936 12922 38988 12928
rect 41248 12850 41276 13126
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 68112 13025 68140 13262
rect 68098 13016 68154 13025
rect 68098 12951 68154 12960
rect 38844 12844 38896 12850
rect 38844 12786 38896 12792
rect 41236 12844 41288 12850
rect 41236 12786 41288 12792
rect 41248 12238 41276 12786
rect 65654 12540 65962 12549
rect 65654 12538 65660 12540
rect 65716 12538 65740 12540
rect 65796 12538 65820 12540
rect 65876 12538 65900 12540
rect 65956 12538 65962 12540
rect 65716 12486 65718 12538
rect 65898 12486 65900 12538
rect 65654 12484 65660 12486
rect 65716 12484 65740 12486
rect 65796 12484 65820 12486
rect 65876 12484 65900 12486
rect 65956 12484 65962 12486
rect 65654 12475 65962 12484
rect 40500 12232 40552 12238
rect 40500 12174 40552 12180
rect 41236 12232 41288 12238
rect 41236 12174 41288 12180
rect 40512 11762 40540 12174
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 40500 11756 40552 11762
rect 40500 11698 40552 11704
rect 40512 10674 40540 11698
rect 67638 11656 67694 11665
rect 67638 11591 67640 11600
rect 67692 11591 67694 11600
rect 67640 11562 67692 11568
rect 65654 11452 65962 11461
rect 65654 11450 65660 11452
rect 65716 11450 65740 11452
rect 65796 11450 65820 11452
rect 65876 11450 65900 11452
rect 65956 11450 65962 11452
rect 65716 11398 65718 11450
rect 65898 11398 65900 11450
rect 65654 11396 65660 11398
rect 65716 11396 65740 11398
rect 65796 11396 65820 11398
rect 65876 11396 65900 11398
rect 65956 11396 65962 11398
rect 65654 11387 65962 11396
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 40500 10668 40552 10674
rect 40500 10610 40552 10616
rect 67640 10464 67692 10470
rect 67640 10406 67692 10412
rect 65654 10364 65962 10373
rect 65654 10362 65660 10364
rect 65716 10362 65740 10364
rect 65796 10362 65820 10364
rect 65876 10362 65900 10364
rect 65956 10362 65962 10364
rect 65716 10310 65718 10362
rect 65898 10310 65900 10362
rect 65654 10308 65660 10310
rect 65716 10308 65740 10310
rect 65796 10308 65820 10310
rect 65876 10308 65900 10310
rect 65956 10308 65962 10310
rect 65654 10299 65962 10308
rect 67652 10305 67680 10406
rect 67638 10296 67694 10305
rect 67638 10231 67694 10240
rect 39028 10124 39080 10130
rect 39028 10066 39080 10072
rect 39040 9586 39068 10066
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 39028 9580 39080 9586
rect 39028 9522 39080 9528
rect 38844 8832 38896 8838
rect 38844 8774 38896 8780
rect 38752 8560 38804 8566
rect 38752 8502 38804 8508
rect 38568 8356 38620 8362
rect 38568 8298 38620 8304
rect 38292 7880 38344 7886
rect 38292 7822 38344 7828
rect 38200 7268 38252 7274
rect 38200 7210 38252 7216
rect 38212 7002 38240 7210
rect 38200 6996 38252 7002
rect 38200 6938 38252 6944
rect 38028 6854 38148 6882
rect 37648 6656 37700 6662
rect 37648 6598 37700 6604
rect 37660 6390 37688 6598
rect 37648 6384 37700 6390
rect 37648 6326 37700 6332
rect 38120 6322 38148 6854
rect 38108 6316 38160 6322
rect 38108 6258 38160 6264
rect 38120 5642 38148 6258
rect 38304 5778 38332 7822
rect 38384 7744 38436 7750
rect 38384 7686 38436 7692
rect 38396 7342 38424 7686
rect 38476 7540 38528 7546
rect 38476 7482 38528 7488
rect 38488 7410 38516 7482
rect 38476 7404 38528 7410
rect 38476 7346 38528 7352
rect 38384 7336 38436 7342
rect 38384 7278 38436 7284
rect 38488 6322 38516 7346
rect 38580 6798 38608 8298
rect 38764 7546 38792 8502
rect 38856 7954 38884 8774
rect 39040 8634 39068 9522
rect 65654 9276 65962 9285
rect 65654 9274 65660 9276
rect 65716 9274 65740 9276
rect 65796 9274 65820 9276
rect 65876 9274 65900 9276
rect 65956 9274 65962 9276
rect 65716 9222 65718 9274
rect 65898 9222 65900 9274
rect 65654 9220 65660 9222
rect 65716 9220 65740 9222
rect 65796 9220 65820 9222
rect 65876 9220 65900 9222
rect 65956 9220 65962 9222
rect 65654 9211 65962 9220
rect 68100 8968 68152 8974
rect 68098 8936 68100 8945
rect 68152 8936 68154 8945
rect 41236 8900 41288 8906
rect 68098 8871 68154 8880
rect 41236 8842 41288 8848
rect 39028 8628 39080 8634
rect 39028 8570 39080 8576
rect 39856 8628 39908 8634
rect 39856 8570 39908 8576
rect 39868 7954 39896 8570
rect 41248 8090 41276 8842
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 65654 8188 65962 8197
rect 65654 8186 65660 8188
rect 65716 8186 65740 8188
rect 65796 8186 65820 8188
rect 65876 8186 65900 8188
rect 65956 8186 65962 8188
rect 65716 8134 65718 8186
rect 65898 8134 65900 8186
rect 65654 8132 65660 8134
rect 65716 8132 65740 8134
rect 65796 8132 65820 8134
rect 65876 8132 65900 8134
rect 65956 8132 65962 8134
rect 65654 8123 65962 8132
rect 41236 8084 41288 8090
rect 41236 8026 41288 8032
rect 38844 7948 38896 7954
rect 38844 7890 38896 7896
rect 39856 7948 39908 7954
rect 39856 7890 39908 7896
rect 38752 7540 38804 7546
rect 38752 7482 38804 7488
rect 39868 6866 39896 7890
rect 68100 7880 68152 7886
rect 68100 7822 68152 7828
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 68112 7585 68140 7822
rect 68098 7576 68154 7585
rect 68098 7511 68154 7520
rect 39948 7200 40000 7206
rect 39948 7142 40000 7148
rect 39856 6860 39908 6866
rect 39856 6802 39908 6808
rect 39960 6798 39988 7142
rect 65654 7100 65962 7109
rect 65654 7098 65660 7100
rect 65716 7098 65740 7100
rect 65796 7098 65820 7100
rect 65876 7098 65900 7100
rect 65956 7098 65962 7100
rect 65716 7046 65718 7098
rect 65898 7046 65900 7098
rect 65654 7044 65660 7046
rect 65716 7044 65740 7046
rect 65796 7044 65820 7046
rect 65876 7044 65900 7046
rect 65956 7044 65962 7046
rect 65654 7035 65962 7044
rect 38568 6792 38620 6798
rect 38568 6734 38620 6740
rect 39948 6792 40000 6798
rect 39948 6734 40000 6740
rect 38580 6458 38608 6734
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 38568 6452 38620 6458
rect 38568 6394 38620 6400
rect 38660 6384 38712 6390
rect 38660 6326 38712 6332
rect 38476 6316 38528 6322
rect 38476 6258 38528 6264
rect 38488 5914 38516 6258
rect 38476 5908 38528 5914
rect 38476 5850 38528 5856
rect 38292 5772 38344 5778
rect 38292 5714 38344 5720
rect 38108 5636 38160 5642
rect 38108 5578 38160 5584
rect 37740 5568 37792 5574
rect 37740 5510 37792 5516
rect 37464 5296 37516 5302
rect 37464 5238 37516 5244
rect 36268 5228 36320 5234
rect 36268 5170 36320 5176
rect 36452 5228 36504 5234
rect 36452 5170 36504 5176
rect 37372 5228 37424 5234
rect 37372 5170 37424 5176
rect 36280 4826 36308 5170
rect 37476 4826 37504 5238
rect 36268 4820 36320 4826
rect 36268 4762 36320 4768
rect 37464 4820 37516 4826
rect 37464 4762 37516 4768
rect 37752 4622 37780 5510
rect 38672 5370 38700 6326
rect 67638 6216 67694 6225
rect 67638 6151 67640 6160
rect 67692 6151 67694 6160
rect 67640 6122 67692 6128
rect 38752 6112 38804 6118
rect 38752 6054 38804 6060
rect 38660 5364 38712 5370
rect 38660 5306 38712 5312
rect 38764 5302 38792 6054
rect 65654 6012 65962 6021
rect 65654 6010 65660 6012
rect 65716 6010 65740 6012
rect 65796 6010 65820 6012
rect 65876 6010 65900 6012
rect 65956 6010 65962 6012
rect 65716 5958 65718 6010
rect 65898 5958 65900 6010
rect 65654 5956 65660 5958
rect 65716 5956 65740 5958
rect 65796 5956 65820 5958
rect 65876 5956 65900 5958
rect 65956 5956 65962 5958
rect 65654 5947 65962 5956
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 38752 5296 38804 5302
rect 38752 5238 38804 5244
rect 38752 5160 38804 5166
rect 38752 5102 38804 5108
rect 58808 5160 58860 5166
rect 58808 5102 58860 5108
rect 38764 4690 38792 5102
rect 58716 5024 58768 5030
rect 58716 4966 58768 4972
rect 57244 4752 57296 4758
rect 57244 4694 57296 4700
rect 58256 4752 58308 4758
rect 58256 4694 58308 4700
rect 38752 4684 38804 4690
rect 38752 4626 38804 4632
rect 36084 4616 36136 4622
rect 36084 4558 36136 4564
rect 37740 4616 37792 4622
rect 37740 4558 37792 4564
rect 36096 4282 36124 4558
rect 36084 4276 36136 4282
rect 36084 4218 36136 4224
rect 38764 4214 38792 4626
rect 57152 4616 57204 4622
rect 57152 4558 57204 4564
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 35900 4208 35952 4214
rect 35900 4150 35952 4156
rect 38752 4208 38804 4214
rect 38752 4150 38804 4156
rect 33140 4140 33192 4146
rect 33140 4082 33192 4088
rect 33784 4140 33836 4146
rect 33784 4082 33836 4088
rect 35624 4140 35676 4146
rect 35624 4082 35676 4088
rect 33152 3602 33180 4082
rect 56140 3936 56192 3942
rect 56140 3878 56192 3884
rect 56324 3936 56376 3942
rect 56324 3878 56376 3884
rect 56968 3936 57020 3942
rect 56968 3878 57020 3884
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 41144 3664 41196 3670
rect 41144 3606 41196 3612
rect 33140 3596 33192 3602
rect 33140 3538 33192 3544
rect 32864 3528 32916 3534
rect 32864 3470 32916 3476
rect 39212 3528 39264 3534
rect 39212 3470 39264 3476
rect 40040 3528 40092 3534
rect 40040 3470 40092 3476
rect 40868 3528 40920 3534
rect 40868 3470 40920 3476
rect 37280 2984 37332 2990
rect 37280 2926 37332 2932
rect 33140 2848 33192 2854
rect 33140 2790 33192 2796
rect 33692 2848 33744 2854
rect 33692 2790 33744 2796
rect 34244 2848 34296 2854
rect 34244 2790 34296 2796
rect 34520 2848 34572 2854
rect 34520 2790 34572 2796
rect 35348 2848 35400 2854
rect 35348 2790 35400 2796
rect 36176 2848 36228 2854
rect 36176 2790 36228 2796
rect 36728 2848 36780 2854
rect 36728 2790 36780 2796
rect 32864 2576 32916 2582
rect 32864 2518 32916 2524
rect 32876 800 32904 2518
rect 33152 800 33180 2790
rect 33416 2440 33468 2446
rect 33416 2382 33468 2388
rect 33428 800 33456 2382
rect 33704 800 33732 2790
rect 33968 2440 34020 2446
rect 33968 2382 34020 2388
rect 33980 800 34008 2382
rect 34256 800 34284 2790
rect 34532 800 34560 2790
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34796 2440 34848 2446
rect 34796 2382 34848 2388
rect 35072 2440 35124 2446
rect 35072 2382 35124 2388
rect 34808 800 34836 2382
rect 35084 800 35112 2382
rect 35360 800 35388 2790
rect 35624 2440 35676 2446
rect 35624 2382 35676 2388
rect 35900 2440 35952 2446
rect 35900 2382 35952 2388
rect 35636 800 35664 2382
rect 35912 800 35940 2382
rect 36188 800 36216 2790
rect 36452 2440 36504 2446
rect 36452 2382 36504 2388
rect 36464 800 36492 2382
rect 36740 800 36768 2790
rect 37004 2508 37056 2514
rect 37004 2450 37056 2456
rect 37016 800 37044 2450
rect 37292 800 37320 2926
rect 38384 2916 38436 2922
rect 38384 2858 38436 2864
rect 37832 2848 37884 2854
rect 37832 2790 37884 2796
rect 37556 2440 37608 2446
rect 37556 2382 37608 2388
rect 37568 800 37596 2382
rect 37844 800 37872 2790
rect 38108 2508 38160 2514
rect 38108 2450 38160 2456
rect 38120 800 38148 2450
rect 38396 800 38424 2858
rect 38936 2848 38988 2854
rect 38936 2790 38988 2796
rect 38660 2440 38712 2446
rect 38660 2382 38712 2388
rect 38672 800 38700 2382
rect 38948 800 38976 2790
rect 39224 800 39252 3470
rect 39764 2916 39816 2922
rect 39764 2858 39816 2864
rect 39488 2372 39540 2378
rect 39488 2314 39540 2320
rect 39500 800 39528 2314
rect 39776 800 39804 2858
rect 40052 800 40080 3470
rect 40316 2848 40368 2854
rect 40316 2790 40368 2796
rect 40328 800 40356 2790
rect 40592 2576 40644 2582
rect 40592 2518 40644 2524
rect 40604 800 40632 2518
rect 40880 800 40908 3470
rect 41156 800 41184 3606
rect 55772 3596 55824 3602
rect 55772 3538 55824 3544
rect 42524 3528 42576 3534
rect 42524 3470 42576 3476
rect 43076 3528 43128 3534
rect 43076 3470 43128 3476
rect 45008 3528 45060 3534
rect 45008 3470 45060 3476
rect 45284 3528 45336 3534
rect 45284 3470 45336 3476
rect 46112 3528 46164 3534
rect 46112 3470 46164 3476
rect 46940 3528 46992 3534
rect 46940 3470 46992 3476
rect 47768 3528 47820 3534
rect 47768 3470 47820 3476
rect 48872 3528 48924 3534
rect 48872 3470 48924 3476
rect 50160 3528 50212 3534
rect 50160 3470 50212 3476
rect 50804 3528 50856 3534
rect 50804 3470 50856 3476
rect 51356 3528 51408 3534
rect 51356 3470 51408 3476
rect 52736 3528 52788 3534
rect 52736 3470 52788 3476
rect 53012 3528 53064 3534
rect 53012 3470 53064 3476
rect 54668 3528 54720 3534
rect 54668 3470 54720 3476
rect 55496 3528 55548 3534
rect 55496 3470 55548 3476
rect 42248 2916 42300 2922
rect 42248 2858 42300 2864
rect 41696 2848 41748 2854
rect 41696 2790 41748 2796
rect 41420 2508 41472 2514
rect 41420 2450 41472 2456
rect 41432 800 41460 2450
rect 41708 800 41736 2790
rect 41972 2440 42024 2446
rect 41972 2382 42024 2388
rect 41984 800 42012 2382
rect 42260 800 42288 2858
rect 42536 800 42564 3470
rect 42800 2848 42852 2854
rect 42800 2790 42852 2796
rect 42812 800 42840 2790
rect 43088 800 43116 3470
rect 44732 2984 44784 2990
rect 44732 2926 44784 2932
rect 43628 2916 43680 2922
rect 43628 2858 43680 2864
rect 43352 2508 43404 2514
rect 43352 2450 43404 2456
rect 43364 800 43392 2450
rect 43640 800 43668 2858
rect 44180 2848 44232 2854
rect 44180 2790 44232 2796
rect 43904 2372 43956 2378
rect 43904 2314 43956 2320
rect 43916 800 43944 2314
rect 44192 800 44220 2790
rect 44456 2576 44508 2582
rect 44456 2518 44508 2524
rect 44468 800 44496 2518
rect 44744 800 44772 2926
rect 45020 800 45048 3470
rect 45296 800 45324 3470
rect 45560 2848 45612 2854
rect 45560 2790 45612 2796
rect 45572 800 45600 2790
rect 45836 2440 45888 2446
rect 45836 2382 45888 2388
rect 45848 800 45876 2382
rect 46124 800 46152 3470
rect 46664 2848 46716 2854
rect 46664 2790 46716 2796
rect 46388 2508 46440 2514
rect 46388 2450 46440 2456
rect 46400 800 46428 2450
rect 46676 800 46704 2790
rect 46952 800 46980 3470
rect 47492 2916 47544 2922
rect 47492 2858 47544 2864
rect 47216 2372 47268 2378
rect 47216 2314 47268 2320
rect 47228 800 47256 2314
rect 47504 800 47532 2858
rect 47780 800 47808 3470
rect 48596 2984 48648 2990
rect 48596 2926 48648 2932
rect 48044 2848 48096 2854
rect 48044 2790 48096 2796
rect 48056 800 48084 2790
rect 48320 2576 48372 2582
rect 48320 2518 48372 2524
rect 48332 800 48360 2518
rect 48608 800 48636 2926
rect 48884 800 48912 3470
rect 49424 2916 49476 2922
rect 49424 2858 49476 2864
rect 49148 2508 49200 2514
rect 49148 2450 49200 2456
rect 49160 800 49188 2450
rect 49436 800 49464 2858
rect 49976 2848 50028 2854
rect 49976 2790 50028 2796
rect 49700 2440 49752 2446
rect 49700 2382 49752 2388
rect 49712 800 49740 2382
rect 49988 800 50016 2790
rect 50172 1850 50200 3470
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 50620 2916 50672 2922
rect 50620 2858 50672 2864
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 50172 1822 50292 1850
rect 50264 800 50292 1822
rect 50632 1442 50660 2858
rect 50540 1414 50660 1442
rect 50540 800 50568 1414
rect 50816 800 50844 3470
rect 51080 2508 51132 2514
rect 51080 2450 51132 2456
rect 51092 800 51120 2450
rect 51368 800 51396 3470
rect 52460 2984 52512 2990
rect 52460 2926 52512 2932
rect 51908 2848 51960 2854
rect 51908 2790 51960 2796
rect 51632 2440 51684 2446
rect 51632 2382 51684 2388
rect 51644 800 51672 2382
rect 51920 800 51948 2790
rect 52184 2576 52236 2582
rect 52184 2518 52236 2524
rect 52196 800 52224 2518
rect 52472 800 52500 2926
rect 52748 800 52776 3470
rect 53024 800 53052 3470
rect 53564 2984 53616 2990
rect 53564 2926 53616 2932
rect 53288 2916 53340 2922
rect 53288 2858 53340 2864
rect 53300 800 53328 2858
rect 53576 800 53604 2926
rect 54392 2916 54444 2922
rect 54392 2858 54444 2864
rect 53840 2848 53892 2854
rect 53840 2790 53892 2796
rect 53852 800 53880 2790
rect 54116 2372 54168 2378
rect 54116 2314 54168 2320
rect 54128 800 54156 2314
rect 54404 800 54432 2858
rect 54680 800 54708 3470
rect 55220 2984 55272 2990
rect 55220 2926 55272 2932
rect 55232 2650 55260 2926
rect 55404 2848 55456 2854
rect 55404 2790 55456 2796
rect 55220 2644 55272 2650
rect 55220 2586 55272 2592
rect 54944 2508 54996 2514
rect 54944 2450 54996 2456
rect 54956 800 54984 2450
rect 55416 1442 55444 2790
rect 55232 1414 55444 1442
rect 55232 800 55260 1414
rect 55508 800 55536 3470
rect 55680 2916 55732 2922
rect 55680 2858 55732 2864
rect 55692 800 55720 2858
rect 55784 800 55812 3538
rect 55956 3188 56008 3194
rect 55956 3130 56008 3136
rect 55864 2576 55916 2582
rect 55864 2518 55916 2524
rect 55876 800 55904 2518
rect 55968 800 55996 3130
rect 56048 2848 56100 2854
rect 56048 2790 56100 2796
rect 56060 800 56088 2790
rect 56152 800 56180 3878
rect 56232 3528 56284 3534
rect 56232 3470 56284 3476
rect 56244 800 56272 3470
rect 56336 800 56364 3878
rect 56508 3664 56560 3670
rect 56508 3606 56560 3612
rect 56416 2440 56468 2446
rect 56416 2382 56468 2388
rect 56428 800 56456 2382
rect 56520 800 56548 3606
rect 56784 3596 56836 3602
rect 56784 3538 56836 3544
rect 56692 2984 56744 2990
rect 56692 2926 56744 2932
rect 56704 1442 56732 2926
rect 56612 1414 56732 1442
rect 56612 800 56640 1414
rect 56796 1306 56824 3538
rect 56876 2304 56928 2310
rect 56876 2246 56928 2252
rect 56704 1278 56824 1306
rect 56704 800 56732 1278
rect 56784 1216 56836 1222
rect 56784 1158 56836 1164
rect 56796 800 56824 1158
rect 56888 800 56916 2246
rect 56980 800 57008 3878
rect 57060 2916 57112 2922
rect 57060 2858 57112 2864
rect 57072 1222 57100 2858
rect 57060 1216 57112 1222
rect 57060 1158 57112 1164
rect 57060 1080 57112 1086
rect 57060 1022 57112 1028
rect 57072 800 57100 1022
rect 57164 800 57192 4558
rect 57256 800 57284 4694
rect 57612 4616 57664 4622
rect 57612 4558 57664 4564
rect 57520 4004 57572 4010
rect 57520 3946 57572 3952
rect 57336 3528 57388 3534
rect 57336 3470 57388 3476
rect 57348 800 57376 3470
rect 57428 2644 57480 2650
rect 57428 2586 57480 2592
rect 57440 800 57468 2586
rect 57532 800 57560 3946
rect 57624 800 57652 4558
rect 57980 4140 58032 4146
rect 57980 4082 58032 4088
rect 57796 3732 57848 3738
rect 57796 3674 57848 3680
rect 57704 3120 57756 3126
rect 57704 3062 57756 3068
rect 57716 800 57744 3062
rect 57808 800 57836 3674
rect 57886 3224 57942 3233
rect 57886 3159 57942 3168
rect 57900 800 57928 3159
rect 57992 800 58020 4082
rect 58072 3936 58124 3942
rect 58072 3878 58124 3884
rect 58084 3738 58112 3878
rect 58072 3732 58124 3738
rect 58072 3674 58124 3680
rect 58072 3188 58124 3194
rect 58072 3130 58124 3136
rect 58084 2582 58112 3130
rect 58164 3052 58216 3058
rect 58164 2994 58216 3000
rect 58072 2576 58124 2582
rect 58072 2518 58124 2524
rect 58072 2100 58124 2106
rect 58072 2042 58124 2048
rect 58084 800 58112 2042
rect 58176 800 58204 2994
rect 58268 800 58296 4694
rect 58624 4004 58676 4010
rect 58624 3946 58676 3952
rect 58348 3664 58400 3670
rect 58348 3606 58400 3612
rect 58360 800 58388 3606
rect 58440 2984 58492 2990
rect 58440 2926 58492 2932
rect 58452 800 58480 2926
rect 58532 1964 58584 1970
rect 58532 1906 58584 1912
rect 58544 800 58572 1906
rect 58636 800 58664 3946
rect 58728 800 58756 4966
rect 58820 800 58848 5102
rect 59268 5092 59320 5098
rect 59268 5034 59320 5040
rect 58900 4684 58952 4690
rect 58900 4626 58952 4632
rect 58912 800 58940 4626
rect 59176 4072 59228 4078
rect 59176 4014 59228 4020
rect 58992 3596 59044 3602
rect 58992 3538 59044 3544
rect 59004 800 59032 3538
rect 59084 2032 59136 2038
rect 59084 1974 59136 1980
rect 59096 800 59124 1974
rect 59188 800 59216 4014
rect 59280 800 59308 5034
rect 67640 5024 67692 5030
rect 67640 4966 67692 4972
rect 65654 4924 65962 4933
rect 65654 4922 65660 4924
rect 65716 4922 65740 4924
rect 65796 4922 65820 4924
rect 65876 4922 65900 4924
rect 65956 4922 65962 4924
rect 65716 4870 65718 4922
rect 65898 4870 65900 4922
rect 65654 4868 65660 4870
rect 65716 4868 65740 4870
rect 65796 4868 65820 4870
rect 65876 4868 65900 4870
rect 65956 4868 65962 4870
rect 65654 4859 65962 4868
rect 67652 4865 67680 4966
rect 67638 4856 67694 4865
rect 67638 4791 67694 4800
rect 65654 3836 65962 3845
rect 65654 3834 65660 3836
rect 65716 3834 65740 3836
rect 65796 3834 65820 3836
rect 65876 3834 65900 3836
rect 65956 3834 65962 3836
rect 65716 3782 65718 3834
rect 65898 3782 65900 3834
rect 65654 3780 65660 3782
rect 65716 3780 65740 3782
rect 65796 3780 65820 3782
rect 65876 3780 65900 3782
rect 65956 3780 65962 3782
rect 65654 3771 65962 3780
rect 60464 3528 60516 3534
rect 68100 3528 68152 3534
rect 60464 3470 60516 3476
rect 68098 3496 68100 3505
rect 68152 3496 68154 3505
rect 60476 3233 60504 3470
rect 68098 3431 68154 3440
rect 60462 3224 60518 3233
rect 60462 3159 60518 3168
rect 60464 3120 60516 3126
rect 60464 3062 60516 3068
rect 59360 2916 59412 2922
rect 59360 2858 59412 2864
rect 59372 800 59400 2858
rect 60476 2854 60504 3062
rect 59452 2848 59504 2854
rect 59452 2790 59504 2796
rect 60464 2848 60516 2854
rect 60464 2790 60516 2796
rect 59464 1086 59492 2790
rect 65654 2748 65962 2757
rect 65654 2746 65660 2748
rect 65716 2746 65740 2748
rect 65796 2746 65820 2748
rect 65876 2746 65900 2748
rect 65956 2746 65962 2748
rect 65716 2694 65718 2746
rect 65898 2694 65900 2746
rect 65654 2692 65660 2694
rect 65716 2692 65740 2694
rect 65796 2692 65820 2694
rect 65876 2692 65900 2694
rect 65956 2692 65962 2694
rect 65654 2683 65962 2692
rect 63684 2508 63736 2514
rect 63684 2450 63736 2456
rect 61752 2440 61804 2446
rect 61752 2382 61804 2388
rect 63040 2440 63092 2446
rect 63040 2382 63092 2388
rect 61764 2106 61792 2382
rect 61752 2100 61804 2106
rect 61752 2042 61804 2048
rect 63052 1970 63080 2382
rect 63696 2038 63724 2450
rect 66996 2440 67048 2446
rect 66996 2382 67048 2388
rect 67548 2440 67600 2446
rect 67548 2382 67600 2388
rect 67008 2145 67036 2382
rect 66994 2136 67050 2145
rect 66994 2071 67050 2080
rect 63684 2032 63736 2038
rect 63684 1974 63736 1980
rect 63040 1964 63092 1970
rect 63040 1906 63092 1912
rect 59452 1080 59504 1086
rect 59452 1022 59504 1028
rect 10244 734 10548 762
rect 2504 196 2556 202
rect 2504 138 2556 144
rect 9680 196 9732 202
rect 9680 138 9732 144
rect 10598 0 10654 800
rect 10690 0 10746 800
rect 10782 0 10838 800
rect 10874 0 10930 800
rect 10966 0 11022 800
rect 11058 0 11114 800
rect 11150 0 11206 800
rect 11242 0 11298 800
rect 11334 0 11390 800
rect 11426 0 11482 800
rect 11518 0 11574 800
rect 11610 0 11666 800
rect 11702 0 11758 800
rect 11794 0 11850 800
rect 11886 0 11942 800
rect 11978 0 12034 800
rect 12070 0 12126 800
rect 12162 0 12218 800
rect 12254 0 12310 800
rect 12346 0 12402 800
rect 12438 0 12494 800
rect 12530 0 12586 800
rect 12622 0 12678 800
rect 12714 0 12770 800
rect 12806 0 12862 800
rect 12898 0 12954 800
rect 12990 0 13046 800
rect 13082 0 13138 800
rect 13174 0 13230 800
rect 13266 0 13322 800
rect 13358 0 13414 800
rect 13450 0 13506 800
rect 13542 0 13598 800
rect 13634 0 13690 800
rect 13726 0 13782 800
rect 13818 0 13874 800
rect 13910 0 13966 800
rect 14002 0 14058 800
rect 14094 0 14150 800
rect 14186 0 14242 800
rect 14278 0 14334 800
rect 14370 0 14426 800
rect 14462 0 14518 800
rect 14554 0 14610 800
rect 14646 0 14702 800
rect 14738 0 14794 800
rect 14830 0 14886 800
rect 14922 0 14978 800
rect 15014 0 15070 800
rect 15106 0 15162 800
rect 15198 0 15254 800
rect 15290 0 15346 800
rect 15382 0 15438 800
rect 15474 0 15530 800
rect 15566 0 15622 800
rect 15658 0 15714 800
rect 15750 0 15806 800
rect 15842 0 15898 800
rect 15934 0 15990 800
rect 16026 0 16082 800
rect 16118 0 16174 800
rect 16210 0 16266 800
rect 16302 0 16358 800
rect 16394 0 16450 800
rect 16486 0 16542 800
rect 16578 0 16634 800
rect 16670 0 16726 800
rect 16762 0 16818 800
rect 16854 0 16910 800
rect 16946 0 17002 800
rect 17038 0 17094 800
rect 17130 0 17186 800
rect 17222 0 17278 800
rect 17314 0 17370 800
rect 17406 0 17462 800
rect 17498 0 17554 800
rect 17590 0 17646 800
rect 17682 0 17738 800
rect 17774 0 17830 800
rect 17866 0 17922 800
rect 17958 0 18014 800
rect 18050 0 18106 800
rect 18142 0 18198 800
rect 18234 0 18290 800
rect 18326 0 18382 800
rect 18418 0 18474 800
rect 18510 0 18566 800
rect 18602 0 18658 800
rect 18694 0 18750 800
rect 18786 0 18842 800
rect 18878 0 18934 800
rect 18970 0 19026 800
rect 19062 0 19118 800
rect 19154 0 19210 800
rect 19246 0 19302 800
rect 19338 0 19394 800
rect 19430 0 19486 800
rect 19522 0 19578 800
rect 19614 0 19670 800
rect 19706 0 19762 800
rect 19798 0 19854 800
rect 19890 0 19946 800
rect 19982 0 20038 800
rect 20074 0 20130 800
rect 20166 0 20222 800
rect 20258 0 20314 800
rect 20350 0 20406 800
rect 20442 0 20498 800
rect 20534 0 20590 800
rect 20626 0 20682 800
rect 20718 0 20774 800
rect 20810 0 20866 800
rect 20902 0 20958 800
rect 20994 0 21050 800
rect 21086 0 21142 800
rect 21178 0 21234 800
rect 21270 0 21326 800
rect 21362 0 21418 800
rect 21454 0 21510 800
rect 21546 0 21602 800
rect 21638 0 21694 800
rect 21730 0 21786 800
rect 21822 0 21878 800
rect 21914 0 21970 800
rect 22006 0 22062 800
rect 22098 0 22154 800
rect 22190 0 22246 800
rect 22282 0 22338 800
rect 22374 0 22430 800
rect 22466 0 22522 800
rect 22558 0 22614 800
rect 22650 0 22706 800
rect 22742 0 22798 800
rect 22834 0 22890 800
rect 22926 0 22982 800
rect 23018 0 23074 800
rect 23110 0 23166 800
rect 23202 0 23258 800
rect 23294 0 23350 800
rect 23386 0 23442 800
rect 23478 0 23534 800
rect 23570 0 23626 800
rect 23662 0 23718 800
rect 23754 0 23810 800
rect 23846 0 23902 800
rect 23938 0 23994 800
rect 24030 0 24086 800
rect 24122 0 24178 800
rect 24214 0 24270 800
rect 24306 0 24362 800
rect 24398 0 24454 800
rect 24490 0 24546 800
rect 24582 0 24638 800
rect 24674 0 24730 800
rect 24766 0 24822 800
rect 24858 0 24914 800
rect 24950 0 25006 800
rect 25042 0 25098 800
rect 25134 0 25190 800
rect 25226 0 25282 800
rect 25318 0 25374 800
rect 25410 0 25466 800
rect 25502 0 25558 800
rect 25594 0 25650 800
rect 25686 0 25742 800
rect 25778 0 25834 800
rect 25870 0 25926 800
rect 25962 0 26018 800
rect 26054 0 26110 800
rect 26146 0 26202 800
rect 26238 0 26294 800
rect 26330 0 26386 800
rect 26422 0 26478 800
rect 26514 0 26570 800
rect 26606 0 26662 800
rect 26698 0 26754 800
rect 26790 0 26846 800
rect 26882 0 26938 800
rect 26974 0 27030 800
rect 27066 0 27122 800
rect 27158 0 27214 800
rect 27250 0 27306 800
rect 27342 0 27398 800
rect 27434 0 27490 800
rect 27526 0 27582 800
rect 27618 0 27674 800
rect 27710 0 27766 800
rect 27802 0 27858 800
rect 27894 0 27950 800
rect 27986 0 28042 800
rect 28078 0 28134 800
rect 28170 0 28226 800
rect 28262 0 28318 800
rect 28354 0 28410 800
rect 28446 0 28502 800
rect 28538 0 28594 800
rect 28630 0 28686 800
rect 28722 0 28778 800
rect 28814 0 28870 800
rect 28906 0 28962 800
rect 28998 0 29054 800
rect 29090 0 29146 800
rect 29182 0 29238 800
rect 29274 0 29330 800
rect 29366 0 29422 800
rect 29458 0 29514 800
rect 29550 0 29606 800
rect 29642 0 29698 800
rect 29734 0 29790 800
rect 29826 0 29882 800
rect 29918 0 29974 800
rect 30010 0 30066 800
rect 30102 0 30158 800
rect 30194 0 30250 800
rect 30286 0 30342 800
rect 30378 0 30434 800
rect 30470 0 30526 800
rect 30562 0 30618 800
rect 30654 0 30710 800
rect 30746 0 30802 800
rect 30838 0 30894 800
rect 30930 0 30986 800
rect 31022 0 31078 800
rect 31114 0 31170 800
rect 31206 0 31262 800
rect 31298 0 31354 800
rect 31390 0 31446 800
rect 31482 0 31538 800
rect 31574 0 31630 800
rect 31666 0 31722 800
rect 31758 0 31814 800
rect 31850 0 31906 800
rect 31942 0 31998 800
rect 32034 0 32090 800
rect 32126 0 32182 800
rect 32218 0 32274 800
rect 32310 0 32366 800
rect 32402 0 32458 800
rect 32494 0 32550 800
rect 32586 0 32642 800
rect 32678 0 32734 800
rect 32770 0 32826 800
rect 32862 0 32918 800
rect 32954 0 33010 800
rect 33046 0 33102 800
rect 33138 0 33194 800
rect 33230 0 33286 800
rect 33322 0 33378 800
rect 33414 0 33470 800
rect 33506 0 33562 800
rect 33598 0 33654 800
rect 33690 0 33746 800
rect 33782 0 33838 800
rect 33874 0 33930 800
rect 33966 0 34022 800
rect 34058 0 34114 800
rect 34150 0 34206 800
rect 34242 0 34298 800
rect 34334 0 34390 800
rect 34426 0 34482 800
rect 34518 0 34574 800
rect 34610 0 34666 800
rect 34702 0 34758 800
rect 34794 0 34850 800
rect 34886 0 34942 800
rect 34978 0 35034 800
rect 35070 0 35126 800
rect 35162 0 35218 800
rect 35254 0 35310 800
rect 35346 0 35402 800
rect 35438 0 35494 800
rect 35530 0 35586 800
rect 35622 0 35678 800
rect 35714 0 35770 800
rect 35806 0 35862 800
rect 35898 0 35954 800
rect 35990 0 36046 800
rect 36082 0 36138 800
rect 36174 0 36230 800
rect 36266 0 36322 800
rect 36358 0 36414 800
rect 36450 0 36506 800
rect 36542 0 36598 800
rect 36634 0 36690 800
rect 36726 0 36782 800
rect 36818 0 36874 800
rect 36910 0 36966 800
rect 37002 0 37058 800
rect 37094 0 37150 800
rect 37186 0 37242 800
rect 37278 0 37334 800
rect 37370 0 37426 800
rect 37462 0 37518 800
rect 37554 0 37610 800
rect 37646 0 37702 800
rect 37738 0 37794 800
rect 37830 0 37886 800
rect 37922 0 37978 800
rect 38014 0 38070 800
rect 38106 0 38162 800
rect 38198 0 38254 800
rect 38290 0 38346 800
rect 38382 0 38438 800
rect 38474 0 38530 800
rect 38566 0 38622 800
rect 38658 0 38714 800
rect 38750 0 38806 800
rect 38842 0 38898 800
rect 38934 0 38990 800
rect 39026 0 39082 800
rect 39118 0 39174 800
rect 39210 0 39266 800
rect 39302 0 39358 800
rect 39394 0 39450 800
rect 39486 0 39542 800
rect 39578 0 39634 800
rect 39670 0 39726 800
rect 39762 0 39818 800
rect 39854 0 39910 800
rect 39946 0 40002 800
rect 40038 0 40094 800
rect 40130 0 40186 800
rect 40222 0 40278 800
rect 40314 0 40370 800
rect 40406 0 40462 800
rect 40498 0 40554 800
rect 40590 0 40646 800
rect 40682 0 40738 800
rect 40774 0 40830 800
rect 40866 0 40922 800
rect 40958 0 41014 800
rect 41050 0 41106 800
rect 41142 0 41198 800
rect 41234 0 41290 800
rect 41326 0 41382 800
rect 41418 0 41474 800
rect 41510 0 41566 800
rect 41602 0 41658 800
rect 41694 0 41750 800
rect 41786 0 41842 800
rect 41878 0 41934 800
rect 41970 0 42026 800
rect 42062 0 42118 800
rect 42154 0 42210 800
rect 42246 0 42302 800
rect 42338 0 42394 800
rect 42430 0 42486 800
rect 42522 0 42578 800
rect 42614 0 42670 800
rect 42706 0 42762 800
rect 42798 0 42854 800
rect 42890 0 42946 800
rect 42982 0 43038 800
rect 43074 0 43130 800
rect 43166 0 43222 800
rect 43258 0 43314 800
rect 43350 0 43406 800
rect 43442 0 43498 800
rect 43534 0 43590 800
rect 43626 0 43682 800
rect 43718 0 43774 800
rect 43810 0 43866 800
rect 43902 0 43958 800
rect 43994 0 44050 800
rect 44086 0 44142 800
rect 44178 0 44234 800
rect 44270 0 44326 800
rect 44362 0 44418 800
rect 44454 0 44510 800
rect 44546 0 44602 800
rect 44638 0 44694 800
rect 44730 0 44786 800
rect 44822 0 44878 800
rect 44914 0 44970 800
rect 45006 0 45062 800
rect 45098 0 45154 800
rect 45190 0 45246 800
rect 45282 0 45338 800
rect 45374 0 45430 800
rect 45466 0 45522 800
rect 45558 0 45614 800
rect 45650 0 45706 800
rect 45742 0 45798 800
rect 45834 0 45890 800
rect 45926 0 45982 800
rect 46018 0 46074 800
rect 46110 0 46166 800
rect 46202 0 46258 800
rect 46294 0 46350 800
rect 46386 0 46442 800
rect 46478 0 46534 800
rect 46570 0 46626 800
rect 46662 0 46718 800
rect 46754 0 46810 800
rect 46846 0 46902 800
rect 46938 0 46994 800
rect 47030 0 47086 800
rect 47122 0 47178 800
rect 47214 0 47270 800
rect 47306 0 47362 800
rect 47398 0 47454 800
rect 47490 0 47546 800
rect 47582 0 47638 800
rect 47674 0 47730 800
rect 47766 0 47822 800
rect 47858 0 47914 800
rect 47950 0 48006 800
rect 48042 0 48098 800
rect 48134 0 48190 800
rect 48226 0 48282 800
rect 48318 0 48374 800
rect 48410 0 48466 800
rect 48502 0 48558 800
rect 48594 0 48650 800
rect 48686 0 48742 800
rect 48778 0 48834 800
rect 48870 0 48926 800
rect 48962 0 49018 800
rect 49054 0 49110 800
rect 49146 0 49202 800
rect 49238 0 49294 800
rect 49330 0 49386 800
rect 49422 0 49478 800
rect 49514 0 49570 800
rect 49606 0 49662 800
rect 49698 0 49754 800
rect 49790 0 49846 800
rect 49882 0 49938 800
rect 49974 0 50030 800
rect 50066 0 50122 800
rect 50158 0 50214 800
rect 50250 0 50306 800
rect 50342 0 50398 800
rect 50434 0 50490 800
rect 50526 0 50582 800
rect 50618 0 50674 800
rect 50710 0 50766 800
rect 50802 0 50858 800
rect 50894 0 50950 800
rect 50986 0 51042 800
rect 51078 0 51134 800
rect 51170 0 51226 800
rect 51262 0 51318 800
rect 51354 0 51410 800
rect 51446 0 51502 800
rect 51538 0 51594 800
rect 51630 0 51686 800
rect 51722 0 51778 800
rect 51814 0 51870 800
rect 51906 0 51962 800
rect 51998 0 52054 800
rect 52090 0 52146 800
rect 52182 0 52238 800
rect 52274 0 52330 800
rect 52366 0 52422 800
rect 52458 0 52514 800
rect 52550 0 52606 800
rect 52642 0 52698 800
rect 52734 0 52790 800
rect 52826 0 52882 800
rect 52918 0 52974 800
rect 53010 0 53066 800
rect 53102 0 53158 800
rect 53194 0 53250 800
rect 53286 0 53342 800
rect 53378 0 53434 800
rect 53470 0 53526 800
rect 53562 0 53618 800
rect 53654 0 53710 800
rect 53746 0 53802 800
rect 53838 0 53894 800
rect 53930 0 53986 800
rect 54022 0 54078 800
rect 54114 0 54170 800
rect 54206 0 54262 800
rect 54298 0 54354 800
rect 54390 0 54446 800
rect 54482 0 54538 800
rect 54574 0 54630 800
rect 54666 0 54722 800
rect 54758 0 54814 800
rect 54850 0 54906 800
rect 54942 0 54998 800
rect 55034 0 55090 800
rect 55126 0 55182 800
rect 55218 0 55274 800
rect 55310 0 55366 800
rect 55402 0 55458 800
rect 55494 0 55550 800
rect 55586 0 55642 800
rect 55678 0 55734 800
rect 55770 0 55826 800
rect 55862 0 55918 800
rect 55954 0 56010 800
rect 56046 0 56102 800
rect 56138 0 56194 800
rect 56230 0 56286 800
rect 56322 0 56378 800
rect 56414 0 56470 800
rect 56506 0 56562 800
rect 56598 0 56654 800
rect 56690 0 56746 800
rect 56782 0 56838 800
rect 56874 0 56930 800
rect 56966 0 57022 800
rect 57058 0 57114 800
rect 57150 0 57206 800
rect 57242 0 57298 800
rect 57334 0 57390 800
rect 57426 0 57482 800
rect 57518 0 57574 800
rect 57610 0 57666 800
rect 57702 0 57758 800
rect 57794 0 57850 800
rect 57886 0 57942 800
rect 57978 0 58034 800
rect 58070 0 58126 800
rect 58162 0 58218 800
rect 58254 0 58310 800
rect 58346 0 58402 800
rect 58438 0 58494 800
rect 58530 0 58586 800
rect 58622 0 58678 800
rect 58714 0 58770 800
rect 58806 0 58862 800
rect 58898 0 58954 800
rect 58990 0 59046 800
rect 59082 0 59138 800
rect 59174 0 59230 800
rect 59266 0 59322 800
rect 59358 0 59414 800
rect 67560 785 67588 2382
rect 67546 776 67602 785
rect 67546 711 67602 720
<< via2 >>
rect 67546 59200 67602 59256
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 66994 57840 67050 57896
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 65660 57146 65716 57148
rect 65740 57146 65796 57148
rect 65820 57146 65876 57148
rect 65900 57146 65956 57148
rect 65660 57094 65706 57146
rect 65706 57094 65716 57146
rect 65740 57094 65770 57146
rect 65770 57094 65782 57146
rect 65782 57094 65796 57146
rect 65820 57094 65834 57146
rect 65834 57094 65846 57146
rect 65846 57094 65876 57146
rect 65900 57094 65910 57146
rect 65910 57094 65956 57146
rect 65660 57092 65716 57094
rect 65740 57092 65796 57094
rect 65820 57092 65876 57094
rect 65900 57092 65956 57094
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 68098 56480 68154 56536
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 65660 56058 65716 56060
rect 65740 56058 65796 56060
rect 65820 56058 65876 56060
rect 65900 56058 65956 56060
rect 65660 56006 65706 56058
rect 65706 56006 65716 56058
rect 65740 56006 65770 56058
rect 65770 56006 65782 56058
rect 65782 56006 65796 56058
rect 65820 56006 65834 56058
rect 65834 56006 65846 56058
rect 65846 56006 65876 56058
rect 65900 56006 65910 56058
rect 65910 56006 65956 56058
rect 65660 56004 65716 56006
rect 65740 56004 65796 56006
rect 65820 56004 65876 56006
rect 65900 56004 65956 56006
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 67638 55140 67694 55176
rect 67638 55120 67640 55140
rect 67640 55120 67692 55140
rect 67692 55120 67694 55140
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 65660 54970 65716 54972
rect 65740 54970 65796 54972
rect 65820 54970 65876 54972
rect 65900 54970 65956 54972
rect 65660 54918 65706 54970
rect 65706 54918 65716 54970
rect 65740 54918 65770 54970
rect 65770 54918 65782 54970
rect 65782 54918 65796 54970
rect 65820 54918 65834 54970
rect 65834 54918 65846 54970
rect 65846 54918 65876 54970
rect 65900 54918 65910 54970
rect 65910 54918 65956 54970
rect 65660 54916 65716 54918
rect 65740 54916 65796 54918
rect 65820 54916 65876 54918
rect 65900 54916 65956 54918
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 65660 53882 65716 53884
rect 65740 53882 65796 53884
rect 65820 53882 65876 53884
rect 65900 53882 65956 53884
rect 65660 53830 65706 53882
rect 65706 53830 65716 53882
rect 65740 53830 65770 53882
rect 65770 53830 65782 53882
rect 65782 53830 65796 53882
rect 65820 53830 65834 53882
rect 65834 53830 65846 53882
rect 65846 53830 65876 53882
rect 65900 53830 65910 53882
rect 65910 53830 65956 53882
rect 65660 53828 65716 53830
rect 65740 53828 65796 53830
rect 65820 53828 65876 53830
rect 65900 53828 65956 53830
rect 67546 53760 67602 53816
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 65660 52794 65716 52796
rect 65740 52794 65796 52796
rect 65820 52794 65876 52796
rect 65900 52794 65956 52796
rect 65660 52742 65706 52794
rect 65706 52742 65716 52794
rect 65740 52742 65770 52794
rect 65770 52742 65782 52794
rect 65782 52742 65796 52794
rect 65820 52742 65834 52794
rect 65834 52742 65846 52794
rect 65846 52742 65876 52794
rect 65900 52742 65910 52794
rect 65910 52742 65956 52794
rect 65660 52740 65716 52742
rect 65740 52740 65796 52742
rect 65820 52740 65876 52742
rect 65900 52740 65956 52742
rect 68098 52436 68100 52456
rect 68100 52436 68152 52456
rect 68152 52436 68154 52456
rect 68098 52400 68154 52436
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 65660 51706 65716 51708
rect 65740 51706 65796 51708
rect 65820 51706 65876 51708
rect 65900 51706 65956 51708
rect 65660 51654 65706 51706
rect 65706 51654 65716 51706
rect 65740 51654 65770 51706
rect 65770 51654 65782 51706
rect 65782 51654 65796 51706
rect 65820 51654 65834 51706
rect 65834 51654 65846 51706
rect 65846 51654 65876 51706
rect 65900 51654 65910 51706
rect 65910 51654 65956 51706
rect 65660 51652 65716 51654
rect 65740 51652 65796 51654
rect 65820 51652 65876 51654
rect 65900 51652 65956 51654
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 68098 51040 68154 51096
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 65660 50618 65716 50620
rect 65740 50618 65796 50620
rect 65820 50618 65876 50620
rect 65900 50618 65956 50620
rect 65660 50566 65706 50618
rect 65706 50566 65716 50618
rect 65740 50566 65770 50618
rect 65770 50566 65782 50618
rect 65782 50566 65796 50618
rect 65820 50566 65834 50618
rect 65834 50566 65846 50618
rect 65846 50566 65876 50618
rect 65900 50566 65910 50618
rect 65910 50566 65956 50618
rect 65660 50564 65716 50566
rect 65740 50564 65796 50566
rect 65820 50564 65876 50566
rect 65900 50564 65956 50566
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 67638 49716 67640 49736
rect 67640 49716 67692 49736
rect 67692 49716 67694 49736
rect 67638 49680 67694 49716
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 65660 49530 65716 49532
rect 65740 49530 65796 49532
rect 65820 49530 65876 49532
rect 65900 49530 65956 49532
rect 65660 49478 65706 49530
rect 65706 49478 65716 49530
rect 65740 49478 65770 49530
rect 65770 49478 65782 49530
rect 65782 49478 65796 49530
rect 65820 49478 65834 49530
rect 65834 49478 65846 49530
rect 65846 49478 65876 49530
rect 65900 49478 65910 49530
rect 65910 49478 65956 49530
rect 65660 49476 65716 49478
rect 65740 49476 65796 49478
rect 65820 49476 65876 49478
rect 65900 49476 65956 49478
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 65660 48442 65716 48444
rect 65740 48442 65796 48444
rect 65820 48442 65876 48444
rect 65900 48442 65956 48444
rect 65660 48390 65706 48442
rect 65706 48390 65716 48442
rect 65740 48390 65770 48442
rect 65770 48390 65782 48442
rect 65782 48390 65796 48442
rect 65820 48390 65834 48442
rect 65834 48390 65846 48442
rect 65846 48390 65876 48442
rect 65900 48390 65910 48442
rect 65910 48390 65956 48442
rect 65660 48388 65716 48390
rect 65740 48388 65796 48390
rect 65820 48388 65876 48390
rect 65900 48388 65956 48390
rect 67638 48320 67694 48376
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 65660 47354 65716 47356
rect 65740 47354 65796 47356
rect 65820 47354 65876 47356
rect 65900 47354 65956 47356
rect 65660 47302 65706 47354
rect 65706 47302 65716 47354
rect 65740 47302 65770 47354
rect 65770 47302 65782 47354
rect 65782 47302 65796 47354
rect 65820 47302 65834 47354
rect 65834 47302 65846 47354
rect 65846 47302 65876 47354
rect 65900 47302 65910 47354
rect 65910 47302 65956 47354
rect 65660 47300 65716 47302
rect 65740 47300 65796 47302
rect 65820 47300 65876 47302
rect 65900 47300 65956 47302
rect 68098 46996 68100 47016
rect 68100 46996 68152 47016
rect 68152 46996 68154 47016
rect 68098 46960 68154 46996
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 65660 46266 65716 46268
rect 65740 46266 65796 46268
rect 65820 46266 65876 46268
rect 65900 46266 65956 46268
rect 65660 46214 65706 46266
rect 65706 46214 65716 46266
rect 65740 46214 65770 46266
rect 65770 46214 65782 46266
rect 65782 46214 65796 46266
rect 65820 46214 65834 46266
rect 65834 46214 65846 46266
rect 65846 46214 65876 46266
rect 65900 46214 65910 46266
rect 65910 46214 65956 46266
rect 65660 46212 65716 46214
rect 65740 46212 65796 46214
rect 65820 46212 65876 46214
rect 65900 46212 65956 46214
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 68098 45600 68154 45656
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 65660 45178 65716 45180
rect 65740 45178 65796 45180
rect 65820 45178 65876 45180
rect 65900 45178 65956 45180
rect 65660 45126 65706 45178
rect 65706 45126 65716 45178
rect 65740 45126 65770 45178
rect 65770 45126 65782 45178
rect 65782 45126 65796 45178
rect 65820 45126 65834 45178
rect 65834 45126 65846 45178
rect 65846 45126 65876 45178
rect 65900 45126 65910 45178
rect 65910 45126 65956 45178
rect 65660 45124 65716 45126
rect 65740 45124 65796 45126
rect 65820 45124 65876 45126
rect 65900 45124 65956 45126
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 67638 44260 67694 44296
rect 67638 44240 67640 44260
rect 67640 44240 67692 44260
rect 67692 44240 67694 44260
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 65660 44090 65716 44092
rect 65740 44090 65796 44092
rect 65820 44090 65876 44092
rect 65900 44090 65956 44092
rect 65660 44038 65706 44090
rect 65706 44038 65716 44090
rect 65740 44038 65770 44090
rect 65770 44038 65782 44090
rect 65782 44038 65796 44090
rect 65820 44038 65834 44090
rect 65834 44038 65846 44090
rect 65846 44038 65876 44090
rect 65900 44038 65910 44090
rect 65910 44038 65956 44090
rect 65660 44036 65716 44038
rect 65740 44036 65796 44038
rect 65820 44036 65876 44038
rect 65900 44036 65956 44038
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 65660 43002 65716 43004
rect 65740 43002 65796 43004
rect 65820 43002 65876 43004
rect 65900 43002 65956 43004
rect 65660 42950 65706 43002
rect 65706 42950 65716 43002
rect 65740 42950 65770 43002
rect 65770 42950 65782 43002
rect 65782 42950 65796 43002
rect 65820 42950 65834 43002
rect 65834 42950 65846 43002
rect 65846 42950 65876 43002
rect 65900 42950 65910 43002
rect 65910 42950 65956 43002
rect 65660 42948 65716 42950
rect 65740 42948 65796 42950
rect 65820 42948 65876 42950
rect 65900 42948 65956 42950
rect 67638 42880 67694 42936
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 65660 41914 65716 41916
rect 65740 41914 65796 41916
rect 65820 41914 65876 41916
rect 65900 41914 65956 41916
rect 65660 41862 65706 41914
rect 65706 41862 65716 41914
rect 65740 41862 65770 41914
rect 65770 41862 65782 41914
rect 65782 41862 65796 41914
rect 65820 41862 65834 41914
rect 65834 41862 65846 41914
rect 65846 41862 65876 41914
rect 65900 41862 65910 41914
rect 65910 41862 65956 41914
rect 65660 41860 65716 41862
rect 65740 41860 65796 41862
rect 65820 41860 65876 41862
rect 65900 41860 65956 41862
rect 68098 41556 68100 41576
rect 68100 41556 68152 41576
rect 68152 41556 68154 41576
rect 68098 41520 68154 41556
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 65660 40826 65716 40828
rect 65740 40826 65796 40828
rect 65820 40826 65876 40828
rect 65900 40826 65956 40828
rect 65660 40774 65706 40826
rect 65706 40774 65716 40826
rect 65740 40774 65770 40826
rect 65770 40774 65782 40826
rect 65782 40774 65796 40826
rect 65820 40774 65834 40826
rect 65834 40774 65846 40826
rect 65846 40774 65876 40826
rect 65900 40774 65910 40826
rect 65910 40774 65956 40826
rect 65660 40772 65716 40774
rect 65740 40772 65796 40774
rect 65820 40772 65876 40774
rect 65900 40772 65956 40774
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 68098 40160 68154 40216
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 65660 39738 65716 39740
rect 65740 39738 65796 39740
rect 65820 39738 65876 39740
rect 65900 39738 65956 39740
rect 65660 39686 65706 39738
rect 65706 39686 65716 39738
rect 65740 39686 65770 39738
rect 65770 39686 65782 39738
rect 65782 39686 65796 39738
rect 65820 39686 65834 39738
rect 65834 39686 65846 39738
rect 65846 39686 65876 39738
rect 65900 39686 65910 39738
rect 65910 39686 65956 39738
rect 65660 39684 65716 39686
rect 65740 39684 65796 39686
rect 65820 39684 65876 39686
rect 65900 39684 65956 39686
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 67638 38820 67694 38856
rect 67638 38800 67640 38820
rect 67640 38800 67692 38820
rect 67692 38800 67694 38820
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 65660 38650 65716 38652
rect 65740 38650 65796 38652
rect 65820 38650 65876 38652
rect 65900 38650 65956 38652
rect 65660 38598 65706 38650
rect 65706 38598 65716 38650
rect 65740 38598 65770 38650
rect 65770 38598 65782 38650
rect 65782 38598 65796 38650
rect 65820 38598 65834 38650
rect 65834 38598 65846 38650
rect 65846 38598 65876 38650
rect 65900 38598 65910 38650
rect 65910 38598 65956 38650
rect 65660 38596 65716 38598
rect 65740 38596 65796 38598
rect 65820 38596 65876 38598
rect 65900 38596 65956 38598
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 65660 37562 65716 37564
rect 65740 37562 65796 37564
rect 65820 37562 65876 37564
rect 65900 37562 65956 37564
rect 65660 37510 65706 37562
rect 65706 37510 65716 37562
rect 65740 37510 65770 37562
rect 65770 37510 65782 37562
rect 65782 37510 65796 37562
rect 65820 37510 65834 37562
rect 65834 37510 65846 37562
rect 65846 37510 65876 37562
rect 65900 37510 65910 37562
rect 65910 37510 65956 37562
rect 65660 37508 65716 37510
rect 65740 37508 65796 37510
rect 65820 37508 65876 37510
rect 65900 37508 65956 37510
rect 67638 37440 67694 37496
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 65660 36474 65716 36476
rect 65740 36474 65796 36476
rect 65820 36474 65876 36476
rect 65900 36474 65956 36476
rect 65660 36422 65706 36474
rect 65706 36422 65716 36474
rect 65740 36422 65770 36474
rect 65770 36422 65782 36474
rect 65782 36422 65796 36474
rect 65820 36422 65834 36474
rect 65834 36422 65846 36474
rect 65846 36422 65876 36474
rect 65900 36422 65910 36474
rect 65910 36422 65956 36474
rect 65660 36420 65716 36422
rect 65740 36420 65796 36422
rect 65820 36420 65876 36422
rect 65900 36420 65956 36422
rect 68098 36116 68100 36136
rect 68100 36116 68152 36136
rect 68152 36116 68154 36136
rect 68098 36080 68154 36116
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 65660 35386 65716 35388
rect 65740 35386 65796 35388
rect 65820 35386 65876 35388
rect 65900 35386 65956 35388
rect 65660 35334 65706 35386
rect 65706 35334 65716 35386
rect 65740 35334 65770 35386
rect 65770 35334 65782 35386
rect 65782 35334 65796 35386
rect 65820 35334 65834 35386
rect 65834 35334 65846 35386
rect 65846 35334 65876 35386
rect 65900 35334 65910 35386
rect 65910 35334 65956 35386
rect 65660 35332 65716 35334
rect 65740 35332 65796 35334
rect 65820 35332 65876 35334
rect 65900 35332 65956 35334
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 68098 34720 68154 34776
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 65660 34298 65716 34300
rect 65740 34298 65796 34300
rect 65820 34298 65876 34300
rect 65900 34298 65956 34300
rect 65660 34246 65706 34298
rect 65706 34246 65716 34298
rect 65740 34246 65770 34298
rect 65770 34246 65782 34298
rect 65782 34246 65796 34298
rect 65820 34246 65834 34298
rect 65834 34246 65846 34298
rect 65846 34246 65876 34298
rect 65900 34246 65910 34298
rect 65910 34246 65956 34298
rect 65660 34244 65716 34246
rect 65740 34244 65796 34246
rect 65820 34244 65876 34246
rect 65900 34244 65956 34246
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 67638 33380 67694 33416
rect 67638 33360 67640 33380
rect 67640 33360 67692 33380
rect 67692 33360 67694 33380
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 65660 33210 65716 33212
rect 65740 33210 65796 33212
rect 65820 33210 65876 33212
rect 65900 33210 65956 33212
rect 65660 33158 65706 33210
rect 65706 33158 65716 33210
rect 65740 33158 65770 33210
rect 65770 33158 65782 33210
rect 65782 33158 65796 33210
rect 65820 33158 65834 33210
rect 65834 33158 65846 33210
rect 65846 33158 65876 33210
rect 65900 33158 65910 33210
rect 65910 33158 65956 33210
rect 65660 33156 65716 33158
rect 65740 33156 65796 33158
rect 65820 33156 65876 33158
rect 65900 33156 65956 33158
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 5814 30116 5870 30152
rect 5814 30096 5816 30116
rect 5816 30096 5868 30116
rect 5868 30096 5870 30116
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 7286 29588 7288 29608
rect 7288 29588 7340 29608
rect 7340 29588 7342 29608
rect 7286 29552 7342 29588
rect 5446 29028 5502 29064
rect 5446 29008 5448 29028
rect 5448 29008 5500 29028
rect 5500 29008 5502 29028
rect 1950 20304 2006 20360
rect 2134 19352 2190 19408
rect 1858 17196 1914 17232
rect 1858 17176 1860 17196
rect 1860 17176 1912 17196
rect 1912 17176 1914 17196
rect 2502 13368 2558 13424
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4618 22500 4674 22536
rect 4618 22480 4620 22500
rect 4620 22480 4672 22500
rect 4672 22480 4674 22500
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 5170 23024 5226 23080
rect 5078 22072 5134 22128
rect 2226 3340 2228 3360
rect 2228 3340 2280 3360
rect 2280 3340 2282 3360
rect 2226 3304 2282 3340
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4158 20324 4214 20360
rect 4158 20304 4160 20324
rect 4160 20304 4212 20324
rect 4212 20304 4214 20324
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4802 19352 4858 19408
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 8114 29552 8170 29608
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 5446 15972 5502 16008
rect 5446 15952 5448 15972
rect 5448 15952 5500 15972
rect 5500 15952 5502 15972
rect 5630 14884 5686 14920
rect 5630 14864 5632 14884
rect 5632 14864 5684 14884
rect 5684 14864 5686 14884
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 3238 5752 3294 5808
rect 2410 2352 2466 2408
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4250 3984 4306 4040
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 5078 3712 5134 3768
rect 5262 3032 5318 3088
rect 6274 17196 6330 17232
rect 6274 17176 6276 17196
rect 6276 17176 6328 17196
rect 6328 17176 6330 17196
rect 7010 16496 7066 16552
rect 7102 13388 7158 13424
rect 7102 13368 7104 13388
rect 7104 13368 7156 13388
rect 7156 13368 7158 13388
rect 6734 5752 6790 5808
rect 6734 3848 6790 3904
rect 6550 2896 6606 2952
rect 5630 2760 5686 2816
rect 5446 2488 5502 2544
rect 3330 2216 3386 2272
rect 7194 3848 7250 3904
rect 9586 26852 9642 26888
rect 9586 26832 9588 26852
rect 9588 26832 9640 26852
rect 9640 26832 9642 26852
rect 9034 20440 9090 20496
rect 8482 19372 8538 19408
rect 9218 19388 9220 19408
rect 9220 19388 9272 19408
rect 9272 19388 9274 19408
rect 8482 19352 8484 19372
rect 8484 19352 8536 19372
rect 8536 19352 8538 19372
rect 9218 19352 9274 19388
rect 7562 12144 7618 12200
rect 7838 8372 7840 8392
rect 7840 8372 7892 8392
rect 7892 8372 7894 8392
rect 7838 8336 7894 8372
rect 7470 4684 7526 4720
rect 7470 4664 7472 4684
rect 7472 4664 7524 4684
rect 7524 4664 7526 4684
rect 8390 4428 8392 4448
rect 8392 4428 8444 4448
rect 8444 4428 8446 4448
rect 8390 4392 8446 4428
rect 7930 3848 7986 3904
rect 7930 3612 7932 3632
rect 7932 3612 7984 3632
rect 7984 3612 7986 3632
rect 7930 3576 7986 3612
rect 7286 3168 7342 3224
rect 7654 2624 7710 2680
rect 8390 3612 8392 3632
rect 8392 3612 8444 3632
rect 8444 3612 8446 3632
rect 8390 3576 8446 3612
rect 12990 25220 13046 25256
rect 12990 25200 12992 25220
rect 12992 25200 13044 25220
rect 13044 25200 13046 25220
rect 11058 22072 11114 22128
rect 10966 21412 11022 21448
rect 10966 21392 10968 21412
rect 10968 21392 11020 21412
rect 11020 21392 11022 21412
rect 11058 17584 11114 17640
rect 9954 13776 10010 13832
rect 10046 10648 10102 10704
rect 9770 9424 9826 9480
rect 6826 2080 6882 2136
rect 9678 6568 9734 6624
rect 9770 4140 9826 4176
rect 9770 4120 9772 4140
rect 9772 4120 9824 4140
rect 9824 4120 9826 4140
rect 9678 3576 9734 3632
rect 10046 3304 10102 3360
rect 10046 2216 10102 2272
rect 10782 12280 10838 12336
rect 12162 15444 12164 15464
rect 12164 15444 12216 15464
rect 12216 15444 12218 15464
rect 12162 15408 12218 15444
rect 12070 13232 12126 13288
rect 12070 12708 12126 12744
rect 12070 12688 12072 12708
rect 12072 12688 12124 12708
rect 12124 12688 12126 12708
rect 10690 10532 10746 10568
rect 10690 10512 10692 10532
rect 10692 10512 10744 10532
rect 10744 10512 10746 10532
rect 12070 11620 12126 11656
rect 12070 11600 12072 11620
rect 12072 11600 12124 11620
rect 12124 11600 12126 11620
rect 10506 9324 10508 9344
rect 10508 9324 10560 9344
rect 10560 9324 10562 9344
rect 10506 9288 10562 9324
rect 10966 9968 11022 10024
rect 10414 3460 10470 3496
rect 10414 3440 10416 3460
rect 10416 3440 10468 3460
rect 10468 3440 10470 3460
rect 11610 9560 11666 9616
rect 10966 3712 11022 3768
rect 10414 2216 10470 2272
rect 12438 12144 12494 12200
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 13910 22480 13966 22536
rect 13450 20168 13506 20224
rect 12622 12180 12624 12200
rect 12624 12180 12676 12200
rect 12676 12180 12678 12200
rect 12622 12144 12678 12180
rect 11610 4392 11666 4448
rect 11518 2760 11574 2816
rect 12254 2896 12310 2952
rect 14186 12588 14188 12608
rect 14188 12588 14240 12608
rect 14240 12588 14242 12608
rect 14186 12552 14242 12588
rect 15382 23044 15438 23080
rect 15382 23024 15384 23044
rect 15384 23024 15436 23044
rect 15436 23024 15438 23044
rect 14186 11892 14242 11928
rect 14186 11872 14188 11892
rect 14188 11872 14240 11892
rect 14240 11872 14242 11892
rect 12898 3984 12954 4040
rect 13910 10376 13966 10432
rect 13542 8336 13598 8392
rect 13542 6568 13598 6624
rect 13634 6160 13690 6216
rect 13542 5616 13598 5672
rect 13358 4800 13414 4856
rect 13358 4120 13414 4176
rect 13450 3168 13506 3224
rect 13266 3032 13322 3088
rect 13266 2916 13322 2952
rect 13266 2896 13268 2916
rect 13268 2896 13320 2916
rect 13320 2896 13322 2916
rect 13266 2760 13322 2816
rect 12990 2352 13046 2408
rect 14370 9560 14426 9616
rect 15290 22208 15346 22264
rect 15842 20032 15898 20088
rect 17314 30096 17370 30152
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 17130 29008 17186 29064
rect 17130 26832 17186 26888
rect 17406 26288 17462 26344
rect 17406 25220 17462 25256
rect 17406 25200 17408 25220
rect 17408 25200 17460 25220
rect 17460 25200 17462 25220
rect 17682 24928 17738 24984
rect 17314 23724 17370 23760
rect 17314 23704 17316 23724
rect 17316 23704 17368 23724
rect 17368 23704 17370 23724
rect 15842 17196 15898 17232
rect 15842 17176 15844 17196
rect 15844 17176 15896 17196
rect 15896 17176 15898 17196
rect 13726 4936 13782 4992
rect 13726 3984 13782 4040
rect 14370 3576 14426 3632
rect 14922 5616 14978 5672
rect 14830 2488 14886 2544
rect 17130 18284 17186 18320
rect 17130 18264 17132 18284
rect 17132 18264 17184 18284
rect 17184 18264 17186 18284
rect 16578 13812 16580 13832
rect 16580 13812 16632 13832
rect 16632 13812 16634 13832
rect 16578 13776 16634 13812
rect 16670 13676 16672 13696
rect 16672 13676 16724 13696
rect 16724 13676 16726 13696
rect 16670 13640 16726 13676
rect 16762 13404 16764 13424
rect 16764 13404 16816 13424
rect 16816 13404 16818 13424
rect 16762 13368 16818 13404
rect 17314 18128 17370 18184
rect 15106 3848 15162 3904
rect 16854 9424 16910 9480
rect 16026 4684 16082 4720
rect 16026 4664 16028 4684
rect 16028 4664 16080 4684
rect 16080 4664 16082 4684
rect 17498 12144 17554 12200
rect 17498 10920 17554 10976
rect 17682 13504 17738 13560
rect 17682 9560 17738 9616
rect 17130 9152 17186 9208
rect 18234 23704 18290 23760
rect 18234 11872 18290 11928
rect 17958 9560 18014 9616
rect 17774 9016 17830 9072
rect 19614 29572 19670 29608
rect 19614 29552 19616 29572
rect 19616 29552 19668 29572
rect 19668 29552 19670 29572
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 18970 20204 18972 20224
rect 18972 20204 19024 20224
rect 19024 20204 19026 20224
rect 18970 20168 19026 20204
rect 18970 19372 19026 19408
rect 18970 19352 18972 19372
rect 18972 19352 19024 19372
rect 19024 19352 19026 19372
rect 19338 23296 19394 23352
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19798 20304 19854 20360
rect 19522 20032 19578 20088
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19062 15680 19118 15736
rect 18326 10240 18382 10296
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 18418 9424 18474 9480
rect 17222 4936 17278 4992
rect 17130 2896 17186 2952
rect 16762 2080 16818 2136
rect 17682 4800 17738 4856
rect 17590 2760 17646 2816
rect 17774 2896 17830 2952
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19798 12844 19854 12880
rect 19798 12824 19800 12844
rect 19800 12824 19852 12844
rect 19852 12824 19854 12844
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19706 11772 19708 11792
rect 19708 11772 19760 11792
rect 19760 11772 19762 11792
rect 19706 11736 19762 11772
rect 19706 11328 19762 11384
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 65660 32122 65716 32124
rect 65740 32122 65796 32124
rect 65820 32122 65876 32124
rect 65900 32122 65956 32124
rect 65660 32070 65706 32122
rect 65706 32070 65716 32122
rect 65740 32070 65770 32122
rect 65770 32070 65782 32122
rect 65782 32070 65796 32122
rect 65820 32070 65834 32122
rect 65834 32070 65846 32122
rect 65846 32070 65876 32122
rect 65900 32070 65910 32122
rect 65910 32070 65956 32122
rect 65660 32068 65716 32070
rect 65740 32068 65796 32070
rect 65820 32068 65876 32070
rect 65900 32068 65956 32070
rect 67638 32000 67694 32056
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 23202 27412 23204 27432
rect 23204 27412 23256 27432
rect 23256 27412 23258 27432
rect 23202 27376 23258 27412
rect 21914 21972 21916 21992
rect 21916 21972 21968 21992
rect 21968 21972 21970 21992
rect 21914 21936 21970 21972
rect 21178 19252 21180 19272
rect 21180 19252 21232 19272
rect 21232 19252 21234 19272
rect 21178 19216 21234 19252
rect 20534 17992 20590 18048
rect 20166 12824 20222 12880
rect 19614 11212 19670 11248
rect 19614 11192 19616 11212
rect 19616 11192 19668 11212
rect 19668 11192 19670 11212
rect 20258 11736 20314 11792
rect 20074 11328 20130 11384
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19706 10124 19762 10160
rect 19706 10104 19708 10124
rect 19708 10104 19760 10124
rect 19760 10104 19762 10124
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19982 9696 20038 9752
rect 20166 9832 20222 9888
rect 19430 8880 19486 8936
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19338 8472 19394 8528
rect 20994 18400 21050 18456
rect 20718 13504 20774 13560
rect 20810 9696 20866 9752
rect 20258 8472 20314 8528
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19982 6160 20038 6216
rect 19614 5652 19616 5672
rect 19616 5652 19668 5672
rect 19668 5652 19670 5672
rect 19614 5616 19670 5652
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19246 3576 19302 3632
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 20074 3460 20130 3496
rect 20074 3440 20076 3460
rect 20076 3440 20128 3460
rect 20128 3440 20130 3460
rect 21086 18300 21088 18320
rect 21088 18300 21140 18320
rect 21140 18300 21142 18320
rect 21086 18264 21142 18300
rect 21362 17604 21418 17640
rect 21362 17584 21364 17604
rect 21364 17584 21416 17604
rect 21416 17584 21418 17604
rect 21822 20168 21878 20224
rect 21822 16360 21878 16416
rect 22006 14864 22062 14920
rect 22742 20884 22744 20904
rect 22744 20884 22796 20904
rect 22796 20884 22798 20904
rect 22742 20848 22798 20884
rect 22558 19352 22614 19408
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 65660 31034 65716 31036
rect 65740 31034 65796 31036
rect 65820 31034 65876 31036
rect 65900 31034 65956 31036
rect 65660 30982 65706 31034
rect 65706 30982 65716 31034
rect 65740 30982 65770 31034
rect 65770 30982 65782 31034
rect 65782 30982 65796 31034
rect 65820 30982 65834 31034
rect 65834 30982 65846 31034
rect 65846 30982 65876 31034
rect 65900 30982 65910 31034
rect 65910 30982 65956 31034
rect 65660 30980 65716 30982
rect 65740 30980 65796 30982
rect 65820 30980 65876 30982
rect 65900 30980 65956 30982
rect 68098 30676 68100 30696
rect 68100 30676 68152 30696
rect 68152 30676 68154 30696
rect 68098 30640 68154 30676
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 65660 29946 65716 29948
rect 65740 29946 65796 29948
rect 65820 29946 65876 29948
rect 65900 29946 65956 29948
rect 65660 29894 65706 29946
rect 65706 29894 65716 29946
rect 65740 29894 65770 29946
rect 65770 29894 65782 29946
rect 65782 29894 65796 29946
rect 65820 29894 65834 29946
rect 65834 29894 65846 29946
rect 65846 29894 65876 29946
rect 65900 29894 65910 29946
rect 65910 29894 65956 29946
rect 65660 29892 65716 29894
rect 65740 29892 65796 29894
rect 65820 29892 65876 29894
rect 65900 29892 65956 29894
rect 24214 27412 24216 27432
rect 24216 27412 24268 27432
rect 24268 27412 24270 27432
rect 24214 27376 24270 27412
rect 23478 21392 23534 21448
rect 23570 20476 23572 20496
rect 23572 20476 23624 20496
rect 23624 20476 23626 20496
rect 23570 20440 23626 20476
rect 23110 17176 23166 17232
rect 23202 16632 23258 16688
rect 22282 15952 22338 16008
rect 22282 15020 22338 15056
rect 22282 15000 22284 15020
rect 22284 15000 22336 15020
rect 22336 15000 22338 15020
rect 21362 11092 21364 11112
rect 21364 11092 21416 11112
rect 21416 11092 21418 11112
rect 21362 11056 21418 11092
rect 23202 15408 23258 15464
rect 22650 10240 22706 10296
rect 23570 13232 23626 13288
rect 23478 12688 23534 12744
rect 22466 8880 22522 8936
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 68098 29280 68154 29336
rect 24858 15680 24914 15736
rect 24950 13932 25006 13968
rect 24950 13912 24952 13932
rect 24952 13912 25004 13932
rect 25004 13912 25006 13932
rect 24674 12824 24730 12880
rect 25410 20884 25412 20904
rect 25412 20884 25464 20904
rect 25464 20884 25466 20904
rect 25410 20848 25466 20884
rect 25686 20576 25742 20632
rect 26146 23296 26202 23352
rect 24950 11192 25006 11248
rect 24950 10784 25006 10840
rect 24950 10376 25006 10432
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 65660 28858 65716 28860
rect 65740 28858 65796 28860
rect 65820 28858 65876 28860
rect 65900 28858 65956 28860
rect 65660 28806 65706 28858
rect 65706 28806 65716 28858
rect 65740 28806 65770 28858
rect 65770 28806 65782 28858
rect 65782 28806 65796 28858
rect 65820 28806 65834 28858
rect 65834 28806 65846 28858
rect 65846 28806 65876 28858
rect 65900 28806 65910 28858
rect 65910 28806 65956 28858
rect 65660 28804 65716 28806
rect 65740 28804 65796 28806
rect 65820 28804 65876 28806
rect 65900 28804 65956 28806
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 26330 18400 26386 18456
rect 26514 17992 26570 18048
rect 26514 17212 26516 17232
rect 26516 17212 26568 17232
rect 26568 17212 26570 17232
rect 26514 17176 26570 17212
rect 26330 16224 26386 16280
rect 27250 16496 27306 16552
rect 25410 10784 25466 10840
rect 24490 9152 24546 9208
rect 24214 8336 24270 8392
rect 26974 11600 27030 11656
rect 27710 14184 27766 14240
rect 27894 13368 27950 13424
rect 67638 27940 67694 27976
rect 67638 27920 67640 27940
rect 67640 27920 67692 27940
rect 67692 27920 67694 27940
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 65660 27770 65716 27772
rect 65740 27770 65796 27772
rect 65820 27770 65876 27772
rect 65900 27770 65956 27772
rect 65660 27718 65706 27770
rect 65706 27718 65716 27770
rect 65740 27718 65770 27770
rect 65770 27718 65782 27770
rect 65782 27718 65796 27770
rect 65820 27718 65834 27770
rect 65834 27718 65846 27770
rect 65846 27718 65876 27770
rect 65900 27718 65910 27770
rect 65910 27718 65956 27770
rect 65660 27716 65716 27718
rect 65740 27716 65796 27718
rect 65820 27716 65876 27718
rect 65900 27716 65956 27718
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 65660 26682 65716 26684
rect 65740 26682 65796 26684
rect 65820 26682 65876 26684
rect 65900 26682 65956 26684
rect 65660 26630 65706 26682
rect 65706 26630 65716 26682
rect 65740 26630 65770 26682
rect 65770 26630 65782 26682
rect 65782 26630 65796 26682
rect 65820 26630 65834 26682
rect 65834 26630 65846 26682
rect 65846 26630 65876 26682
rect 65900 26630 65910 26682
rect 65910 26630 65956 26682
rect 65660 26628 65716 26630
rect 65740 26628 65796 26630
rect 65820 26628 65876 26630
rect 65900 26628 65956 26630
rect 67638 26560 67694 26616
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 28630 17212 28632 17232
rect 28632 17212 28684 17232
rect 28684 17212 28686 17232
rect 28630 17176 28686 17212
rect 28630 16496 28686 16552
rect 28722 13368 28778 13424
rect 29642 17448 29698 17504
rect 27986 12280 28042 12336
rect 28446 12144 28502 12200
rect 27986 9288 28042 9344
rect 28814 10668 28870 10704
rect 28814 10648 28816 10668
rect 28816 10648 28868 10668
rect 28868 10648 28870 10668
rect 28998 10512 29054 10568
rect 28538 10140 28540 10160
rect 28540 10140 28592 10160
rect 28592 10140 28594 10160
rect 28538 10104 28594 10140
rect 28446 9560 28502 9616
rect 28906 9968 28962 10024
rect 29366 9016 29422 9072
rect 30562 21936 30618 21992
rect 30378 16360 30434 16416
rect 30838 19216 30894 19272
rect 31022 18128 31078 18184
rect 31114 16516 31170 16552
rect 31114 16496 31116 16516
rect 31116 16496 31168 16516
rect 31168 16496 31170 16516
rect 31482 21936 31538 21992
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 65660 25594 65716 25596
rect 65740 25594 65796 25596
rect 65820 25594 65876 25596
rect 65900 25594 65956 25596
rect 65660 25542 65706 25594
rect 65706 25542 65716 25594
rect 65740 25542 65770 25594
rect 65770 25542 65782 25594
rect 65782 25542 65796 25594
rect 65820 25542 65834 25594
rect 65834 25542 65846 25594
rect 65846 25542 65876 25594
rect 65900 25542 65910 25594
rect 65910 25542 65956 25594
rect 65660 25540 65716 25542
rect 65740 25540 65796 25542
rect 65820 25540 65876 25542
rect 65900 25540 65956 25542
rect 68098 25236 68100 25256
rect 68100 25236 68152 25256
rect 68152 25236 68154 25256
rect 68098 25200 68154 25236
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 65660 24506 65716 24508
rect 65740 24506 65796 24508
rect 65820 24506 65876 24508
rect 65900 24506 65956 24508
rect 65660 24454 65706 24506
rect 65706 24454 65716 24506
rect 65740 24454 65770 24506
rect 65770 24454 65782 24506
rect 65782 24454 65796 24506
rect 65820 24454 65834 24506
rect 65834 24454 65846 24506
rect 65846 24454 65876 24506
rect 65900 24454 65910 24506
rect 65910 24454 65956 24506
rect 65660 24452 65716 24454
rect 65740 24452 65796 24454
rect 65820 24452 65876 24454
rect 65900 24452 65956 24454
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 68098 23840 68154 23896
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 65660 23418 65716 23420
rect 65740 23418 65796 23420
rect 65820 23418 65876 23420
rect 65900 23418 65956 23420
rect 65660 23366 65706 23418
rect 65706 23366 65716 23418
rect 65740 23366 65770 23418
rect 65770 23366 65782 23418
rect 65782 23366 65796 23418
rect 65820 23366 65834 23418
rect 65834 23366 65846 23418
rect 65846 23366 65876 23418
rect 65900 23366 65910 23418
rect 65910 23366 65956 23418
rect 65660 23364 65716 23366
rect 65740 23364 65796 23366
rect 65820 23364 65876 23366
rect 65900 23364 65956 23366
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 67638 22500 67694 22536
rect 67638 22480 67640 22500
rect 67640 22480 67692 22500
rect 67692 22480 67694 22500
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 65660 22330 65716 22332
rect 65740 22330 65796 22332
rect 65820 22330 65876 22332
rect 65900 22330 65956 22332
rect 65660 22278 65706 22330
rect 65706 22278 65716 22330
rect 65740 22278 65770 22330
rect 65770 22278 65782 22330
rect 65782 22278 65796 22330
rect 65820 22278 65834 22330
rect 65834 22278 65846 22330
rect 65846 22278 65876 22330
rect 65900 22278 65910 22330
rect 65910 22278 65956 22330
rect 65660 22276 65716 22278
rect 65740 22276 65796 22278
rect 65820 22276 65876 22278
rect 65900 22276 65956 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 33322 18300 33324 18320
rect 33324 18300 33376 18320
rect 33376 18300 33378 18320
rect 33322 18264 33378 18300
rect 30838 9172 30894 9208
rect 30838 9152 30840 9172
rect 30840 9152 30892 9172
rect 30892 9152 30894 9172
rect 32954 14220 32956 14240
rect 32956 14220 33008 14240
rect 33008 14220 33010 14240
rect 32954 14184 33010 14220
rect 33046 13368 33102 13424
rect 33690 16224 33746 16280
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 65660 21242 65716 21244
rect 65740 21242 65796 21244
rect 65820 21242 65876 21244
rect 65900 21242 65956 21244
rect 65660 21190 65706 21242
rect 65706 21190 65716 21242
rect 65740 21190 65770 21242
rect 65770 21190 65782 21242
rect 65782 21190 65796 21242
rect 65820 21190 65834 21242
rect 65834 21190 65846 21242
rect 65846 21190 65876 21242
rect 65900 21190 65910 21242
rect 65910 21190 65956 21242
rect 65660 21188 65716 21190
rect 65740 21188 65796 21190
rect 65820 21188 65876 21190
rect 65900 21188 65956 21190
rect 67638 21120 67694 21176
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34702 13912 34758 13968
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 36634 17448 36690 17504
rect 35990 15272 36046 15328
rect 35990 15000 36046 15056
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 33874 8356 33930 8392
rect 33874 8336 33876 8356
rect 33876 8336 33928 8356
rect 33928 8336 33930 8356
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 26330 2896 26386 2952
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 65660 20154 65716 20156
rect 65740 20154 65796 20156
rect 65820 20154 65876 20156
rect 65900 20154 65956 20156
rect 65660 20102 65706 20154
rect 65706 20102 65716 20154
rect 65740 20102 65770 20154
rect 65770 20102 65782 20154
rect 65782 20102 65796 20154
rect 65820 20102 65834 20154
rect 65834 20102 65846 20154
rect 65846 20102 65876 20154
rect 65900 20102 65910 20154
rect 65910 20102 65956 20154
rect 65660 20100 65716 20102
rect 65740 20100 65796 20102
rect 65820 20100 65876 20102
rect 65900 20100 65956 20102
rect 68098 19796 68100 19816
rect 68100 19796 68152 19816
rect 68152 19796 68154 19816
rect 38014 17620 38016 17640
rect 38016 17620 38068 17640
rect 38068 17620 38070 17640
rect 38014 17584 38070 17620
rect 37922 16496 37978 16552
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 68098 19760 68154 19796
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 65660 19066 65716 19068
rect 65740 19066 65796 19068
rect 65820 19066 65876 19068
rect 65900 19066 65956 19068
rect 65660 19014 65706 19066
rect 65706 19014 65716 19066
rect 65740 19014 65770 19066
rect 65770 19014 65782 19066
rect 65782 19014 65796 19066
rect 65820 19014 65834 19066
rect 65834 19014 65846 19066
rect 65846 19014 65876 19066
rect 65900 19014 65910 19066
rect 65910 19014 65956 19066
rect 65660 19012 65716 19014
rect 65740 19012 65796 19014
rect 65820 19012 65876 19014
rect 65900 19012 65956 19014
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 68098 18400 68154 18456
rect 65660 17978 65716 17980
rect 65740 17978 65796 17980
rect 65820 17978 65876 17980
rect 65900 17978 65956 17980
rect 65660 17926 65706 17978
rect 65706 17926 65716 17978
rect 65740 17926 65770 17978
rect 65770 17926 65782 17978
rect 65782 17926 65796 17978
rect 65820 17926 65834 17978
rect 65834 17926 65846 17978
rect 65846 17926 65876 17978
rect 65900 17926 65910 17978
rect 65910 17926 65956 17978
rect 65660 17924 65716 17926
rect 65740 17924 65796 17926
rect 65820 17924 65876 17926
rect 65900 17924 65956 17926
rect 39302 17604 39358 17640
rect 39302 17584 39304 17604
rect 39304 17584 39356 17604
rect 39356 17584 39358 17604
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 67638 17060 67694 17096
rect 67638 17040 67640 17060
rect 67640 17040 67692 17060
rect 67692 17040 67694 17060
rect 65660 16890 65716 16892
rect 65740 16890 65796 16892
rect 65820 16890 65876 16892
rect 65900 16890 65956 16892
rect 65660 16838 65706 16890
rect 65706 16838 65716 16890
rect 65740 16838 65770 16890
rect 65770 16838 65782 16890
rect 65782 16838 65796 16890
rect 65820 16838 65834 16890
rect 65834 16838 65846 16890
rect 65846 16838 65876 16890
rect 65900 16838 65910 16890
rect 65910 16838 65956 16890
rect 65660 16836 65716 16838
rect 65740 16836 65796 16838
rect 65820 16836 65876 16838
rect 65900 16836 65956 16838
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 65660 15802 65716 15804
rect 65740 15802 65796 15804
rect 65820 15802 65876 15804
rect 65900 15802 65956 15804
rect 65660 15750 65706 15802
rect 65706 15750 65716 15802
rect 65740 15750 65770 15802
rect 65770 15750 65782 15802
rect 65782 15750 65796 15802
rect 65820 15750 65834 15802
rect 65834 15750 65846 15802
rect 65846 15750 65876 15802
rect 65900 15750 65910 15802
rect 65910 15750 65956 15802
rect 65660 15748 65716 15750
rect 65740 15748 65796 15750
rect 65820 15748 65876 15750
rect 65900 15748 65956 15750
rect 67638 15680 67694 15736
rect 38934 15272 38990 15328
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 65660 14714 65716 14716
rect 65740 14714 65796 14716
rect 65820 14714 65876 14716
rect 65900 14714 65956 14716
rect 65660 14662 65706 14714
rect 65706 14662 65716 14714
rect 65740 14662 65770 14714
rect 65770 14662 65782 14714
rect 65782 14662 65796 14714
rect 65820 14662 65834 14714
rect 65834 14662 65846 14714
rect 65846 14662 65876 14714
rect 65900 14662 65910 14714
rect 65910 14662 65956 14714
rect 65660 14660 65716 14662
rect 65740 14660 65796 14662
rect 65820 14660 65876 14662
rect 65900 14660 65956 14662
rect 68098 14356 68100 14376
rect 68100 14356 68152 14376
rect 68152 14356 68154 14376
rect 68098 14320 68154 14356
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 65660 13626 65716 13628
rect 65740 13626 65796 13628
rect 65820 13626 65876 13628
rect 65900 13626 65956 13628
rect 65660 13574 65706 13626
rect 65706 13574 65716 13626
rect 65740 13574 65770 13626
rect 65770 13574 65782 13626
rect 65782 13574 65796 13626
rect 65820 13574 65834 13626
rect 65834 13574 65846 13626
rect 65846 13574 65876 13626
rect 65900 13574 65910 13626
rect 65910 13574 65956 13626
rect 65660 13572 65716 13574
rect 65740 13572 65796 13574
rect 65820 13572 65876 13574
rect 65900 13572 65956 13574
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 68098 12960 68154 13016
rect 65660 12538 65716 12540
rect 65740 12538 65796 12540
rect 65820 12538 65876 12540
rect 65900 12538 65956 12540
rect 65660 12486 65706 12538
rect 65706 12486 65716 12538
rect 65740 12486 65770 12538
rect 65770 12486 65782 12538
rect 65782 12486 65796 12538
rect 65820 12486 65834 12538
rect 65834 12486 65846 12538
rect 65846 12486 65876 12538
rect 65900 12486 65910 12538
rect 65910 12486 65956 12538
rect 65660 12484 65716 12486
rect 65740 12484 65796 12486
rect 65820 12484 65876 12486
rect 65900 12484 65956 12486
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 67638 11620 67694 11656
rect 67638 11600 67640 11620
rect 67640 11600 67692 11620
rect 67692 11600 67694 11620
rect 65660 11450 65716 11452
rect 65740 11450 65796 11452
rect 65820 11450 65876 11452
rect 65900 11450 65956 11452
rect 65660 11398 65706 11450
rect 65706 11398 65716 11450
rect 65740 11398 65770 11450
rect 65770 11398 65782 11450
rect 65782 11398 65796 11450
rect 65820 11398 65834 11450
rect 65834 11398 65846 11450
rect 65846 11398 65876 11450
rect 65900 11398 65910 11450
rect 65910 11398 65956 11450
rect 65660 11396 65716 11398
rect 65740 11396 65796 11398
rect 65820 11396 65876 11398
rect 65900 11396 65956 11398
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 65660 10362 65716 10364
rect 65740 10362 65796 10364
rect 65820 10362 65876 10364
rect 65900 10362 65956 10364
rect 65660 10310 65706 10362
rect 65706 10310 65716 10362
rect 65740 10310 65770 10362
rect 65770 10310 65782 10362
rect 65782 10310 65796 10362
rect 65820 10310 65834 10362
rect 65834 10310 65846 10362
rect 65846 10310 65876 10362
rect 65900 10310 65910 10362
rect 65910 10310 65956 10362
rect 65660 10308 65716 10310
rect 65740 10308 65796 10310
rect 65820 10308 65876 10310
rect 65900 10308 65956 10310
rect 67638 10240 67694 10296
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 65660 9274 65716 9276
rect 65740 9274 65796 9276
rect 65820 9274 65876 9276
rect 65900 9274 65956 9276
rect 65660 9222 65706 9274
rect 65706 9222 65716 9274
rect 65740 9222 65770 9274
rect 65770 9222 65782 9274
rect 65782 9222 65796 9274
rect 65820 9222 65834 9274
rect 65834 9222 65846 9274
rect 65846 9222 65876 9274
rect 65900 9222 65910 9274
rect 65910 9222 65956 9274
rect 65660 9220 65716 9222
rect 65740 9220 65796 9222
rect 65820 9220 65876 9222
rect 65900 9220 65956 9222
rect 68098 8916 68100 8936
rect 68100 8916 68152 8936
rect 68152 8916 68154 8936
rect 68098 8880 68154 8916
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 65660 8186 65716 8188
rect 65740 8186 65796 8188
rect 65820 8186 65876 8188
rect 65900 8186 65956 8188
rect 65660 8134 65706 8186
rect 65706 8134 65716 8186
rect 65740 8134 65770 8186
rect 65770 8134 65782 8186
rect 65782 8134 65796 8186
rect 65820 8134 65834 8186
rect 65834 8134 65846 8186
rect 65846 8134 65876 8186
rect 65900 8134 65910 8186
rect 65910 8134 65956 8186
rect 65660 8132 65716 8134
rect 65740 8132 65796 8134
rect 65820 8132 65876 8134
rect 65900 8132 65956 8134
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 68098 7520 68154 7576
rect 65660 7098 65716 7100
rect 65740 7098 65796 7100
rect 65820 7098 65876 7100
rect 65900 7098 65956 7100
rect 65660 7046 65706 7098
rect 65706 7046 65716 7098
rect 65740 7046 65770 7098
rect 65770 7046 65782 7098
rect 65782 7046 65796 7098
rect 65820 7046 65834 7098
rect 65834 7046 65846 7098
rect 65846 7046 65876 7098
rect 65900 7046 65910 7098
rect 65910 7046 65956 7098
rect 65660 7044 65716 7046
rect 65740 7044 65796 7046
rect 65820 7044 65876 7046
rect 65900 7044 65956 7046
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 67638 6180 67694 6216
rect 67638 6160 67640 6180
rect 67640 6160 67692 6180
rect 67692 6160 67694 6180
rect 65660 6010 65716 6012
rect 65740 6010 65796 6012
rect 65820 6010 65876 6012
rect 65900 6010 65956 6012
rect 65660 5958 65706 6010
rect 65706 5958 65716 6010
rect 65740 5958 65770 6010
rect 65770 5958 65782 6010
rect 65782 5958 65796 6010
rect 65820 5958 65834 6010
rect 65834 5958 65846 6010
rect 65846 5958 65876 6010
rect 65900 5958 65910 6010
rect 65910 5958 65956 6010
rect 65660 5956 65716 5958
rect 65740 5956 65796 5958
rect 65820 5956 65876 5958
rect 65900 5956 65956 5958
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 57886 3168 57942 3224
rect 65660 4922 65716 4924
rect 65740 4922 65796 4924
rect 65820 4922 65876 4924
rect 65900 4922 65956 4924
rect 65660 4870 65706 4922
rect 65706 4870 65716 4922
rect 65740 4870 65770 4922
rect 65770 4870 65782 4922
rect 65782 4870 65796 4922
rect 65820 4870 65834 4922
rect 65834 4870 65846 4922
rect 65846 4870 65876 4922
rect 65900 4870 65910 4922
rect 65910 4870 65956 4922
rect 65660 4868 65716 4870
rect 65740 4868 65796 4870
rect 65820 4868 65876 4870
rect 65900 4868 65956 4870
rect 67638 4800 67694 4856
rect 65660 3834 65716 3836
rect 65740 3834 65796 3836
rect 65820 3834 65876 3836
rect 65900 3834 65956 3836
rect 65660 3782 65706 3834
rect 65706 3782 65716 3834
rect 65740 3782 65770 3834
rect 65770 3782 65782 3834
rect 65782 3782 65796 3834
rect 65820 3782 65834 3834
rect 65834 3782 65846 3834
rect 65846 3782 65876 3834
rect 65900 3782 65910 3834
rect 65910 3782 65956 3834
rect 65660 3780 65716 3782
rect 65740 3780 65796 3782
rect 65820 3780 65876 3782
rect 65900 3780 65956 3782
rect 68098 3476 68100 3496
rect 68100 3476 68152 3496
rect 68152 3476 68154 3496
rect 68098 3440 68154 3476
rect 60462 3168 60518 3224
rect 65660 2746 65716 2748
rect 65740 2746 65796 2748
rect 65820 2746 65876 2748
rect 65900 2746 65956 2748
rect 65660 2694 65706 2746
rect 65706 2694 65716 2746
rect 65740 2694 65770 2746
rect 65770 2694 65782 2746
rect 65782 2694 65796 2746
rect 65820 2694 65834 2746
rect 65834 2694 65846 2746
rect 65846 2694 65876 2746
rect 65900 2694 65910 2746
rect 65910 2694 65956 2746
rect 65660 2692 65716 2694
rect 65740 2692 65796 2694
rect 65820 2692 65876 2694
rect 65900 2692 65956 2694
rect 66994 2080 67050 2136
rect 67546 720 67602 776
<< metal3 >>
rect 67541 59258 67607 59261
rect 69200 59258 70000 59288
rect 67541 59256 70000 59258
rect 67541 59200 67546 59256
rect 67602 59200 70000 59256
rect 67541 59198 70000 59200
rect 67541 59195 67607 59198
rect 69200 59168 70000 59198
rect 66989 57898 67055 57901
rect 69200 57898 70000 57928
rect 66989 57896 70000 57898
rect 66989 57840 66994 57896
rect 67050 57840 70000 57896
rect 66989 57838 70000 57840
rect 66989 57835 67055 57838
rect 69200 57808 70000 57838
rect 19570 57696 19886 57697
rect 0 57536 800 57656
rect 19570 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19886 57696
rect 19570 57631 19886 57632
rect 50290 57696 50606 57697
rect 50290 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50606 57696
rect 50290 57631 50606 57632
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 34930 57087 35246 57088
rect 65650 57152 65966 57153
rect 65650 57088 65656 57152
rect 65720 57088 65736 57152
rect 65800 57088 65816 57152
rect 65880 57088 65896 57152
rect 65960 57088 65966 57152
rect 65650 57087 65966 57088
rect 19570 56608 19886 56609
rect 19570 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19886 56608
rect 19570 56543 19886 56544
rect 50290 56608 50606 56609
rect 50290 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50606 56608
rect 50290 56543 50606 56544
rect 68093 56538 68159 56541
rect 69200 56538 70000 56568
rect 68093 56536 70000 56538
rect 68093 56480 68098 56536
rect 68154 56480 70000 56536
rect 68093 56478 70000 56480
rect 68093 56475 68159 56478
rect 69200 56448 70000 56478
rect 0 56040 800 56160
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 34930 55999 35246 56000
rect 65650 56064 65966 56065
rect 65650 56000 65656 56064
rect 65720 56000 65736 56064
rect 65800 56000 65816 56064
rect 65880 56000 65896 56064
rect 65960 56000 65966 56064
rect 65650 55999 65966 56000
rect 19570 55520 19886 55521
rect 19570 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19886 55520
rect 19570 55455 19886 55456
rect 50290 55520 50606 55521
rect 50290 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50606 55520
rect 50290 55455 50606 55456
rect 67633 55178 67699 55181
rect 69200 55178 70000 55208
rect 67633 55176 70000 55178
rect 67633 55120 67638 55176
rect 67694 55120 70000 55176
rect 67633 55118 70000 55120
rect 67633 55115 67699 55118
rect 69200 55088 70000 55118
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 34930 54911 35246 54912
rect 65650 54976 65966 54977
rect 65650 54912 65656 54976
rect 65720 54912 65736 54976
rect 65800 54912 65816 54976
rect 65880 54912 65896 54976
rect 65960 54912 65966 54976
rect 65650 54911 65966 54912
rect 0 54544 800 54664
rect 19570 54432 19886 54433
rect 19570 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19886 54432
rect 19570 54367 19886 54368
rect 50290 54432 50606 54433
rect 50290 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50606 54432
rect 50290 54367 50606 54368
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 34930 53823 35246 53824
rect 65650 53888 65966 53889
rect 65650 53824 65656 53888
rect 65720 53824 65736 53888
rect 65800 53824 65816 53888
rect 65880 53824 65896 53888
rect 65960 53824 65966 53888
rect 65650 53823 65966 53824
rect 67541 53818 67607 53821
rect 69200 53818 70000 53848
rect 67541 53816 70000 53818
rect 67541 53760 67546 53816
rect 67602 53760 70000 53816
rect 67541 53758 70000 53760
rect 67541 53755 67607 53758
rect 69200 53728 70000 53758
rect 19570 53344 19886 53345
rect 19570 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19886 53344
rect 19570 53279 19886 53280
rect 50290 53344 50606 53345
rect 50290 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50606 53344
rect 50290 53279 50606 53280
rect 0 53048 800 53168
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 34930 52735 35246 52736
rect 65650 52800 65966 52801
rect 65650 52736 65656 52800
rect 65720 52736 65736 52800
rect 65800 52736 65816 52800
rect 65880 52736 65896 52800
rect 65960 52736 65966 52800
rect 65650 52735 65966 52736
rect 68093 52458 68159 52461
rect 69200 52458 70000 52488
rect 68093 52456 70000 52458
rect 68093 52400 68098 52456
rect 68154 52400 70000 52456
rect 68093 52398 70000 52400
rect 68093 52395 68159 52398
rect 69200 52368 70000 52398
rect 19570 52256 19886 52257
rect 19570 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19886 52256
rect 19570 52191 19886 52192
rect 50290 52256 50606 52257
rect 50290 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50606 52256
rect 50290 52191 50606 52192
rect 4210 51712 4526 51713
rect 0 51552 800 51672
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 34930 51647 35246 51648
rect 65650 51712 65966 51713
rect 65650 51648 65656 51712
rect 65720 51648 65736 51712
rect 65800 51648 65816 51712
rect 65880 51648 65896 51712
rect 65960 51648 65966 51712
rect 65650 51647 65966 51648
rect 19570 51168 19886 51169
rect 19570 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19886 51168
rect 19570 51103 19886 51104
rect 50290 51168 50606 51169
rect 50290 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50606 51168
rect 50290 51103 50606 51104
rect 68093 51098 68159 51101
rect 69200 51098 70000 51128
rect 68093 51096 70000 51098
rect 68093 51040 68098 51096
rect 68154 51040 70000 51096
rect 68093 51038 70000 51040
rect 68093 51035 68159 51038
rect 69200 51008 70000 51038
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 34930 50559 35246 50560
rect 65650 50624 65966 50625
rect 65650 50560 65656 50624
rect 65720 50560 65736 50624
rect 65800 50560 65816 50624
rect 65880 50560 65896 50624
rect 65960 50560 65966 50624
rect 65650 50559 65966 50560
rect 0 50056 800 50176
rect 19570 50080 19886 50081
rect 19570 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19886 50080
rect 19570 50015 19886 50016
rect 50290 50080 50606 50081
rect 50290 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50606 50080
rect 50290 50015 50606 50016
rect 67633 49738 67699 49741
rect 69200 49738 70000 49768
rect 67633 49736 70000 49738
rect 67633 49680 67638 49736
rect 67694 49680 70000 49736
rect 67633 49678 70000 49680
rect 67633 49675 67699 49678
rect 69200 49648 70000 49678
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 34930 49471 35246 49472
rect 65650 49536 65966 49537
rect 65650 49472 65656 49536
rect 65720 49472 65736 49536
rect 65800 49472 65816 49536
rect 65880 49472 65896 49536
rect 65960 49472 65966 49536
rect 65650 49471 65966 49472
rect 19570 48992 19886 48993
rect 19570 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19886 48992
rect 19570 48927 19886 48928
rect 50290 48992 50606 48993
rect 50290 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50606 48992
rect 50290 48927 50606 48928
rect 0 48560 800 48680
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 34930 48383 35246 48384
rect 65650 48448 65966 48449
rect 65650 48384 65656 48448
rect 65720 48384 65736 48448
rect 65800 48384 65816 48448
rect 65880 48384 65896 48448
rect 65960 48384 65966 48448
rect 65650 48383 65966 48384
rect 67633 48378 67699 48381
rect 69200 48378 70000 48408
rect 67633 48376 70000 48378
rect 67633 48320 67638 48376
rect 67694 48320 70000 48376
rect 67633 48318 70000 48320
rect 67633 48315 67699 48318
rect 69200 48288 70000 48318
rect 19570 47904 19886 47905
rect 19570 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19886 47904
rect 19570 47839 19886 47840
rect 50290 47904 50606 47905
rect 50290 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50606 47904
rect 50290 47839 50606 47840
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 65650 47360 65966 47361
rect 65650 47296 65656 47360
rect 65720 47296 65736 47360
rect 65800 47296 65816 47360
rect 65880 47296 65896 47360
rect 65960 47296 65966 47360
rect 65650 47295 65966 47296
rect 0 47064 800 47184
rect 68093 47018 68159 47021
rect 69200 47018 70000 47048
rect 68093 47016 70000 47018
rect 68093 46960 68098 47016
rect 68154 46960 70000 47016
rect 68093 46958 70000 46960
rect 68093 46955 68159 46958
rect 69200 46928 70000 46958
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 50290 46816 50606 46817
rect 50290 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50606 46816
rect 50290 46751 50606 46752
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 65650 46272 65966 46273
rect 65650 46208 65656 46272
rect 65720 46208 65736 46272
rect 65800 46208 65816 46272
rect 65880 46208 65896 46272
rect 65960 46208 65966 46272
rect 65650 46207 65966 46208
rect 19570 45728 19886 45729
rect 0 45568 800 45688
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 50290 45728 50606 45729
rect 50290 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50606 45728
rect 50290 45663 50606 45664
rect 68093 45658 68159 45661
rect 69200 45658 70000 45688
rect 68093 45656 70000 45658
rect 68093 45600 68098 45656
rect 68154 45600 70000 45656
rect 68093 45598 70000 45600
rect 68093 45595 68159 45598
rect 69200 45568 70000 45598
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 65650 45184 65966 45185
rect 65650 45120 65656 45184
rect 65720 45120 65736 45184
rect 65800 45120 65816 45184
rect 65880 45120 65896 45184
rect 65960 45120 65966 45184
rect 65650 45119 65966 45120
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 50290 44640 50606 44641
rect 50290 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50606 44640
rect 50290 44575 50606 44576
rect 67633 44298 67699 44301
rect 69200 44298 70000 44328
rect 67633 44296 70000 44298
rect 67633 44240 67638 44296
rect 67694 44240 70000 44296
rect 67633 44238 70000 44240
rect 67633 44235 67699 44238
rect 69200 44208 70000 44238
rect 0 44072 800 44192
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 65650 44096 65966 44097
rect 65650 44032 65656 44096
rect 65720 44032 65736 44096
rect 65800 44032 65816 44096
rect 65880 44032 65896 44096
rect 65960 44032 65966 44096
rect 65650 44031 65966 44032
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 50290 43552 50606 43553
rect 50290 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50606 43552
rect 50290 43487 50606 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 65650 43008 65966 43009
rect 65650 42944 65656 43008
rect 65720 42944 65736 43008
rect 65800 42944 65816 43008
rect 65880 42944 65896 43008
rect 65960 42944 65966 43008
rect 65650 42943 65966 42944
rect 67633 42938 67699 42941
rect 69200 42938 70000 42968
rect 67633 42936 70000 42938
rect 67633 42880 67638 42936
rect 67694 42880 70000 42936
rect 67633 42878 70000 42880
rect 67633 42875 67699 42878
rect 69200 42848 70000 42878
rect 0 42576 800 42696
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 50290 42464 50606 42465
rect 50290 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50606 42464
rect 50290 42399 50606 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 65650 41920 65966 41921
rect 65650 41856 65656 41920
rect 65720 41856 65736 41920
rect 65800 41856 65816 41920
rect 65880 41856 65896 41920
rect 65960 41856 65966 41920
rect 65650 41855 65966 41856
rect 68093 41578 68159 41581
rect 69200 41578 70000 41608
rect 68093 41576 70000 41578
rect 68093 41520 68098 41576
rect 68154 41520 70000 41576
rect 68093 41518 70000 41520
rect 68093 41515 68159 41518
rect 69200 41488 70000 41518
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 50290 41376 50606 41377
rect 50290 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50606 41376
rect 50290 41311 50606 41312
rect 0 41080 800 41200
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 65650 40832 65966 40833
rect 65650 40768 65656 40832
rect 65720 40768 65736 40832
rect 65800 40768 65816 40832
rect 65880 40768 65896 40832
rect 65960 40768 65966 40832
rect 65650 40767 65966 40768
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 50290 40288 50606 40289
rect 50290 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50606 40288
rect 50290 40223 50606 40224
rect 68093 40218 68159 40221
rect 69200 40218 70000 40248
rect 68093 40216 70000 40218
rect 68093 40160 68098 40216
rect 68154 40160 70000 40216
rect 68093 40158 70000 40160
rect 68093 40155 68159 40158
rect 69200 40128 70000 40158
rect 4210 39744 4526 39745
rect 0 39584 800 39704
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 65650 39744 65966 39745
rect 65650 39680 65656 39744
rect 65720 39680 65736 39744
rect 65800 39680 65816 39744
rect 65880 39680 65896 39744
rect 65960 39680 65966 39744
rect 65650 39679 65966 39680
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 50290 39135 50606 39136
rect 67633 38858 67699 38861
rect 69200 38858 70000 38888
rect 67633 38856 70000 38858
rect 67633 38800 67638 38856
rect 67694 38800 70000 38856
rect 67633 38798 70000 38800
rect 67633 38795 67699 38798
rect 69200 38768 70000 38798
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 65650 38656 65966 38657
rect 65650 38592 65656 38656
rect 65720 38592 65736 38656
rect 65800 38592 65816 38656
rect 65880 38592 65896 38656
rect 65960 38592 65966 38656
rect 65650 38591 65966 38592
rect 0 38088 800 38208
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 50290 38047 50606 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 65650 37568 65966 37569
rect 65650 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65966 37568
rect 65650 37503 65966 37504
rect 67633 37498 67699 37501
rect 69200 37498 70000 37528
rect 67633 37496 70000 37498
rect 67633 37440 67638 37496
rect 67694 37440 70000 37496
rect 67633 37438 70000 37440
rect 67633 37435 67699 37438
rect 69200 37408 70000 37438
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 50290 36959 50606 36960
rect 0 36592 800 36712
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 65650 36480 65966 36481
rect 65650 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65966 36480
rect 65650 36415 65966 36416
rect 68093 36138 68159 36141
rect 69200 36138 70000 36168
rect 68093 36136 70000 36138
rect 68093 36080 68098 36136
rect 68154 36080 70000 36136
rect 68093 36078 70000 36080
rect 68093 36075 68159 36078
rect 69200 36048 70000 36078
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 50290 35871 50606 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 65650 35392 65966 35393
rect 65650 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65966 35392
rect 65650 35327 65966 35328
rect 0 35096 800 35216
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 50290 34783 50606 34784
rect 68093 34778 68159 34781
rect 69200 34778 70000 34808
rect 68093 34776 70000 34778
rect 68093 34720 68098 34776
rect 68154 34720 70000 34776
rect 68093 34718 70000 34720
rect 68093 34715 68159 34718
rect 69200 34688 70000 34718
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 65650 34304 65966 34305
rect 65650 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65966 34304
rect 65650 34239 65966 34240
rect 19570 33760 19886 33761
rect 0 33600 800 33720
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 50290 33695 50606 33696
rect 67633 33418 67699 33421
rect 69200 33418 70000 33448
rect 67633 33416 70000 33418
rect 67633 33360 67638 33416
rect 67694 33360 70000 33416
rect 67633 33358 70000 33360
rect 67633 33355 67699 33358
rect 69200 33328 70000 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 65650 33216 65966 33217
rect 65650 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65966 33216
rect 65650 33151 65966 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 50290 32607 50606 32608
rect 0 32104 800 32224
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 65650 32128 65966 32129
rect 65650 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65966 32128
rect 65650 32063 65966 32064
rect 67633 32058 67699 32061
rect 69200 32058 70000 32088
rect 67633 32056 70000 32058
rect 67633 32000 67638 32056
rect 67694 32000 70000 32056
rect 67633 31998 70000 32000
rect 67633 31995 67699 31998
rect 69200 31968 70000 31998
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 50290 31519 50606 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 65650 31040 65966 31041
rect 65650 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65966 31040
rect 65650 30975 65966 30976
rect 0 30608 800 30728
rect 68093 30698 68159 30701
rect 69200 30698 70000 30728
rect 68093 30696 70000 30698
rect 68093 30640 68098 30696
rect 68154 30640 70000 30696
rect 68093 30638 70000 30640
rect 68093 30635 68159 30638
rect 69200 30608 70000 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 50290 30431 50606 30432
rect 5809 30154 5875 30157
rect 17309 30154 17375 30157
rect 5809 30152 17375 30154
rect 5809 30096 5814 30152
rect 5870 30096 17314 30152
rect 17370 30096 17375 30152
rect 5809 30094 17375 30096
rect 5809 30091 5875 30094
rect 17309 30091 17375 30094
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 65650 29952 65966 29953
rect 65650 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65966 29952
rect 65650 29887 65966 29888
rect 7281 29610 7347 29613
rect 8109 29610 8175 29613
rect 19609 29610 19675 29613
rect 7281 29608 19675 29610
rect 7281 29552 7286 29608
rect 7342 29552 8114 29608
rect 8170 29552 19614 29608
rect 19670 29552 19675 29608
rect 7281 29550 19675 29552
rect 7281 29547 7347 29550
rect 8109 29547 8175 29550
rect 19609 29547 19675 29550
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 50290 29343 50606 29344
rect 68093 29338 68159 29341
rect 69200 29338 70000 29368
rect 68093 29336 70000 29338
rect 68093 29280 68098 29336
rect 68154 29280 70000 29336
rect 68093 29278 70000 29280
rect 68093 29275 68159 29278
rect 69200 29248 70000 29278
rect 0 29112 800 29232
rect 5441 29066 5507 29069
rect 17125 29066 17191 29069
rect 5441 29064 17191 29066
rect 5441 29008 5446 29064
rect 5502 29008 17130 29064
rect 17186 29008 17191 29064
rect 5441 29006 17191 29008
rect 5441 29003 5507 29006
rect 17125 29003 17191 29006
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 65650 28864 65966 28865
rect 65650 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65966 28864
rect 65650 28799 65966 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 50290 28255 50606 28256
rect 67633 27978 67699 27981
rect 69200 27978 70000 28008
rect 67633 27976 70000 27978
rect 67633 27920 67638 27976
rect 67694 27920 70000 27976
rect 67633 27918 70000 27920
rect 67633 27915 67699 27918
rect 69200 27888 70000 27918
rect 4210 27776 4526 27777
rect 0 27616 800 27736
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 65650 27776 65966 27777
rect 65650 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65966 27776
rect 65650 27711 65966 27712
rect 23197 27434 23263 27437
rect 24209 27434 24275 27437
rect 23197 27432 24275 27434
rect 23197 27376 23202 27432
rect 23258 27376 24214 27432
rect 24270 27376 24275 27432
rect 23197 27374 24275 27376
rect 23197 27371 23263 27374
rect 24209 27371 24275 27374
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 50290 27167 50606 27168
rect 9581 26890 9647 26893
rect 17125 26890 17191 26893
rect 9581 26888 17191 26890
rect 9581 26832 9586 26888
rect 9642 26832 17130 26888
rect 17186 26832 17191 26888
rect 9581 26830 17191 26832
rect 9581 26827 9647 26830
rect 17125 26827 17191 26830
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 65650 26688 65966 26689
rect 65650 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65966 26688
rect 65650 26623 65966 26624
rect 67633 26618 67699 26621
rect 69200 26618 70000 26648
rect 67633 26616 70000 26618
rect 67633 26560 67638 26616
rect 67694 26560 70000 26616
rect 67633 26558 70000 26560
rect 67633 26555 67699 26558
rect 69200 26528 70000 26558
rect 17401 26346 17467 26349
rect 17534 26346 17540 26348
rect 17401 26344 17540 26346
rect 17401 26288 17406 26344
rect 17462 26288 17540 26344
rect 17401 26286 17540 26288
rect 17401 26283 17467 26286
rect 17534 26284 17540 26286
rect 17604 26284 17610 26348
rect 0 26120 800 26240
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 50290 26079 50606 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 65650 25600 65966 25601
rect 65650 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65966 25600
rect 65650 25535 65966 25536
rect 12985 25258 13051 25261
rect 17401 25258 17467 25261
rect 12985 25256 17467 25258
rect 12985 25200 12990 25256
rect 13046 25200 17406 25256
rect 17462 25200 17467 25256
rect 12985 25198 17467 25200
rect 12985 25195 13051 25198
rect 17401 25195 17467 25198
rect 68093 25258 68159 25261
rect 69200 25258 70000 25288
rect 68093 25256 70000 25258
rect 68093 25200 68098 25256
rect 68154 25200 70000 25256
rect 68093 25198 70000 25200
rect 68093 25195 68159 25198
rect 69200 25168 70000 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 50290 24991 50606 24992
rect 17677 24988 17743 24989
rect 17677 24984 17724 24988
rect 17788 24986 17794 24988
rect 17677 24928 17682 24984
rect 17677 24924 17724 24928
rect 17788 24926 17834 24986
rect 17788 24924 17794 24926
rect 17677 24923 17743 24924
rect 0 24624 800 24744
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 65650 24512 65966 24513
rect 65650 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65966 24512
rect 65650 24447 65966 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 50290 23903 50606 23904
rect 68093 23898 68159 23901
rect 69200 23898 70000 23928
rect 68093 23896 70000 23898
rect 68093 23840 68098 23896
rect 68154 23840 70000 23896
rect 68093 23838 70000 23840
rect 68093 23835 68159 23838
rect 69200 23808 70000 23838
rect 17309 23762 17375 23765
rect 18229 23762 18295 23765
rect 17309 23760 18295 23762
rect 17309 23704 17314 23760
rect 17370 23704 18234 23760
rect 18290 23704 18295 23760
rect 17309 23702 18295 23704
rect 17309 23699 17375 23702
rect 18229 23699 18295 23702
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 65650 23424 65966 23425
rect 65650 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65966 23424
rect 65650 23359 65966 23360
rect 19333 23354 19399 23357
rect 26141 23354 26207 23357
rect 19333 23352 26207 23354
rect 19333 23296 19338 23352
rect 19394 23296 26146 23352
rect 26202 23296 26207 23352
rect 19333 23294 26207 23296
rect 19333 23291 19399 23294
rect 26141 23291 26207 23294
rect 0 23128 800 23248
rect 5165 23082 5231 23085
rect 15377 23082 15443 23085
rect 5165 23080 15443 23082
rect 5165 23024 5170 23080
rect 5226 23024 15382 23080
rect 15438 23024 15443 23080
rect 5165 23022 15443 23024
rect 5165 23019 5231 23022
rect 15377 23019 15443 23022
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 50290 22815 50606 22816
rect 4613 22538 4679 22541
rect 13905 22538 13971 22541
rect 4613 22536 13971 22538
rect 4613 22480 4618 22536
rect 4674 22480 13910 22536
rect 13966 22480 13971 22536
rect 4613 22478 13971 22480
rect 4613 22475 4679 22478
rect 13905 22475 13971 22478
rect 67633 22538 67699 22541
rect 69200 22538 70000 22568
rect 67633 22536 70000 22538
rect 67633 22480 67638 22536
rect 67694 22480 70000 22536
rect 67633 22478 70000 22480
rect 67633 22475 67699 22478
rect 69200 22448 70000 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 65650 22336 65966 22337
rect 65650 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65966 22336
rect 65650 22271 65966 22272
rect 15285 22268 15351 22269
rect 15285 22264 15332 22268
rect 15396 22266 15402 22268
rect 15285 22208 15290 22264
rect 15285 22204 15332 22208
rect 15396 22206 15442 22266
rect 15396 22204 15402 22206
rect 15285 22203 15351 22204
rect 5073 22130 5139 22133
rect 11053 22130 11119 22133
rect 5073 22128 11119 22130
rect 5073 22072 5078 22128
rect 5134 22072 11058 22128
rect 11114 22072 11119 22128
rect 5073 22070 11119 22072
rect 5073 22067 5139 22070
rect 11053 22067 11119 22070
rect 21909 21994 21975 21997
rect 30557 21994 30623 21997
rect 31477 21994 31543 21997
rect 21909 21992 31543 21994
rect 21909 21936 21914 21992
rect 21970 21936 30562 21992
rect 30618 21936 31482 21992
rect 31538 21936 31543 21992
rect 21909 21934 31543 21936
rect 21909 21931 21975 21934
rect 30557 21931 30623 21934
rect 31477 21931 31543 21934
rect 19570 21792 19886 21793
rect 0 21632 800 21752
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 50290 21727 50606 21728
rect 10961 21450 11027 21453
rect 23473 21450 23539 21453
rect 10961 21448 23539 21450
rect 10961 21392 10966 21448
rect 11022 21392 23478 21448
rect 23534 21392 23539 21448
rect 10961 21390 23539 21392
rect 10961 21387 11027 21390
rect 23473 21387 23539 21390
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 65650 21248 65966 21249
rect 65650 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65966 21248
rect 65650 21183 65966 21184
rect 67633 21178 67699 21181
rect 69200 21178 70000 21208
rect 67633 21176 70000 21178
rect 67633 21120 67638 21176
rect 67694 21120 70000 21176
rect 67633 21118 70000 21120
rect 67633 21115 67699 21118
rect 69200 21088 70000 21118
rect 22737 20906 22803 20909
rect 25405 20906 25471 20909
rect 22737 20904 25471 20906
rect 22737 20848 22742 20904
rect 22798 20848 25410 20904
rect 25466 20848 25471 20904
rect 22737 20846 25471 20848
rect 22737 20843 22803 20846
rect 25405 20843 25471 20846
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 50290 20639 50606 20640
rect 25681 20634 25747 20637
rect 23798 20632 25747 20634
rect 23798 20576 25686 20632
rect 25742 20576 25747 20632
rect 23798 20574 25747 20576
rect 9029 20498 9095 20501
rect 23565 20498 23631 20501
rect 9029 20496 23631 20498
rect 9029 20440 9034 20496
rect 9090 20440 23570 20496
rect 23626 20440 23631 20496
rect 9029 20438 23631 20440
rect 9029 20435 9095 20438
rect 23565 20435 23631 20438
rect 1945 20362 2011 20365
rect 4153 20362 4219 20365
rect 1945 20360 4219 20362
rect 1945 20304 1950 20360
rect 2006 20304 4158 20360
rect 4214 20304 4219 20360
rect 1945 20302 4219 20304
rect 1945 20299 2011 20302
rect 4153 20299 4219 20302
rect 19793 20362 19859 20365
rect 23798 20362 23858 20574
rect 25681 20571 25747 20574
rect 19793 20360 23858 20362
rect 19793 20304 19798 20360
rect 19854 20304 23858 20360
rect 19793 20302 23858 20304
rect 19793 20299 19859 20302
rect 0 20136 800 20256
rect 13445 20226 13511 20229
rect 18965 20226 19031 20229
rect 21817 20226 21883 20229
rect 13445 20224 21883 20226
rect 13445 20168 13450 20224
rect 13506 20168 18970 20224
rect 19026 20168 21822 20224
rect 21878 20168 21883 20224
rect 13445 20166 21883 20168
rect 13445 20163 13511 20166
rect 18965 20163 19031 20166
rect 21817 20163 21883 20166
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 65650 20160 65966 20161
rect 65650 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65966 20160
rect 65650 20095 65966 20096
rect 15837 20090 15903 20093
rect 19517 20090 19583 20093
rect 15837 20088 19583 20090
rect 15837 20032 15842 20088
rect 15898 20032 19522 20088
rect 19578 20032 19583 20088
rect 15837 20030 19583 20032
rect 15837 20027 15903 20030
rect 19517 20027 19583 20030
rect 68093 19818 68159 19821
rect 69200 19818 70000 19848
rect 68093 19816 70000 19818
rect 68093 19760 68098 19816
rect 68154 19760 70000 19816
rect 68093 19758 70000 19760
rect 68093 19755 68159 19758
rect 69200 19728 70000 19758
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 50290 19551 50606 19552
rect 2129 19410 2195 19413
rect 4797 19410 4863 19413
rect 2129 19408 4863 19410
rect 2129 19352 2134 19408
rect 2190 19352 4802 19408
rect 4858 19352 4863 19408
rect 2129 19350 4863 19352
rect 2129 19347 2195 19350
rect 4797 19347 4863 19350
rect 8477 19410 8543 19413
rect 9213 19410 9279 19413
rect 8477 19408 9279 19410
rect 8477 19352 8482 19408
rect 8538 19352 9218 19408
rect 9274 19352 9279 19408
rect 8477 19350 9279 19352
rect 8477 19347 8543 19350
rect 9213 19347 9279 19350
rect 18965 19410 19031 19413
rect 22553 19410 22619 19413
rect 18965 19408 22619 19410
rect 18965 19352 18970 19408
rect 19026 19352 22558 19408
rect 22614 19352 22619 19408
rect 18965 19350 22619 19352
rect 18965 19347 19031 19350
rect 22553 19347 22619 19350
rect 21173 19274 21239 19277
rect 30833 19274 30899 19277
rect 21173 19272 30899 19274
rect 21173 19216 21178 19272
rect 21234 19216 30838 19272
rect 30894 19216 30899 19272
rect 21173 19214 30899 19216
rect 21173 19211 21239 19214
rect 30833 19211 30899 19214
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 65650 19072 65966 19073
rect 65650 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65966 19072
rect 65650 19007 65966 19008
rect 0 18640 800 18760
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 50290 18463 50606 18464
rect 20989 18458 21055 18461
rect 26325 18458 26391 18461
rect 20118 18456 26391 18458
rect 20118 18400 20994 18456
rect 21050 18400 26330 18456
rect 26386 18400 26391 18456
rect 20118 18398 26391 18400
rect 17125 18322 17191 18325
rect 20118 18322 20178 18398
rect 20989 18395 21055 18398
rect 26325 18395 26391 18398
rect 68093 18458 68159 18461
rect 69200 18458 70000 18488
rect 68093 18456 70000 18458
rect 68093 18400 68098 18456
rect 68154 18400 70000 18456
rect 68093 18398 70000 18400
rect 68093 18395 68159 18398
rect 69200 18368 70000 18398
rect 17125 18320 20178 18322
rect 17125 18264 17130 18320
rect 17186 18264 20178 18320
rect 17125 18262 20178 18264
rect 21081 18322 21147 18325
rect 33317 18322 33383 18325
rect 21081 18320 33383 18322
rect 21081 18264 21086 18320
rect 21142 18264 33322 18320
rect 33378 18264 33383 18320
rect 21081 18262 33383 18264
rect 17125 18259 17191 18262
rect 21081 18259 21147 18262
rect 33317 18259 33383 18262
rect 17309 18186 17375 18189
rect 31017 18186 31083 18189
rect 17309 18184 31083 18186
rect 17309 18128 17314 18184
rect 17370 18128 31022 18184
rect 31078 18128 31083 18184
rect 17309 18126 31083 18128
rect 17309 18123 17375 18126
rect 31017 18123 31083 18126
rect 20529 18050 20595 18053
rect 26509 18050 26575 18053
rect 20529 18048 26575 18050
rect 20529 17992 20534 18048
rect 20590 17992 26514 18048
rect 26570 17992 26575 18048
rect 20529 17990 26575 17992
rect 20529 17987 20595 17990
rect 26509 17987 26575 17990
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 65650 17984 65966 17985
rect 65650 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65966 17984
rect 65650 17919 65966 17920
rect 11053 17642 11119 17645
rect 21357 17642 21423 17645
rect 11053 17640 21423 17642
rect 11053 17584 11058 17640
rect 11114 17584 21362 17640
rect 21418 17584 21423 17640
rect 11053 17582 21423 17584
rect 11053 17579 11119 17582
rect 21357 17579 21423 17582
rect 38009 17642 38075 17645
rect 39297 17642 39363 17645
rect 38009 17640 39363 17642
rect 38009 17584 38014 17640
rect 38070 17584 39302 17640
rect 39358 17584 39363 17640
rect 38009 17582 39363 17584
rect 38009 17579 38075 17582
rect 39297 17579 39363 17582
rect 29637 17506 29703 17509
rect 36629 17506 36695 17509
rect 29637 17504 36695 17506
rect 29637 17448 29642 17504
rect 29698 17448 36634 17504
rect 36690 17448 36695 17504
rect 29637 17446 36695 17448
rect 29637 17443 29703 17446
rect 36629 17443 36695 17446
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 50290 17375 50606 17376
rect 0 17144 800 17264
rect 1853 17234 1919 17237
rect 6269 17234 6335 17237
rect 1853 17232 6335 17234
rect 1853 17176 1858 17232
rect 1914 17176 6274 17232
rect 6330 17176 6335 17232
rect 1853 17174 6335 17176
rect 1853 17171 1919 17174
rect 6269 17171 6335 17174
rect 15837 17234 15903 17237
rect 23105 17234 23171 17237
rect 15837 17232 23171 17234
rect 15837 17176 15842 17232
rect 15898 17176 23110 17232
rect 23166 17176 23171 17232
rect 15837 17174 23171 17176
rect 15837 17171 15903 17174
rect 23105 17171 23171 17174
rect 26509 17234 26575 17237
rect 28625 17234 28691 17237
rect 26509 17232 28691 17234
rect 26509 17176 26514 17232
rect 26570 17176 28630 17232
rect 28686 17176 28691 17232
rect 26509 17174 28691 17176
rect 26509 17171 26575 17174
rect 28625 17171 28691 17174
rect 67633 17098 67699 17101
rect 69200 17098 70000 17128
rect 67633 17096 70000 17098
rect 67633 17040 67638 17096
rect 67694 17040 70000 17096
rect 67633 17038 70000 17040
rect 67633 17035 67699 17038
rect 69200 17008 70000 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 65650 16896 65966 16897
rect 65650 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65966 16896
rect 65650 16831 65966 16832
rect 23197 16690 23263 16693
rect 23197 16688 28642 16690
rect 23197 16632 23202 16688
rect 23258 16632 28642 16688
rect 23197 16630 28642 16632
rect 23197 16627 23263 16630
rect 28582 16557 28642 16630
rect 7005 16554 7071 16557
rect 27245 16554 27311 16557
rect 7005 16552 27311 16554
rect 7005 16496 7010 16552
rect 7066 16496 27250 16552
rect 27306 16496 27311 16552
rect 7005 16494 27311 16496
rect 28582 16552 28691 16557
rect 28582 16496 28630 16552
rect 28686 16496 28691 16552
rect 28582 16494 28691 16496
rect 7005 16491 7071 16494
rect 27245 16491 27311 16494
rect 28625 16491 28691 16494
rect 31109 16554 31175 16557
rect 37917 16554 37983 16557
rect 31109 16552 37983 16554
rect 31109 16496 31114 16552
rect 31170 16496 37922 16552
rect 37978 16496 37983 16552
rect 31109 16494 37983 16496
rect 31109 16491 31175 16494
rect 37917 16491 37983 16494
rect 21817 16418 21883 16421
rect 30373 16418 30439 16421
rect 21817 16416 30439 16418
rect 21817 16360 21822 16416
rect 21878 16360 30378 16416
rect 30434 16360 30439 16416
rect 21817 16358 30439 16360
rect 21817 16355 21883 16358
rect 30373 16355 30439 16358
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 50290 16287 50606 16288
rect 26325 16282 26391 16285
rect 33685 16282 33751 16285
rect 26325 16280 33751 16282
rect 26325 16224 26330 16280
rect 26386 16224 33690 16280
rect 33746 16224 33751 16280
rect 26325 16222 33751 16224
rect 26325 16219 26391 16222
rect 33685 16219 33751 16222
rect 5441 16010 5507 16013
rect 22277 16010 22343 16013
rect 5441 16008 22343 16010
rect 5441 15952 5446 16008
rect 5502 15952 22282 16008
rect 22338 15952 22343 16008
rect 5441 15950 22343 15952
rect 5441 15947 5507 15950
rect 22277 15947 22343 15950
rect 4210 15808 4526 15809
rect 0 15648 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 65650 15808 65966 15809
rect 65650 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65966 15808
rect 65650 15743 65966 15744
rect 19057 15738 19123 15741
rect 24853 15738 24919 15741
rect 19057 15736 24919 15738
rect 19057 15680 19062 15736
rect 19118 15680 24858 15736
rect 24914 15680 24919 15736
rect 19057 15678 24919 15680
rect 19057 15675 19123 15678
rect 24853 15675 24919 15678
rect 67633 15738 67699 15741
rect 69200 15738 70000 15768
rect 67633 15736 70000 15738
rect 67633 15680 67638 15736
rect 67694 15680 70000 15736
rect 67633 15678 70000 15680
rect 67633 15675 67699 15678
rect 69200 15648 70000 15678
rect 12157 15466 12223 15469
rect 23197 15466 23263 15469
rect 12157 15464 23263 15466
rect 12157 15408 12162 15464
rect 12218 15408 23202 15464
rect 23258 15408 23263 15464
rect 12157 15406 23263 15408
rect 12157 15403 12223 15406
rect 23197 15403 23263 15406
rect 35985 15330 36051 15333
rect 38929 15330 38995 15333
rect 35985 15328 38995 15330
rect 35985 15272 35990 15328
rect 36046 15272 38934 15328
rect 38990 15272 38995 15328
rect 35985 15270 38995 15272
rect 35985 15267 36051 15270
rect 38929 15267 38995 15270
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 50290 15199 50606 15200
rect 22277 15058 22343 15061
rect 35985 15058 36051 15061
rect 22277 15056 36051 15058
rect 22277 15000 22282 15056
rect 22338 15000 35990 15056
rect 36046 15000 36051 15056
rect 22277 14998 36051 15000
rect 22277 14995 22343 14998
rect 35985 14995 36051 14998
rect 5625 14922 5691 14925
rect 22001 14922 22067 14925
rect 5625 14920 22067 14922
rect 5625 14864 5630 14920
rect 5686 14864 22006 14920
rect 22062 14864 22067 14920
rect 5625 14862 22067 14864
rect 5625 14859 5691 14862
rect 22001 14859 22067 14862
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 65650 14720 65966 14721
rect 65650 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65966 14720
rect 65650 14655 65966 14656
rect 68093 14378 68159 14381
rect 69200 14378 70000 14408
rect 68093 14376 70000 14378
rect 68093 14320 68098 14376
rect 68154 14320 70000 14376
rect 68093 14318 70000 14320
rect 68093 14315 68159 14318
rect 69200 14288 70000 14318
rect 0 14152 800 14272
rect 27705 14242 27771 14245
rect 32949 14242 33015 14245
rect 27705 14240 33015 14242
rect 27705 14184 27710 14240
rect 27766 14184 32954 14240
rect 33010 14184 33015 14240
rect 27705 14182 33015 14184
rect 27705 14179 27771 14182
rect 32949 14179 33015 14182
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 50290 14111 50606 14112
rect 24945 13970 25011 13973
rect 34697 13970 34763 13973
rect 24945 13968 34763 13970
rect 24945 13912 24950 13968
rect 25006 13912 34702 13968
rect 34758 13912 34763 13968
rect 24945 13910 34763 13912
rect 24945 13907 25011 13910
rect 34697 13907 34763 13910
rect 9949 13834 10015 13837
rect 16573 13834 16639 13837
rect 9949 13832 16639 13834
rect 9949 13776 9954 13832
rect 10010 13776 16578 13832
rect 16634 13776 16639 13832
rect 9949 13774 16639 13776
rect 9949 13771 10015 13774
rect 16573 13771 16639 13774
rect 15326 13636 15332 13700
rect 15396 13698 15402 13700
rect 16665 13698 16731 13701
rect 15396 13696 16731 13698
rect 15396 13640 16670 13696
rect 16726 13640 16731 13696
rect 15396 13638 16731 13640
rect 15396 13636 15402 13638
rect 16665 13635 16731 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 65650 13632 65966 13633
rect 65650 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65966 13632
rect 65650 13567 65966 13568
rect 17677 13562 17743 13565
rect 20713 13562 20779 13565
rect 17677 13560 20779 13562
rect 17677 13504 17682 13560
rect 17738 13504 20718 13560
rect 20774 13504 20779 13560
rect 17677 13502 20779 13504
rect 17677 13499 17743 13502
rect 20713 13499 20779 13502
rect 2497 13426 2563 13429
rect 7097 13426 7163 13429
rect 2497 13424 7163 13426
rect 2497 13368 2502 13424
rect 2558 13368 7102 13424
rect 7158 13368 7163 13424
rect 2497 13366 7163 13368
rect 2497 13363 2563 13366
rect 7097 13363 7163 13366
rect 16757 13426 16823 13429
rect 27889 13426 27955 13429
rect 16757 13424 27955 13426
rect 16757 13368 16762 13424
rect 16818 13368 27894 13424
rect 27950 13368 27955 13424
rect 16757 13366 27955 13368
rect 16757 13363 16823 13366
rect 27889 13363 27955 13366
rect 28717 13426 28783 13429
rect 33041 13426 33107 13429
rect 28717 13424 33107 13426
rect 28717 13368 28722 13424
rect 28778 13368 33046 13424
rect 33102 13368 33107 13424
rect 28717 13366 33107 13368
rect 28717 13363 28783 13366
rect 33041 13363 33107 13366
rect 12065 13290 12131 13293
rect 23565 13290 23631 13293
rect 12065 13288 23631 13290
rect 12065 13232 12070 13288
rect 12126 13232 23570 13288
rect 23626 13232 23631 13288
rect 12065 13230 23631 13232
rect 12065 13227 12131 13230
rect 23565 13227 23631 13230
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 50290 13023 50606 13024
rect 68093 13018 68159 13021
rect 69200 13018 70000 13048
rect 68093 13016 70000 13018
rect 68093 12960 68098 13016
rect 68154 12960 70000 13016
rect 68093 12958 70000 12960
rect 68093 12955 68159 12958
rect 69200 12928 70000 12958
rect 19793 12882 19859 12885
rect 20161 12882 20227 12885
rect 24669 12882 24735 12885
rect 19793 12880 24735 12882
rect 19793 12824 19798 12880
rect 19854 12824 20166 12880
rect 20222 12824 24674 12880
rect 24730 12824 24735 12880
rect 19793 12822 24735 12824
rect 19793 12819 19859 12822
rect 20161 12819 20227 12822
rect 24669 12819 24735 12822
rect 0 12656 800 12776
rect 12065 12746 12131 12749
rect 23473 12746 23539 12749
rect 12065 12744 23539 12746
rect 12065 12688 12070 12744
rect 12126 12688 23478 12744
rect 23534 12688 23539 12744
rect 12065 12686 23539 12688
rect 12065 12683 12131 12686
rect 23473 12683 23539 12686
rect 14181 12612 14247 12613
rect 14181 12610 14228 12612
rect 14136 12608 14228 12610
rect 14136 12552 14186 12608
rect 14136 12550 14228 12552
rect 14181 12548 14228 12550
rect 14292 12548 14298 12612
rect 14181 12547 14247 12548
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 65650 12544 65966 12545
rect 65650 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65966 12544
rect 65650 12479 65966 12480
rect 10777 12338 10843 12341
rect 27981 12338 28047 12341
rect 10777 12336 28047 12338
rect 10777 12280 10782 12336
rect 10838 12280 27986 12336
rect 28042 12280 28047 12336
rect 10777 12278 28047 12280
rect 10777 12275 10843 12278
rect 27981 12275 28047 12278
rect 7557 12202 7623 12205
rect 12433 12202 12499 12205
rect 7557 12200 12499 12202
rect 7557 12144 7562 12200
rect 7618 12144 12438 12200
rect 12494 12144 12499 12200
rect 7557 12142 12499 12144
rect 7557 12139 7623 12142
rect 12433 12139 12499 12142
rect 12617 12202 12683 12205
rect 16430 12202 16436 12204
rect 12617 12200 16436 12202
rect 12617 12144 12622 12200
rect 12678 12144 16436 12200
rect 12617 12142 16436 12144
rect 12617 12139 12683 12142
rect 16430 12140 16436 12142
rect 16500 12140 16506 12204
rect 17493 12202 17559 12205
rect 28441 12202 28507 12205
rect 17493 12200 28507 12202
rect 17493 12144 17498 12200
rect 17554 12144 28446 12200
rect 28502 12144 28507 12200
rect 17493 12142 28507 12144
rect 17493 12139 17559 12142
rect 28441 12139 28507 12142
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 50290 11935 50606 11936
rect 14181 11930 14247 11933
rect 18229 11930 18295 11933
rect 14181 11928 18295 11930
rect 14181 11872 14186 11928
rect 14242 11872 18234 11928
rect 18290 11872 18295 11928
rect 14181 11870 18295 11872
rect 14181 11867 14247 11870
rect 18229 11867 18295 11870
rect 19701 11794 19767 11797
rect 20253 11794 20319 11797
rect 19701 11792 20319 11794
rect 19701 11736 19706 11792
rect 19762 11736 20258 11792
rect 20314 11736 20319 11792
rect 19701 11734 20319 11736
rect 19701 11731 19767 11734
rect 20253 11731 20319 11734
rect 12065 11658 12131 11661
rect 26969 11658 27035 11661
rect 12065 11656 27035 11658
rect 12065 11600 12070 11656
rect 12126 11600 26974 11656
rect 27030 11600 27035 11656
rect 12065 11598 27035 11600
rect 12065 11595 12131 11598
rect 26969 11595 27035 11598
rect 67633 11658 67699 11661
rect 69200 11658 70000 11688
rect 67633 11656 70000 11658
rect 67633 11600 67638 11656
rect 67694 11600 70000 11656
rect 67633 11598 70000 11600
rect 67633 11595 67699 11598
rect 69200 11568 70000 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 65650 11456 65966 11457
rect 65650 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65966 11456
rect 65650 11391 65966 11392
rect 19701 11386 19767 11389
rect 20069 11386 20135 11389
rect 19701 11384 20135 11386
rect 19701 11328 19706 11384
rect 19762 11328 20074 11384
rect 20130 11328 20135 11384
rect 19701 11326 20135 11328
rect 19701 11323 19767 11326
rect 20069 11323 20135 11326
rect 0 11160 800 11280
rect 19609 11250 19675 11253
rect 24945 11250 25011 11253
rect 19609 11248 25011 11250
rect 19609 11192 19614 11248
rect 19670 11192 24950 11248
rect 25006 11192 25011 11248
rect 19609 11190 25011 11192
rect 19609 11187 19675 11190
rect 24945 11187 25011 11190
rect 20110 11052 20116 11116
rect 20180 11114 20186 11116
rect 21357 11114 21423 11117
rect 20180 11112 21423 11114
rect 20180 11056 21362 11112
rect 21418 11056 21423 11112
rect 20180 11054 21423 11056
rect 20180 11052 20186 11054
rect 21357 11051 21423 11054
rect 17493 10980 17559 10981
rect 17493 10976 17540 10980
rect 17604 10978 17610 10980
rect 17493 10920 17498 10976
rect 17493 10916 17540 10920
rect 17604 10918 17650 10978
rect 17604 10916 17610 10918
rect 17493 10915 17559 10916
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 50290 10847 50606 10848
rect 24945 10842 25011 10845
rect 25405 10842 25471 10845
rect 24945 10840 25471 10842
rect 24945 10784 24950 10840
rect 25006 10784 25410 10840
rect 25466 10784 25471 10840
rect 24945 10782 25471 10784
rect 24945 10779 25011 10782
rect 25405 10779 25471 10782
rect 10041 10706 10107 10709
rect 28809 10706 28875 10709
rect 10041 10704 28875 10706
rect 10041 10648 10046 10704
rect 10102 10648 28814 10704
rect 28870 10648 28875 10704
rect 10041 10646 28875 10648
rect 10041 10643 10107 10646
rect 28809 10643 28875 10646
rect 10685 10570 10751 10573
rect 28993 10570 29059 10573
rect 10685 10568 29059 10570
rect 10685 10512 10690 10568
rect 10746 10512 28998 10568
rect 29054 10512 29059 10568
rect 10685 10510 29059 10512
rect 10685 10507 10751 10510
rect 28993 10507 29059 10510
rect 13905 10434 13971 10437
rect 24945 10434 25011 10437
rect 13905 10432 25011 10434
rect 13905 10376 13910 10432
rect 13966 10376 24950 10432
rect 25006 10376 25011 10432
rect 13905 10374 25011 10376
rect 13905 10371 13971 10374
rect 24945 10371 25011 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 65650 10368 65966 10369
rect 65650 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65966 10368
rect 65650 10303 65966 10304
rect 18321 10298 18387 10301
rect 22645 10298 22711 10301
rect 18321 10296 22711 10298
rect 18321 10240 18326 10296
rect 18382 10240 22650 10296
rect 22706 10240 22711 10296
rect 18321 10238 22711 10240
rect 18321 10235 18387 10238
rect 22645 10235 22711 10238
rect 67633 10298 67699 10301
rect 69200 10298 70000 10328
rect 67633 10296 70000 10298
rect 67633 10240 67638 10296
rect 67694 10240 70000 10296
rect 67633 10238 70000 10240
rect 67633 10235 67699 10238
rect 69200 10208 70000 10238
rect 19701 10162 19767 10165
rect 28533 10162 28599 10165
rect 19701 10160 28599 10162
rect 19701 10104 19706 10160
rect 19762 10104 28538 10160
rect 28594 10104 28599 10160
rect 19701 10102 28599 10104
rect 19701 10099 19767 10102
rect 28533 10099 28599 10102
rect 10961 10026 11027 10029
rect 28901 10026 28967 10029
rect 10961 10024 28967 10026
rect 10961 9968 10966 10024
rect 11022 9968 28906 10024
rect 28962 9968 28967 10024
rect 10961 9966 28967 9968
rect 10961 9963 11027 9966
rect 28901 9963 28967 9966
rect 20161 9890 20227 9893
rect 20294 9890 20300 9892
rect 20161 9888 20300 9890
rect 20161 9832 20166 9888
rect 20222 9832 20300 9888
rect 20161 9830 20300 9832
rect 20161 9827 20227 9830
rect 20294 9828 20300 9830
rect 20364 9828 20370 9892
rect 19570 9824 19886 9825
rect 0 9664 800 9784
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 50290 9759 50606 9760
rect 19977 9754 20043 9757
rect 20805 9754 20871 9757
rect 19977 9752 20871 9754
rect 19977 9696 19982 9752
rect 20038 9696 20810 9752
rect 20866 9696 20871 9752
rect 19977 9694 20871 9696
rect 19977 9691 20043 9694
rect 20805 9691 20871 9694
rect 8150 9556 8156 9620
rect 8220 9618 8226 9620
rect 11605 9618 11671 9621
rect 8220 9616 11671 9618
rect 8220 9560 11610 9616
rect 11666 9560 11671 9616
rect 8220 9558 11671 9560
rect 8220 9556 8226 9558
rect 11605 9555 11671 9558
rect 13118 9556 13124 9620
rect 13188 9618 13194 9620
rect 14365 9618 14431 9621
rect 17677 9620 17743 9621
rect 13188 9616 17602 9618
rect 13188 9560 14370 9616
rect 14426 9560 17602 9616
rect 13188 9558 17602 9560
rect 13188 9556 13194 9558
rect 14365 9555 14431 9558
rect 9765 9482 9831 9485
rect 16849 9482 16915 9485
rect 9765 9480 16915 9482
rect 9765 9424 9770 9480
rect 9826 9424 16854 9480
rect 16910 9424 16915 9480
rect 9765 9422 16915 9424
rect 17542 9482 17602 9558
rect 17677 9616 17724 9620
rect 17788 9618 17794 9620
rect 17953 9618 18019 9621
rect 28441 9618 28507 9621
rect 17677 9560 17682 9616
rect 17677 9556 17724 9560
rect 17788 9558 17834 9618
rect 17953 9616 28507 9618
rect 17953 9560 17958 9616
rect 18014 9560 28446 9616
rect 28502 9560 28507 9616
rect 17953 9558 28507 9560
rect 17788 9556 17794 9558
rect 17677 9555 17743 9556
rect 17953 9555 18019 9558
rect 28441 9555 28507 9558
rect 18413 9482 18479 9485
rect 17542 9480 18479 9482
rect 17542 9424 18418 9480
rect 18474 9424 18479 9480
rect 17542 9422 18479 9424
rect 9765 9419 9831 9422
rect 16849 9419 16915 9422
rect 18413 9419 18479 9422
rect 10501 9346 10567 9349
rect 27981 9346 28047 9349
rect 10501 9344 28047 9346
rect 10501 9288 10506 9344
rect 10562 9288 27986 9344
rect 28042 9288 28047 9344
rect 10501 9286 28047 9288
rect 10501 9283 10567 9286
rect 27981 9283 28047 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 65650 9280 65966 9281
rect 65650 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65966 9280
rect 65650 9215 65966 9216
rect 16982 9148 16988 9212
rect 17052 9210 17058 9212
rect 17125 9210 17191 9213
rect 17052 9208 17191 9210
rect 17052 9152 17130 9208
rect 17186 9152 17191 9208
rect 17052 9150 17191 9152
rect 17052 9148 17058 9150
rect 17125 9147 17191 9150
rect 24485 9210 24551 9213
rect 30833 9210 30899 9213
rect 24485 9208 30899 9210
rect 24485 9152 24490 9208
rect 24546 9152 30838 9208
rect 30894 9152 30899 9208
rect 24485 9150 30899 9152
rect 24485 9147 24551 9150
rect 30833 9147 30899 9150
rect 17769 9074 17835 9077
rect 29361 9074 29427 9077
rect 17769 9072 29427 9074
rect 17769 9016 17774 9072
rect 17830 9016 29366 9072
rect 29422 9016 29427 9072
rect 17769 9014 29427 9016
rect 17769 9011 17835 9014
rect 29361 9011 29427 9014
rect 19425 8938 19491 8941
rect 22461 8938 22527 8941
rect 19425 8936 22527 8938
rect 19425 8880 19430 8936
rect 19486 8880 22466 8936
rect 22522 8880 22527 8936
rect 19425 8878 22527 8880
rect 19425 8875 19491 8878
rect 22461 8875 22527 8878
rect 68093 8938 68159 8941
rect 69200 8938 70000 8968
rect 68093 8936 70000 8938
rect 68093 8880 68098 8936
rect 68154 8880 70000 8936
rect 68093 8878 70000 8880
rect 68093 8875 68159 8878
rect 69200 8848 70000 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 50290 8671 50606 8672
rect 19333 8530 19399 8533
rect 20253 8530 20319 8533
rect 19333 8528 20319 8530
rect 19333 8472 19338 8528
rect 19394 8472 20258 8528
rect 20314 8472 20319 8528
rect 19333 8470 20319 8472
rect 19333 8467 19399 8470
rect 20253 8467 20319 8470
rect 6862 8332 6868 8396
rect 6932 8394 6938 8396
rect 7833 8394 7899 8397
rect 6932 8392 7899 8394
rect 6932 8336 7838 8392
rect 7894 8336 7899 8392
rect 6932 8334 7899 8336
rect 6932 8332 6938 8334
rect 7833 8331 7899 8334
rect 13537 8394 13603 8397
rect 13670 8394 13676 8396
rect 13537 8392 13676 8394
rect 13537 8336 13542 8392
rect 13598 8336 13676 8392
rect 13537 8334 13676 8336
rect 13537 8331 13603 8334
rect 13670 8332 13676 8334
rect 13740 8332 13746 8396
rect 24209 8394 24275 8397
rect 33869 8394 33935 8397
rect 24209 8392 33935 8394
rect 24209 8336 24214 8392
rect 24270 8336 33874 8392
rect 33930 8336 33935 8392
rect 24209 8334 33935 8336
rect 24209 8331 24275 8334
rect 33869 8331 33935 8334
rect 0 8168 800 8288
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 65650 8192 65966 8193
rect 65650 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65966 8192
rect 65650 8127 65966 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 50290 7583 50606 7584
rect 68093 7578 68159 7581
rect 69200 7578 70000 7608
rect 68093 7576 70000 7578
rect 68093 7520 68098 7576
rect 68154 7520 70000 7576
rect 68093 7518 70000 7520
rect 68093 7515 68159 7518
rect 69200 7488 70000 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 65650 7104 65966 7105
rect 65650 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65966 7104
rect 65650 7039 65966 7040
rect 0 6672 800 6792
rect 9673 6626 9739 6629
rect 13537 6626 13603 6629
rect 9673 6624 13603 6626
rect 9673 6568 9678 6624
rect 9734 6568 13542 6624
rect 13598 6568 13603 6624
rect 9673 6566 13603 6568
rect 9673 6563 9739 6566
rect 13537 6563 13603 6566
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 50290 6495 50606 6496
rect 13629 6218 13695 6221
rect 19977 6218 20043 6221
rect 13629 6216 20043 6218
rect 13629 6160 13634 6216
rect 13690 6160 19982 6216
rect 20038 6160 20043 6216
rect 13629 6158 20043 6160
rect 13629 6155 13695 6158
rect 19977 6155 20043 6158
rect 67633 6218 67699 6221
rect 69200 6218 70000 6248
rect 67633 6216 70000 6218
rect 67633 6160 67638 6216
rect 67694 6160 70000 6216
rect 67633 6158 70000 6160
rect 67633 6155 67699 6158
rect 69200 6128 70000 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 65650 6016 65966 6017
rect 65650 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65966 6016
rect 65650 5951 65966 5952
rect 3233 5810 3299 5813
rect 6729 5810 6795 5813
rect 3233 5808 6795 5810
rect 3233 5752 3238 5808
rect 3294 5752 6734 5808
rect 6790 5752 6795 5808
rect 3233 5750 6795 5752
rect 3233 5747 3299 5750
rect 6729 5747 6795 5750
rect 13537 5674 13603 5677
rect 14917 5674 14983 5677
rect 13537 5672 14983 5674
rect 13537 5616 13542 5672
rect 13598 5616 14922 5672
rect 14978 5616 14983 5672
rect 13537 5614 14983 5616
rect 13537 5611 13603 5614
rect 14917 5611 14983 5614
rect 16430 5612 16436 5676
rect 16500 5674 16506 5676
rect 17902 5674 17908 5676
rect 16500 5614 17908 5674
rect 16500 5612 16506 5614
rect 17902 5612 17908 5614
rect 17972 5674 17978 5676
rect 19609 5674 19675 5677
rect 17972 5672 19675 5674
rect 17972 5616 19614 5672
rect 19670 5616 19675 5672
rect 17972 5614 19675 5616
rect 17972 5612 17978 5614
rect 19609 5611 19675 5614
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 50290 5407 50606 5408
rect 0 5176 800 5296
rect 13721 4994 13787 4997
rect 17217 4994 17283 4997
rect 13721 4992 17283 4994
rect 13721 4936 13726 4992
rect 13782 4936 17222 4992
rect 17278 4936 17283 4992
rect 13721 4934 17283 4936
rect 13721 4931 13787 4934
rect 17217 4931 17283 4934
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 65650 4928 65966 4929
rect 65650 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65966 4928
rect 65650 4863 65966 4864
rect 13353 4858 13419 4861
rect 17677 4858 17743 4861
rect 13353 4856 17743 4858
rect 13353 4800 13358 4856
rect 13414 4800 17682 4856
rect 17738 4800 17743 4856
rect 13353 4798 17743 4800
rect 13353 4795 13419 4798
rect 17677 4795 17743 4798
rect 67633 4858 67699 4861
rect 69200 4858 70000 4888
rect 67633 4856 70000 4858
rect 67633 4800 67638 4856
rect 67694 4800 70000 4856
rect 67633 4798 70000 4800
rect 67633 4795 67699 4798
rect 69200 4768 70000 4798
rect 7465 4722 7531 4725
rect 16021 4722 16087 4725
rect 7465 4720 16087 4722
rect 7465 4664 7470 4720
rect 7526 4664 16026 4720
rect 16082 4664 16087 4720
rect 7465 4662 16087 4664
rect 7465 4659 7531 4662
rect 16021 4659 16087 4662
rect 8385 4450 8451 4453
rect 11605 4450 11671 4453
rect 8385 4448 11671 4450
rect 8385 4392 8390 4448
rect 8446 4392 11610 4448
rect 11666 4392 11671 4448
rect 8385 4390 11671 4392
rect 8385 4387 8451 4390
rect 11605 4387 11671 4390
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 50290 4319 50606 4320
rect 9765 4178 9831 4181
rect 13353 4178 13419 4181
rect 9765 4176 13419 4178
rect 9765 4120 9770 4176
rect 9826 4120 13358 4176
rect 13414 4120 13419 4176
rect 9765 4118 13419 4120
rect 9765 4115 9831 4118
rect 13353 4115 13419 4118
rect 4245 4042 4311 4045
rect 6862 4042 6868 4044
rect 4245 4040 6868 4042
rect 4245 3984 4250 4040
rect 4306 3984 6868 4040
rect 4245 3982 6868 3984
rect 4245 3979 4311 3982
rect 6862 3980 6868 3982
rect 6932 3980 6938 4044
rect 12893 4042 12959 4045
rect 13721 4044 13787 4045
rect 13118 4042 13124 4044
rect 12893 4040 13124 4042
rect 12893 3984 12898 4040
rect 12954 3984 13124 4040
rect 12893 3982 13124 3984
rect 12893 3979 12959 3982
rect 13118 3980 13124 3982
rect 13188 3980 13194 4044
rect 13670 3980 13676 4044
rect 13740 4042 13787 4044
rect 13740 4040 13832 4042
rect 13782 3984 13832 4040
rect 13740 3982 13832 3984
rect 13740 3980 13787 3982
rect 13721 3979 13787 3980
rect 6729 3906 6795 3909
rect 7189 3906 7255 3909
rect 7925 3906 7991 3909
rect 15101 3906 15167 3909
rect 6729 3904 15167 3906
rect 6729 3848 6734 3904
rect 6790 3848 7194 3904
rect 7250 3848 7930 3904
rect 7986 3848 15106 3904
rect 15162 3848 15167 3904
rect 6729 3846 15167 3848
rect 6729 3843 6795 3846
rect 7189 3843 7255 3846
rect 7925 3843 7991 3846
rect 15101 3843 15167 3846
rect 4210 3840 4526 3841
rect 0 3680 800 3800
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 65650 3840 65966 3841
rect 65650 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65966 3840
rect 65650 3775 65966 3776
rect 5073 3770 5139 3773
rect 10961 3770 11027 3773
rect 5073 3768 11027 3770
rect 5073 3712 5078 3768
rect 5134 3712 10966 3768
rect 11022 3712 11027 3768
rect 5073 3710 11027 3712
rect 5073 3707 5139 3710
rect 10961 3707 11027 3710
rect 7925 3634 7991 3637
rect 8385 3634 8451 3637
rect 7925 3632 8451 3634
rect 7925 3576 7930 3632
rect 7986 3576 8390 3632
rect 8446 3576 8451 3632
rect 7925 3574 8451 3576
rect 7925 3571 7991 3574
rect 8385 3571 8451 3574
rect 9673 3634 9739 3637
rect 14365 3634 14431 3637
rect 19241 3634 19307 3637
rect 9673 3632 19307 3634
rect 9673 3576 9678 3632
rect 9734 3576 14370 3632
rect 14426 3576 19246 3632
rect 19302 3576 19307 3632
rect 9673 3574 19307 3576
rect 9673 3571 9739 3574
rect 14365 3571 14431 3574
rect 19241 3571 19307 3574
rect 10409 3498 10475 3501
rect 20069 3498 20135 3501
rect 10409 3496 20135 3498
rect 10409 3440 10414 3496
rect 10470 3440 20074 3496
rect 20130 3440 20135 3496
rect 10409 3438 20135 3440
rect 10409 3435 10475 3438
rect 20069 3435 20135 3438
rect 68093 3498 68159 3501
rect 69200 3498 70000 3528
rect 68093 3496 70000 3498
rect 68093 3440 68098 3496
rect 68154 3440 70000 3496
rect 68093 3438 70000 3440
rect 68093 3435 68159 3438
rect 69200 3408 70000 3438
rect 2221 3362 2287 3365
rect 10041 3362 10107 3365
rect 2221 3360 10107 3362
rect 2221 3304 2226 3360
rect 2282 3304 10046 3360
rect 10102 3304 10107 3360
rect 2221 3302 10107 3304
rect 2221 3299 2287 3302
rect 10041 3299 10107 3302
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 50290 3231 50606 3232
rect 7281 3226 7347 3229
rect 13445 3226 13511 3229
rect 7281 3224 13511 3226
rect 7281 3168 7286 3224
rect 7342 3168 13450 3224
rect 13506 3168 13511 3224
rect 7281 3166 13511 3168
rect 7281 3163 7347 3166
rect 13445 3163 13511 3166
rect 57881 3226 57947 3229
rect 60457 3226 60523 3229
rect 57881 3224 60523 3226
rect 57881 3168 57886 3224
rect 57942 3168 60462 3224
rect 60518 3168 60523 3224
rect 57881 3166 60523 3168
rect 57881 3163 57947 3166
rect 60457 3163 60523 3166
rect 5257 3090 5323 3093
rect 13261 3090 13327 3093
rect 5257 3088 13327 3090
rect 5257 3032 5262 3088
rect 5318 3032 13266 3088
rect 13322 3032 13327 3088
rect 5257 3030 13327 3032
rect 5257 3027 5323 3030
rect 13261 3027 13327 3030
rect 6545 2954 6611 2957
rect 12249 2954 12315 2957
rect 6545 2952 12315 2954
rect 6545 2896 6550 2952
rect 6606 2896 12254 2952
rect 12310 2896 12315 2952
rect 6545 2894 12315 2896
rect 6545 2891 6611 2894
rect 12249 2891 12315 2894
rect 13261 2954 13327 2957
rect 17125 2954 17191 2957
rect 13261 2952 17191 2954
rect 13261 2896 13266 2952
rect 13322 2896 17130 2952
rect 17186 2896 17191 2952
rect 13261 2894 17191 2896
rect 13261 2891 13327 2894
rect 17125 2891 17191 2894
rect 17769 2954 17835 2957
rect 17902 2954 17908 2956
rect 17769 2952 17908 2954
rect 17769 2896 17774 2952
rect 17830 2896 17908 2952
rect 17769 2894 17908 2896
rect 17769 2891 17835 2894
rect 17902 2892 17908 2894
rect 17972 2954 17978 2956
rect 26325 2954 26391 2957
rect 17972 2952 26391 2954
rect 17972 2896 26330 2952
rect 26386 2896 26391 2952
rect 17972 2894 26391 2896
rect 17972 2892 17978 2894
rect 26325 2891 26391 2894
rect 5625 2818 5691 2821
rect 11513 2818 11579 2821
rect 5625 2816 11579 2818
rect 5625 2760 5630 2816
rect 5686 2760 11518 2816
rect 11574 2760 11579 2816
rect 5625 2758 11579 2760
rect 5625 2755 5691 2758
rect 11513 2755 11579 2758
rect 13261 2818 13327 2821
rect 17585 2818 17651 2821
rect 13261 2816 17651 2818
rect 13261 2760 13266 2816
rect 13322 2760 17590 2816
rect 17646 2760 17651 2816
rect 13261 2758 17651 2760
rect 13261 2755 13327 2758
rect 17585 2755 17651 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 65650 2752 65966 2753
rect 65650 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65966 2752
rect 65650 2687 65966 2688
rect 7649 2682 7715 2685
rect 8150 2682 8156 2684
rect 7649 2680 8156 2682
rect 7649 2624 7654 2680
rect 7710 2624 8156 2680
rect 7649 2622 8156 2624
rect 7649 2619 7715 2622
rect 8150 2620 8156 2622
rect 8220 2620 8226 2684
rect 5441 2546 5507 2549
rect 14825 2546 14891 2549
rect 20110 2546 20116 2548
rect 5441 2544 20116 2546
rect 5441 2488 5446 2544
rect 5502 2488 14830 2544
rect 14886 2488 20116 2544
rect 5441 2486 20116 2488
rect 5441 2483 5507 2486
rect 14825 2483 14891 2486
rect 20110 2484 20116 2486
rect 20180 2484 20186 2548
rect 2405 2410 2471 2413
rect 12985 2410 13051 2413
rect 20294 2410 20300 2412
rect 2405 2408 20300 2410
rect 2405 2352 2410 2408
rect 2466 2352 12990 2408
rect 13046 2352 20300 2408
rect 2405 2350 20300 2352
rect 2405 2347 2471 2350
rect 12985 2347 13051 2350
rect 20294 2348 20300 2350
rect 20364 2348 20370 2412
rect 0 2184 800 2304
rect 3325 2274 3391 2277
rect 10041 2274 10107 2277
rect 3325 2272 10107 2274
rect 3325 2216 3330 2272
rect 3386 2216 10046 2272
rect 10102 2216 10107 2272
rect 3325 2214 10107 2216
rect 3325 2211 3391 2214
rect 10041 2211 10107 2214
rect 10409 2274 10475 2277
rect 16982 2274 16988 2276
rect 10409 2272 16988 2274
rect 10409 2216 10414 2272
rect 10470 2216 16988 2272
rect 10409 2214 16988 2216
rect 10409 2211 10475 2214
rect 16982 2212 16988 2214
rect 17052 2212 17058 2276
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 50290 2143 50606 2144
rect 6821 2138 6887 2141
rect 14222 2138 14228 2140
rect 6821 2136 14228 2138
rect 6821 2080 6826 2136
rect 6882 2080 14228 2136
rect 6821 2078 14228 2080
rect 6821 2075 6887 2078
rect 14222 2076 14228 2078
rect 14292 2138 14298 2140
rect 16757 2138 16823 2141
rect 14292 2136 16823 2138
rect 14292 2080 16762 2136
rect 16818 2080 16823 2136
rect 14292 2078 16823 2080
rect 14292 2076 14298 2078
rect 16757 2075 16823 2078
rect 66989 2138 67055 2141
rect 69200 2138 70000 2168
rect 66989 2136 70000 2138
rect 66989 2080 66994 2136
rect 67050 2080 70000 2136
rect 66989 2078 70000 2080
rect 66989 2075 67055 2078
rect 69200 2048 70000 2078
rect 67541 778 67607 781
rect 69200 778 70000 808
rect 67541 776 70000 778
rect 67541 720 67546 776
rect 67602 720 70000 776
rect 67541 718 70000 720
rect 67541 715 67607 718
rect 69200 688 70000 718
<< via3 >>
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 65656 57148 65720 57152
rect 65656 57092 65660 57148
rect 65660 57092 65716 57148
rect 65716 57092 65720 57148
rect 65656 57088 65720 57092
rect 65736 57148 65800 57152
rect 65736 57092 65740 57148
rect 65740 57092 65796 57148
rect 65796 57092 65800 57148
rect 65736 57088 65800 57092
rect 65816 57148 65880 57152
rect 65816 57092 65820 57148
rect 65820 57092 65876 57148
rect 65876 57092 65880 57148
rect 65816 57088 65880 57092
rect 65896 57148 65960 57152
rect 65896 57092 65900 57148
rect 65900 57092 65956 57148
rect 65956 57092 65960 57148
rect 65896 57088 65960 57092
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 65656 56060 65720 56064
rect 65656 56004 65660 56060
rect 65660 56004 65716 56060
rect 65716 56004 65720 56060
rect 65656 56000 65720 56004
rect 65736 56060 65800 56064
rect 65736 56004 65740 56060
rect 65740 56004 65796 56060
rect 65796 56004 65800 56060
rect 65736 56000 65800 56004
rect 65816 56060 65880 56064
rect 65816 56004 65820 56060
rect 65820 56004 65876 56060
rect 65876 56004 65880 56060
rect 65816 56000 65880 56004
rect 65896 56060 65960 56064
rect 65896 56004 65900 56060
rect 65900 56004 65956 56060
rect 65956 56004 65960 56060
rect 65896 56000 65960 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 65656 54972 65720 54976
rect 65656 54916 65660 54972
rect 65660 54916 65716 54972
rect 65716 54916 65720 54972
rect 65656 54912 65720 54916
rect 65736 54972 65800 54976
rect 65736 54916 65740 54972
rect 65740 54916 65796 54972
rect 65796 54916 65800 54972
rect 65736 54912 65800 54916
rect 65816 54972 65880 54976
rect 65816 54916 65820 54972
rect 65820 54916 65876 54972
rect 65876 54916 65880 54972
rect 65816 54912 65880 54916
rect 65896 54972 65960 54976
rect 65896 54916 65900 54972
rect 65900 54916 65956 54972
rect 65956 54916 65960 54972
rect 65896 54912 65960 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 65656 53884 65720 53888
rect 65656 53828 65660 53884
rect 65660 53828 65716 53884
rect 65716 53828 65720 53884
rect 65656 53824 65720 53828
rect 65736 53884 65800 53888
rect 65736 53828 65740 53884
rect 65740 53828 65796 53884
rect 65796 53828 65800 53884
rect 65736 53824 65800 53828
rect 65816 53884 65880 53888
rect 65816 53828 65820 53884
rect 65820 53828 65876 53884
rect 65876 53828 65880 53884
rect 65816 53824 65880 53828
rect 65896 53884 65960 53888
rect 65896 53828 65900 53884
rect 65900 53828 65956 53884
rect 65956 53828 65960 53884
rect 65896 53824 65960 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 65656 52796 65720 52800
rect 65656 52740 65660 52796
rect 65660 52740 65716 52796
rect 65716 52740 65720 52796
rect 65656 52736 65720 52740
rect 65736 52796 65800 52800
rect 65736 52740 65740 52796
rect 65740 52740 65796 52796
rect 65796 52740 65800 52796
rect 65736 52736 65800 52740
rect 65816 52796 65880 52800
rect 65816 52740 65820 52796
rect 65820 52740 65876 52796
rect 65876 52740 65880 52796
rect 65816 52736 65880 52740
rect 65896 52796 65960 52800
rect 65896 52740 65900 52796
rect 65900 52740 65956 52796
rect 65956 52740 65960 52796
rect 65896 52736 65960 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 65656 51708 65720 51712
rect 65656 51652 65660 51708
rect 65660 51652 65716 51708
rect 65716 51652 65720 51708
rect 65656 51648 65720 51652
rect 65736 51708 65800 51712
rect 65736 51652 65740 51708
rect 65740 51652 65796 51708
rect 65796 51652 65800 51708
rect 65736 51648 65800 51652
rect 65816 51708 65880 51712
rect 65816 51652 65820 51708
rect 65820 51652 65876 51708
rect 65876 51652 65880 51708
rect 65816 51648 65880 51652
rect 65896 51708 65960 51712
rect 65896 51652 65900 51708
rect 65900 51652 65956 51708
rect 65956 51652 65960 51708
rect 65896 51648 65960 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 65656 50620 65720 50624
rect 65656 50564 65660 50620
rect 65660 50564 65716 50620
rect 65716 50564 65720 50620
rect 65656 50560 65720 50564
rect 65736 50620 65800 50624
rect 65736 50564 65740 50620
rect 65740 50564 65796 50620
rect 65796 50564 65800 50620
rect 65736 50560 65800 50564
rect 65816 50620 65880 50624
rect 65816 50564 65820 50620
rect 65820 50564 65876 50620
rect 65876 50564 65880 50620
rect 65816 50560 65880 50564
rect 65896 50620 65960 50624
rect 65896 50564 65900 50620
rect 65900 50564 65956 50620
rect 65956 50564 65960 50620
rect 65896 50560 65960 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 65656 49532 65720 49536
rect 65656 49476 65660 49532
rect 65660 49476 65716 49532
rect 65716 49476 65720 49532
rect 65656 49472 65720 49476
rect 65736 49532 65800 49536
rect 65736 49476 65740 49532
rect 65740 49476 65796 49532
rect 65796 49476 65800 49532
rect 65736 49472 65800 49476
rect 65816 49532 65880 49536
rect 65816 49476 65820 49532
rect 65820 49476 65876 49532
rect 65876 49476 65880 49532
rect 65816 49472 65880 49476
rect 65896 49532 65960 49536
rect 65896 49476 65900 49532
rect 65900 49476 65956 49532
rect 65956 49476 65960 49532
rect 65896 49472 65960 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 65656 48444 65720 48448
rect 65656 48388 65660 48444
rect 65660 48388 65716 48444
rect 65716 48388 65720 48444
rect 65656 48384 65720 48388
rect 65736 48444 65800 48448
rect 65736 48388 65740 48444
rect 65740 48388 65796 48444
rect 65796 48388 65800 48444
rect 65736 48384 65800 48388
rect 65816 48444 65880 48448
rect 65816 48388 65820 48444
rect 65820 48388 65876 48444
rect 65876 48388 65880 48444
rect 65816 48384 65880 48388
rect 65896 48444 65960 48448
rect 65896 48388 65900 48444
rect 65900 48388 65956 48444
rect 65956 48388 65960 48444
rect 65896 48384 65960 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 65656 47356 65720 47360
rect 65656 47300 65660 47356
rect 65660 47300 65716 47356
rect 65716 47300 65720 47356
rect 65656 47296 65720 47300
rect 65736 47356 65800 47360
rect 65736 47300 65740 47356
rect 65740 47300 65796 47356
rect 65796 47300 65800 47356
rect 65736 47296 65800 47300
rect 65816 47356 65880 47360
rect 65816 47300 65820 47356
rect 65820 47300 65876 47356
rect 65876 47300 65880 47356
rect 65816 47296 65880 47300
rect 65896 47356 65960 47360
rect 65896 47300 65900 47356
rect 65900 47300 65956 47356
rect 65956 47300 65960 47356
rect 65896 47296 65960 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 65656 46268 65720 46272
rect 65656 46212 65660 46268
rect 65660 46212 65716 46268
rect 65716 46212 65720 46268
rect 65656 46208 65720 46212
rect 65736 46268 65800 46272
rect 65736 46212 65740 46268
rect 65740 46212 65796 46268
rect 65796 46212 65800 46268
rect 65736 46208 65800 46212
rect 65816 46268 65880 46272
rect 65816 46212 65820 46268
rect 65820 46212 65876 46268
rect 65876 46212 65880 46268
rect 65816 46208 65880 46212
rect 65896 46268 65960 46272
rect 65896 46212 65900 46268
rect 65900 46212 65956 46268
rect 65956 46212 65960 46268
rect 65896 46208 65960 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 65656 45180 65720 45184
rect 65656 45124 65660 45180
rect 65660 45124 65716 45180
rect 65716 45124 65720 45180
rect 65656 45120 65720 45124
rect 65736 45180 65800 45184
rect 65736 45124 65740 45180
rect 65740 45124 65796 45180
rect 65796 45124 65800 45180
rect 65736 45120 65800 45124
rect 65816 45180 65880 45184
rect 65816 45124 65820 45180
rect 65820 45124 65876 45180
rect 65876 45124 65880 45180
rect 65816 45120 65880 45124
rect 65896 45180 65960 45184
rect 65896 45124 65900 45180
rect 65900 45124 65956 45180
rect 65956 45124 65960 45180
rect 65896 45120 65960 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 65656 44092 65720 44096
rect 65656 44036 65660 44092
rect 65660 44036 65716 44092
rect 65716 44036 65720 44092
rect 65656 44032 65720 44036
rect 65736 44092 65800 44096
rect 65736 44036 65740 44092
rect 65740 44036 65796 44092
rect 65796 44036 65800 44092
rect 65736 44032 65800 44036
rect 65816 44092 65880 44096
rect 65816 44036 65820 44092
rect 65820 44036 65876 44092
rect 65876 44036 65880 44092
rect 65816 44032 65880 44036
rect 65896 44092 65960 44096
rect 65896 44036 65900 44092
rect 65900 44036 65956 44092
rect 65956 44036 65960 44092
rect 65896 44032 65960 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 65656 43004 65720 43008
rect 65656 42948 65660 43004
rect 65660 42948 65716 43004
rect 65716 42948 65720 43004
rect 65656 42944 65720 42948
rect 65736 43004 65800 43008
rect 65736 42948 65740 43004
rect 65740 42948 65796 43004
rect 65796 42948 65800 43004
rect 65736 42944 65800 42948
rect 65816 43004 65880 43008
rect 65816 42948 65820 43004
rect 65820 42948 65876 43004
rect 65876 42948 65880 43004
rect 65816 42944 65880 42948
rect 65896 43004 65960 43008
rect 65896 42948 65900 43004
rect 65900 42948 65956 43004
rect 65956 42948 65960 43004
rect 65896 42944 65960 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 65656 41916 65720 41920
rect 65656 41860 65660 41916
rect 65660 41860 65716 41916
rect 65716 41860 65720 41916
rect 65656 41856 65720 41860
rect 65736 41916 65800 41920
rect 65736 41860 65740 41916
rect 65740 41860 65796 41916
rect 65796 41860 65800 41916
rect 65736 41856 65800 41860
rect 65816 41916 65880 41920
rect 65816 41860 65820 41916
rect 65820 41860 65876 41916
rect 65876 41860 65880 41916
rect 65816 41856 65880 41860
rect 65896 41916 65960 41920
rect 65896 41860 65900 41916
rect 65900 41860 65956 41916
rect 65956 41860 65960 41916
rect 65896 41856 65960 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 65656 40828 65720 40832
rect 65656 40772 65660 40828
rect 65660 40772 65716 40828
rect 65716 40772 65720 40828
rect 65656 40768 65720 40772
rect 65736 40828 65800 40832
rect 65736 40772 65740 40828
rect 65740 40772 65796 40828
rect 65796 40772 65800 40828
rect 65736 40768 65800 40772
rect 65816 40828 65880 40832
rect 65816 40772 65820 40828
rect 65820 40772 65876 40828
rect 65876 40772 65880 40828
rect 65816 40768 65880 40772
rect 65896 40828 65960 40832
rect 65896 40772 65900 40828
rect 65900 40772 65956 40828
rect 65956 40772 65960 40828
rect 65896 40768 65960 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 65656 39740 65720 39744
rect 65656 39684 65660 39740
rect 65660 39684 65716 39740
rect 65716 39684 65720 39740
rect 65656 39680 65720 39684
rect 65736 39740 65800 39744
rect 65736 39684 65740 39740
rect 65740 39684 65796 39740
rect 65796 39684 65800 39740
rect 65736 39680 65800 39684
rect 65816 39740 65880 39744
rect 65816 39684 65820 39740
rect 65820 39684 65876 39740
rect 65876 39684 65880 39740
rect 65816 39680 65880 39684
rect 65896 39740 65960 39744
rect 65896 39684 65900 39740
rect 65900 39684 65956 39740
rect 65956 39684 65960 39740
rect 65896 39680 65960 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 65656 38652 65720 38656
rect 65656 38596 65660 38652
rect 65660 38596 65716 38652
rect 65716 38596 65720 38652
rect 65656 38592 65720 38596
rect 65736 38652 65800 38656
rect 65736 38596 65740 38652
rect 65740 38596 65796 38652
rect 65796 38596 65800 38652
rect 65736 38592 65800 38596
rect 65816 38652 65880 38656
rect 65816 38596 65820 38652
rect 65820 38596 65876 38652
rect 65876 38596 65880 38652
rect 65816 38592 65880 38596
rect 65896 38652 65960 38656
rect 65896 38596 65900 38652
rect 65900 38596 65956 38652
rect 65956 38596 65960 38652
rect 65896 38592 65960 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 65656 37564 65720 37568
rect 65656 37508 65660 37564
rect 65660 37508 65716 37564
rect 65716 37508 65720 37564
rect 65656 37504 65720 37508
rect 65736 37564 65800 37568
rect 65736 37508 65740 37564
rect 65740 37508 65796 37564
rect 65796 37508 65800 37564
rect 65736 37504 65800 37508
rect 65816 37564 65880 37568
rect 65816 37508 65820 37564
rect 65820 37508 65876 37564
rect 65876 37508 65880 37564
rect 65816 37504 65880 37508
rect 65896 37564 65960 37568
rect 65896 37508 65900 37564
rect 65900 37508 65956 37564
rect 65956 37508 65960 37564
rect 65896 37504 65960 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 65656 36476 65720 36480
rect 65656 36420 65660 36476
rect 65660 36420 65716 36476
rect 65716 36420 65720 36476
rect 65656 36416 65720 36420
rect 65736 36476 65800 36480
rect 65736 36420 65740 36476
rect 65740 36420 65796 36476
rect 65796 36420 65800 36476
rect 65736 36416 65800 36420
rect 65816 36476 65880 36480
rect 65816 36420 65820 36476
rect 65820 36420 65876 36476
rect 65876 36420 65880 36476
rect 65816 36416 65880 36420
rect 65896 36476 65960 36480
rect 65896 36420 65900 36476
rect 65900 36420 65956 36476
rect 65956 36420 65960 36476
rect 65896 36416 65960 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 65656 35388 65720 35392
rect 65656 35332 65660 35388
rect 65660 35332 65716 35388
rect 65716 35332 65720 35388
rect 65656 35328 65720 35332
rect 65736 35388 65800 35392
rect 65736 35332 65740 35388
rect 65740 35332 65796 35388
rect 65796 35332 65800 35388
rect 65736 35328 65800 35332
rect 65816 35388 65880 35392
rect 65816 35332 65820 35388
rect 65820 35332 65876 35388
rect 65876 35332 65880 35388
rect 65816 35328 65880 35332
rect 65896 35388 65960 35392
rect 65896 35332 65900 35388
rect 65900 35332 65956 35388
rect 65956 35332 65960 35388
rect 65896 35328 65960 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 65656 34300 65720 34304
rect 65656 34244 65660 34300
rect 65660 34244 65716 34300
rect 65716 34244 65720 34300
rect 65656 34240 65720 34244
rect 65736 34300 65800 34304
rect 65736 34244 65740 34300
rect 65740 34244 65796 34300
rect 65796 34244 65800 34300
rect 65736 34240 65800 34244
rect 65816 34300 65880 34304
rect 65816 34244 65820 34300
rect 65820 34244 65876 34300
rect 65876 34244 65880 34300
rect 65816 34240 65880 34244
rect 65896 34300 65960 34304
rect 65896 34244 65900 34300
rect 65900 34244 65956 34300
rect 65956 34244 65960 34300
rect 65896 34240 65960 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 65656 33212 65720 33216
rect 65656 33156 65660 33212
rect 65660 33156 65716 33212
rect 65716 33156 65720 33212
rect 65656 33152 65720 33156
rect 65736 33212 65800 33216
rect 65736 33156 65740 33212
rect 65740 33156 65796 33212
rect 65796 33156 65800 33212
rect 65736 33152 65800 33156
rect 65816 33212 65880 33216
rect 65816 33156 65820 33212
rect 65820 33156 65876 33212
rect 65876 33156 65880 33212
rect 65816 33152 65880 33156
rect 65896 33212 65960 33216
rect 65896 33156 65900 33212
rect 65900 33156 65956 33212
rect 65956 33156 65960 33212
rect 65896 33152 65960 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 65656 32124 65720 32128
rect 65656 32068 65660 32124
rect 65660 32068 65716 32124
rect 65716 32068 65720 32124
rect 65656 32064 65720 32068
rect 65736 32124 65800 32128
rect 65736 32068 65740 32124
rect 65740 32068 65796 32124
rect 65796 32068 65800 32124
rect 65736 32064 65800 32068
rect 65816 32124 65880 32128
rect 65816 32068 65820 32124
rect 65820 32068 65876 32124
rect 65876 32068 65880 32124
rect 65816 32064 65880 32068
rect 65896 32124 65960 32128
rect 65896 32068 65900 32124
rect 65900 32068 65956 32124
rect 65956 32068 65960 32124
rect 65896 32064 65960 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 65656 31036 65720 31040
rect 65656 30980 65660 31036
rect 65660 30980 65716 31036
rect 65716 30980 65720 31036
rect 65656 30976 65720 30980
rect 65736 31036 65800 31040
rect 65736 30980 65740 31036
rect 65740 30980 65796 31036
rect 65796 30980 65800 31036
rect 65736 30976 65800 30980
rect 65816 31036 65880 31040
rect 65816 30980 65820 31036
rect 65820 30980 65876 31036
rect 65876 30980 65880 31036
rect 65816 30976 65880 30980
rect 65896 31036 65960 31040
rect 65896 30980 65900 31036
rect 65900 30980 65956 31036
rect 65956 30980 65960 31036
rect 65896 30976 65960 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 65656 29948 65720 29952
rect 65656 29892 65660 29948
rect 65660 29892 65716 29948
rect 65716 29892 65720 29948
rect 65656 29888 65720 29892
rect 65736 29948 65800 29952
rect 65736 29892 65740 29948
rect 65740 29892 65796 29948
rect 65796 29892 65800 29948
rect 65736 29888 65800 29892
rect 65816 29948 65880 29952
rect 65816 29892 65820 29948
rect 65820 29892 65876 29948
rect 65876 29892 65880 29948
rect 65816 29888 65880 29892
rect 65896 29948 65960 29952
rect 65896 29892 65900 29948
rect 65900 29892 65956 29948
rect 65956 29892 65960 29948
rect 65896 29888 65960 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 65656 28860 65720 28864
rect 65656 28804 65660 28860
rect 65660 28804 65716 28860
rect 65716 28804 65720 28860
rect 65656 28800 65720 28804
rect 65736 28860 65800 28864
rect 65736 28804 65740 28860
rect 65740 28804 65796 28860
rect 65796 28804 65800 28860
rect 65736 28800 65800 28804
rect 65816 28860 65880 28864
rect 65816 28804 65820 28860
rect 65820 28804 65876 28860
rect 65876 28804 65880 28860
rect 65816 28800 65880 28804
rect 65896 28860 65960 28864
rect 65896 28804 65900 28860
rect 65900 28804 65956 28860
rect 65956 28804 65960 28860
rect 65896 28800 65960 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 65656 27772 65720 27776
rect 65656 27716 65660 27772
rect 65660 27716 65716 27772
rect 65716 27716 65720 27772
rect 65656 27712 65720 27716
rect 65736 27772 65800 27776
rect 65736 27716 65740 27772
rect 65740 27716 65796 27772
rect 65796 27716 65800 27772
rect 65736 27712 65800 27716
rect 65816 27772 65880 27776
rect 65816 27716 65820 27772
rect 65820 27716 65876 27772
rect 65876 27716 65880 27772
rect 65816 27712 65880 27716
rect 65896 27772 65960 27776
rect 65896 27716 65900 27772
rect 65900 27716 65956 27772
rect 65956 27716 65960 27772
rect 65896 27712 65960 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 65656 26684 65720 26688
rect 65656 26628 65660 26684
rect 65660 26628 65716 26684
rect 65716 26628 65720 26684
rect 65656 26624 65720 26628
rect 65736 26684 65800 26688
rect 65736 26628 65740 26684
rect 65740 26628 65796 26684
rect 65796 26628 65800 26684
rect 65736 26624 65800 26628
rect 65816 26684 65880 26688
rect 65816 26628 65820 26684
rect 65820 26628 65876 26684
rect 65876 26628 65880 26684
rect 65816 26624 65880 26628
rect 65896 26684 65960 26688
rect 65896 26628 65900 26684
rect 65900 26628 65956 26684
rect 65956 26628 65960 26684
rect 65896 26624 65960 26628
rect 17540 26284 17604 26348
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 65656 25596 65720 25600
rect 65656 25540 65660 25596
rect 65660 25540 65716 25596
rect 65716 25540 65720 25596
rect 65656 25536 65720 25540
rect 65736 25596 65800 25600
rect 65736 25540 65740 25596
rect 65740 25540 65796 25596
rect 65796 25540 65800 25596
rect 65736 25536 65800 25540
rect 65816 25596 65880 25600
rect 65816 25540 65820 25596
rect 65820 25540 65876 25596
rect 65876 25540 65880 25596
rect 65816 25536 65880 25540
rect 65896 25596 65960 25600
rect 65896 25540 65900 25596
rect 65900 25540 65956 25596
rect 65956 25540 65960 25596
rect 65896 25536 65960 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 17724 24984 17788 24988
rect 17724 24928 17738 24984
rect 17738 24928 17788 24984
rect 17724 24924 17788 24928
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 65656 24508 65720 24512
rect 65656 24452 65660 24508
rect 65660 24452 65716 24508
rect 65716 24452 65720 24508
rect 65656 24448 65720 24452
rect 65736 24508 65800 24512
rect 65736 24452 65740 24508
rect 65740 24452 65796 24508
rect 65796 24452 65800 24508
rect 65736 24448 65800 24452
rect 65816 24508 65880 24512
rect 65816 24452 65820 24508
rect 65820 24452 65876 24508
rect 65876 24452 65880 24508
rect 65816 24448 65880 24452
rect 65896 24508 65960 24512
rect 65896 24452 65900 24508
rect 65900 24452 65956 24508
rect 65956 24452 65960 24508
rect 65896 24448 65960 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 65656 23420 65720 23424
rect 65656 23364 65660 23420
rect 65660 23364 65716 23420
rect 65716 23364 65720 23420
rect 65656 23360 65720 23364
rect 65736 23420 65800 23424
rect 65736 23364 65740 23420
rect 65740 23364 65796 23420
rect 65796 23364 65800 23420
rect 65736 23360 65800 23364
rect 65816 23420 65880 23424
rect 65816 23364 65820 23420
rect 65820 23364 65876 23420
rect 65876 23364 65880 23420
rect 65816 23360 65880 23364
rect 65896 23420 65960 23424
rect 65896 23364 65900 23420
rect 65900 23364 65956 23420
rect 65956 23364 65960 23420
rect 65896 23360 65960 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 65656 22332 65720 22336
rect 65656 22276 65660 22332
rect 65660 22276 65716 22332
rect 65716 22276 65720 22332
rect 65656 22272 65720 22276
rect 65736 22332 65800 22336
rect 65736 22276 65740 22332
rect 65740 22276 65796 22332
rect 65796 22276 65800 22332
rect 65736 22272 65800 22276
rect 65816 22332 65880 22336
rect 65816 22276 65820 22332
rect 65820 22276 65876 22332
rect 65876 22276 65880 22332
rect 65816 22272 65880 22276
rect 65896 22332 65960 22336
rect 65896 22276 65900 22332
rect 65900 22276 65956 22332
rect 65956 22276 65960 22332
rect 65896 22272 65960 22276
rect 15332 22264 15396 22268
rect 15332 22208 15346 22264
rect 15346 22208 15396 22264
rect 15332 22204 15396 22208
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 65656 21244 65720 21248
rect 65656 21188 65660 21244
rect 65660 21188 65716 21244
rect 65716 21188 65720 21244
rect 65656 21184 65720 21188
rect 65736 21244 65800 21248
rect 65736 21188 65740 21244
rect 65740 21188 65796 21244
rect 65796 21188 65800 21244
rect 65736 21184 65800 21188
rect 65816 21244 65880 21248
rect 65816 21188 65820 21244
rect 65820 21188 65876 21244
rect 65876 21188 65880 21244
rect 65816 21184 65880 21188
rect 65896 21244 65960 21248
rect 65896 21188 65900 21244
rect 65900 21188 65956 21244
rect 65956 21188 65960 21244
rect 65896 21184 65960 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 65656 20156 65720 20160
rect 65656 20100 65660 20156
rect 65660 20100 65716 20156
rect 65716 20100 65720 20156
rect 65656 20096 65720 20100
rect 65736 20156 65800 20160
rect 65736 20100 65740 20156
rect 65740 20100 65796 20156
rect 65796 20100 65800 20156
rect 65736 20096 65800 20100
rect 65816 20156 65880 20160
rect 65816 20100 65820 20156
rect 65820 20100 65876 20156
rect 65876 20100 65880 20156
rect 65816 20096 65880 20100
rect 65896 20156 65960 20160
rect 65896 20100 65900 20156
rect 65900 20100 65956 20156
rect 65956 20100 65960 20156
rect 65896 20096 65960 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 65656 19068 65720 19072
rect 65656 19012 65660 19068
rect 65660 19012 65716 19068
rect 65716 19012 65720 19068
rect 65656 19008 65720 19012
rect 65736 19068 65800 19072
rect 65736 19012 65740 19068
rect 65740 19012 65796 19068
rect 65796 19012 65800 19068
rect 65736 19008 65800 19012
rect 65816 19068 65880 19072
rect 65816 19012 65820 19068
rect 65820 19012 65876 19068
rect 65876 19012 65880 19068
rect 65816 19008 65880 19012
rect 65896 19068 65960 19072
rect 65896 19012 65900 19068
rect 65900 19012 65956 19068
rect 65956 19012 65960 19068
rect 65896 19008 65960 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 65656 17980 65720 17984
rect 65656 17924 65660 17980
rect 65660 17924 65716 17980
rect 65716 17924 65720 17980
rect 65656 17920 65720 17924
rect 65736 17980 65800 17984
rect 65736 17924 65740 17980
rect 65740 17924 65796 17980
rect 65796 17924 65800 17980
rect 65736 17920 65800 17924
rect 65816 17980 65880 17984
rect 65816 17924 65820 17980
rect 65820 17924 65876 17980
rect 65876 17924 65880 17980
rect 65816 17920 65880 17924
rect 65896 17980 65960 17984
rect 65896 17924 65900 17980
rect 65900 17924 65956 17980
rect 65956 17924 65960 17980
rect 65896 17920 65960 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 65656 16892 65720 16896
rect 65656 16836 65660 16892
rect 65660 16836 65716 16892
rect 65716 16836 65720 16892
rect 65656 16832 65720 16836
rect 65736 16892 65800 16896
rect 65736 16836 65740 16892
rect 65740 16836 65796 16892
rect 65796 16836 65800 16892
rect 65736 16832 65800 16836
rect 65816 16892 65880 16896
rect 65816 16836 65820 16892
rect 65820 16836 65876 16892
rect 65876 16836 65880 16892
rect 65816 16832 65880 16836
rect 65896 16892 65960 16896
rect 65896 16836 65900 16892
rect 65900 16836 65956 16892
rect 65956 16836 65960 16892
rect 65896 16832 65960 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 65656 15804 65720 15808
rect 65656 15748 65660 15804
rect 65660 15748 65716 15804
rect 65716 15748 65720 15804
rect 65656 15744 65720 15748
rect 65736 15804 65800 15808
rect 65736 15748 65740 15804
rect 65740 15748 65796 15804
rect 65796 15748 65800 15804
rect 65736 15744 65800 15748
rect 65816 15804 65880 15808
rect 65816 15748 65820 15804
rect 65820 15748 65876 15804
rect 65876 15748 65880 15804
rect 65816 15744 65880 15748
rect 65896 15804 65960 15808
rect 65896 15748 65900 15804
rect 65900 15748 65956 15804
rect 65956 15748 65960 15804
rect 65896 15744 65960 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 65656 14716 65720 14720
rect 65656 14660 65660 14716
rect 65660 14660 65716 14716
rect 65716 14660 65720 14716
rect 65656 14656 65720 14660
rect 65736 14716 65800 14720
rect 65736 14660 65740 14716
rect 65740 14660 65796 14716
rect 65796 14660 65800 14716
rect 65736 14656 65800 14660
rect 65816 14716 65880 14720
rect 65816 14660 65820 14716
rect 65820 14660 65876 14716
rect 65876 14660 65880 14716
rect 65816 14656 65880 14660
rect 65896 14716 65960 14720
rect 65896 14660 65900 14716
rect 65900 14660 65956 14716
rect 65956 14660 65960 14716
rect 65896 14656 65960 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 15332 13636 15396 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 65656 13628 65720 13632
rect 65656 13572 65660 13628
rect 65660 13572 65716 13628
rect 65716 13572 65720 13628
rect 65656 13568 65720 13572
rect 65736 13628 65800 13632
rect 65736 13572 65740 13628
rect 65740 13572 65796 13628
rect 65796 13572 65800 13628
rect 65736 13568 65800 13572
rect 65816 13628 65880 13632
rect 65816 13572 65820 13628
rect 65820 13572 65876 13628
rect 65876 13572 65880 13628
rect 65816 13568 65880 13572
rect 65896 13628 65960 13632
rect 65896 13572 65900 13628
rect 65900 13572 65956 13628
rect 65956 13572 65960 13628
rect 65896 13568 65960 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 14228 12608 14292 12612
rect 14228 12552 14242 12608
rect 14242 12552 14292 12608
rect 14228 12548 14292 12552
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 65656 12540 65720 12544
rect 65656 12484 65660 12540
rect 65660 12484 65716 12540
rect 65716 12484 65720 12540
rect 65656 12480 65720 12484
rect 65736 12540 65800 12544
rect 65736 12484 65740 12540
rect 65740 12484 65796 12540
rect 65796 12484 65800 12540
rect 65736 12480 65800 12484
rect 65816 12540 65880 12544
rect 65816 12484 65820 12540
rect 65820 12484 65876 12540
rect 65876 12484 65880 12540
rect 65816 12480 65880 12484
rect 65896 12540 65960 12544
rect 65896 12484 65900 12540
rect 65900 12484 65956 12540
rect 65956 12484 65960 12540
rect 65896 12480 65960 12484
rect 16436 12140 16500 12204
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 65656 11452 65720 11456
rect 65656 11396 65660 11452
rect 65660 11396 65716 11452
rect 65716 11396 65720 11452
rect 65656 11392 65720 11396
rect 65736 11452 65800 11456
rect 65736 11396 65740 11452
rect 65740 11396 65796 11452
rect 65796 11396 65800 11452
rect 65736 11392 65800 11396
rect 65816 11452 65880 11456
rect 65816 11396 65820 11452
rect 65820 11396 65876 11452
rect 65876 11396 65880 11452
rect 65816 11392 65880 11396
rect 65896 11452 65960 11456
rect 65896 11396 65900 11452
rect 65900 11396 65956 11452
rect 65956 11396 65960 11452
rect 65896 11392 65960 11396
rect 20116 11052 20180 11116
rect 17540 10976 17604 10980
rect 17540 10920 17554 10976
rect 17554 10920 17604 10976
rect 17540 10916 17604 10920
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 65656 10364 65720 10368
rect 65656 10308 65660 10364
rect 65660 10308 65716 10364
rect 65716 10308 65720 10364
rect 65656 10304 65720 10308
rect 65736 10364 65800 10368
rect 65736 10308 65740 10364
rect 65740 10308 65796 10364
rect 65796 10308 65800 10364
rect 65736 10304 65800 10308
rect 65816 10364 65880 10368
rect 65816 10308 65820 10364
rect 65820 10308 65876 10364
rect 65876 10308 65880 10364
rect 65816 10304 65880 10308
rect 65896 10364 65960 10368
rect 65896 10308 65900 10364
rect 65900 10308 65956 10364
rect 65956 10308 65960 10364
rect 65896 10304 65960 10308
rect 20300 9828 20364 9892
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 8156 9556 8220 9620
rect 13124 9556 13188 9620
rect 17724 9616 17788 9620
rect 17724 9560 17738 9616
rect 17738 9560 17788 9616
rect 17724 9556 17788 9560
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 65656 9276 65720 9280
rect 65656 9220 65660 9276
rect 65660 9220 65716 9276
rect 65716 9220 65720 9276
rect 65656 9216 65720 9220
rect 65736 9276 65800 9280
rect 65736 9220 65740 9276
rect 65740 9220 65796 9276
rect 65796 9220 65800 9276
rect 65736 9216 65800 9220
rect 65816 9276 65880 9280
rect 65816 9220 65820 9276
rect 65820 9220 65876 9276
rect 65876 9220 65880 9276
rect 65816 9216 65880 9220
rect 65896 9276 65960 9280
rect 65896 9220 65900 9276
rect 65900 9220 65956 9276
rect 65956 9220 65960 9276
rect 65896 9216 65960 9220
rect 16988 9148 17052 9212
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 6868 8332 6932 8396
rect 13676 8332 13740 8396
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 65656 8188 65720 8192
rect 65656 8132 65660 8188
rect 65660 8132 65716 8188
rect 65716 8132 65720 8188
rect 65656 8128 65720 8132
rect 65736 8188 65800 8192
rect 65736 8132 65740 8188
rect 65740 8132 65796 8188
rect 65796 8132 65800 8188
rect 65736 8128 65800 8132
rect 65816 8188 65880 8192
rect 65816 8132 65820 8188
rect 65820 8132 65876 8188
rect 65876 8132 65880 8188
rect 65816 8128 65880 8132
rect 65896 8188 65960 8192
rect 65896 8132 65900 8188
rect 65900 8132 65956 8188
rect 65956 8132 65960 8188
rect 65896 8128 65960 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 65656 7100 65720 7104
rect 65656 7044 65660 7100
rect 65660 7044 65716 7100
rect 65716 7044 65720 7100
rect 65656 7040 65720 7044
rect 65736 7100 65800 7104
rect 65736 7044 65740 7100
rect 65740 7044 65796 7100
rect 65796 7044 65800 7100
rect 65736 7040 65800 7044
rect 65816 7100 65880 7104
rect 65816 7044 65820 7100
rect 65820 7044 65876 7100
rect 65876 7044 65880 7100
rect 65816 7040 65880 7044
rect 65896 7100 65960 7104
rect 65896 7044 65900 7100
rect 65900 7044 65956 7100
rect 65956 7044 65960 7100
rect 65896 7040 65960 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 65656 6012 65720 6016
rect 65656 5956 65660 6012
rect 65660 5956 65716 6012
rect 65716 5956 65720 6012
rect 65656 5952 65720 5956
rect 65736 6012 65800 6016
rect 65736 5956 65740 6012
rect 65740 5956 65796 6012
rect 65796 5956 65800 6012
rect 65736 5952 65800 5956
rect 65816 6012 65880 6016
rect 65816 5956 65820 6012
rect 65820 5956 65876 6012
rect 65876 5956 65880 6012
rect 65816 5952 65880 5956
rect 65896 6012 65960 6016
rect 65896 5956 65900 6012
rect 65900 5956 65956 6012
rect 65956 5956 65960 6012
rect 65896 5952 65960 5956
rect 16436 5612 16500 5676
rect 17908 5612 17972 5676
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 65656 4924 65720 4928
rect 65656 4868 65660 4924
rect 65660 4868 65716 4924
rect 65716 4868 65720 4924
rect 65656 4864 65720 4868
rect 65736 4924 65800 4928
rect 65736 4868 65740 4924
rect 65740 4868 65796 4924
rect 65796 4868 65800 4924
rect 65736 4864 65800 4868
rect 65816 4924 65880 4928
rect 65816 4868 65820 4924
rect 65820 4868 65876 4924
rect 65876 4868 65880 4924
rect 65816 4864 65880 4868
rect 65896 4924 65960 4928
rect 65896 4868 65900 4924
rect 65900 4868 65956 4924
rect 65956 4868 65960 4924
rect 65896 4864 65960 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 6868 3980 6932 4044
rect 13124 3980 13188 4044
rect 13676 4040 13740 4044
rect 13676 3984 13726 4040
rect 13726 3984 13740 4040
rect 13676 3980 13740 3984
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 65656 3836 65720 3840
rect 65656 3780 65660 3836
rect 65660 3780 65716 3836
rect 65716 3780 65720 3836
rect 65656 3776 65720 3780
rect 65736 3836 65800 3840
rect 65736 3780 65740 3836
rect 65740 3780 65796 3836
rect 65796 3780 65800 3836
rect 65736 3776 65800 3780
rect 65816 3836 65880 3840
rect 65816 3780 65820 3836
rect 65820 3780 65876 3836
rect 65876 3780 65880 3836
rect 65816 3776 65880 3780
rect 65896 3836 65960 3840
rect 65896 3780 65900 3836
rect 65900 3780 65956 3836
rect 65956 3780 65960 3836
rect 65896 3776 65960 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 17908 2892 17972 2956
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 65656 2748 65720 2752
rect 65656 2692 65660 2748
rect 65660 2692 65716 2748
rect 65716 2692 65720 2748
rect 65656 2688 65720 2692
rect 65736 2748 65800 2752
rect 65736 2692 65740 2748
rect 65740 2692 65796 2748
rect 65796 2692 65800 2748
rect 65736 2688 65800 2692
rect 65816 2748 65880 2752
rect 65816 2692 65820 2748
rect 65820 2692 65876 2748
rect 65876 2692 65880 2748
rect 65816 2688 65880 2692
rect 65896 2748 65960 2752
rect 65896 2692 65900 2748
rect 65900 2692 65956 2748
rect 65956 2692 65960 2748
rect 65896 2688 65960 2692
rect 8156 2620 8220 2684
rect 20116 2484 20180 2548
rect 20300 2348 20364 2412
rect 16988 2212 17052 2276
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
rect 14228 2076 14292 2140
<< metal4 >>
rect 4208 57152 4528 57712
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 19568 57696 19888 57712
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 17539 26348 17605 26349
rect 17539 26284 17540 26348
rect 17604 26284 17605 26348
rect 17539 26283 17605 26284
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 15331 22268 15397 22269
rect 15331 22204 15332 22268
rect 15396 22204 15397 22268
rect 15331 22203 15397 22204
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 15334 13701 15394 22203
rect 15331 13700 15397 13701
rect 15331 13636 15332 13700
rect 15396 13636 15397 13700
rect 15331 13635 15397 13636
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 14227 12612 14293 12613
rect 14227 12548 14228 12612
rect 14292 12548 14293 12612
rect 14227 12547 14293 12548
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 8155 9620 8221 9621
rect 8155 9556 8156 9620
rect 8220 9556 8221 9620
rect 8155 9555 8221 9556
rect 13123 9620 13189 9621
rect 13123 9556 13124 9620
rect 13188 9556 13189 9620
rect 13123 9555 13189 9556
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 6867 8396 6933 8397
rect 6867 8332 6868 8396
rect 6932 8332 6933 8396
rect 6867 8331 6933 8332
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 6870 4045 6930 8331
rect 6867 4044 6933 4045
rect 6867 3980 6868 4044
rect 6932 3980 6933 4044
rect 6867 3979 6933 3980
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 8158 2685 8218 9555
rect 13126 4045 13186 9555
rect 13675 8396 13741 8397
rect 13675 8332 13676 8396
rect 13740 8332 13741 8396
rect 13675 8331 13741 8332
rect 13678 4045 13738 8331
rect 13123 4044 13189 4045
rect 13123 3980 13124 4044
rect 13188 3980 13189 4044
rect 13123 3979 13189 3980
rect 13675 4044 13741 4045
rect 13675 3980 13676 4044
rect 13740 3980 13741 4044
rect 13675 3979 13741 3980
rect 8155 2684 8221 2685
rect 8155 2620 8156 2684
rect 8220 2620 8221 2684
rect 8155 2619 8221 2620
rect 14230 2141 14290 12547
rect 16435 12204 16501 12205
rect 16435 12140 16436 12204
rect 16500 12140 16501 12204
rect 16435 12139 16501 12140
rect 16438 5677 16498 12139
rect 17542 10981 17602 26283
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 17723 24988 17789 24989
rect 17723 24924 17724 24988
rect 17788 24924 17789 24988
rect 17723 24923 17789 24924
rect 17539 10980 17605 10981
rect 17539 10916 17540 10980
rect 17604 10916 17605 10980
rect 17539 10915 17605 10916
rect 17726 9621 17786 24923
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 34928 57152 35248 57712
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 20115 11116 20181 11117
rect 20115 11052 20116 11116
rect 20180 11052 20181 11116
rect 20115 11051 20181 11052
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 17723 9620 17789 9621
rect 17723 9556 17724 9620
rect 17788 9556 17789 9620
rect 17723 9555 17789 9556
rect 16987 9212 17053 9213
rect 16987 9148 16988 9212
rect 17052 9148 17053 9212
rect 16987 9147 17053 9148
rect 16435 5676 16501 5677
rect 16435 5612 16436 5676
rect 16500 5612 16501 5676
rect 16435 5611 16501 5612
rect 16990 2277 17050 9147
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 17907 5676 17973 5677
rect 17907 5612 17908 5676
rect 17972 5612 17973 5676
rect 17907 5611 17973 5612
rect 17910 2957 17970 5611
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 17907 2956 17973 2957
rect 17907 2892 17908 2956
rect 17972 2892 17973 2956
rect 17907 2891 17973 2892
rect 16987 2276 17053 2277
rect 16987 2212 16988 2276
rect 17052 2212 17053 2276
rect 16987 2211 17053 2212
rect 19568 2208 19888 3232
rect 20118 2549 20178 11051
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 20299 9892 20365 9893
rect 20299 9828 20300 9892
rect 20364 9828 20365 9892
rect 20299 9827 20365 9828
rect 20115 2548 20181 2549
rect 20115 2484 20116 2548
rect 20180 2484 20181 2548
rect 20115 2483 20181 2484
rect 20302 2413 20362 9827
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 20299 2412 20365 2413
rect 20299 2348 20300 2412
rect 20364 2348 20365 2412
rect 20299 2347 20365 2348
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 14227 2140 14293 2141
rect 14227 2076 14228 2140
rect 14292 2076 14293 2140
rect 19568 2128 19888 2144
rect 34928 2128 35248 2688
rect 50288 57696 50608 57712
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
rect 65648 57152 65968 57712
rect 65648 57088 65656 57152
rect 65720 57088 65736 57152
rect 65800 57088 65816 57152
rect 65880 57088 65896 57152
rect 65960 57088 65968 57152
rect 65648 56064 65968 57088
rect 65648 56000 65656 56064
rect 65720 56000 65736 56064
rect 65800 56000 65816 56064
rect 65880 56000 65896 56064
rect 65960 56000 65968 56064
rect 65648 54976 65968 56000
rect 65648 54912 65656 54976
rect 65720 54912 65736 54976
rect 65800 54912 65816 54976
rect 65880 54912 65896 54976
rect 65960 54912 65968 54976
rect 65648 53888 65968 54912
rect 65648 53824 65656 53888
rect 65720 53824 65736 53888
rect 65800 53824 65816 53888
rect 65880 53824 65896 53888
rect 65960 53824 65968 53888
rect 65648 52800 65968 53824
rect 65648 52736 65656 52800
rect 65720 52736 65736 52800
rect 65800 52736 65816 52800
rect 65880 52736 65896 52800
rect 65960 52736 65968 52800
rect 65648 51712 65968 52736
rect 65648 51648 65656 51712
rect 65720 51648 65736 51712
rect 65800 51648 65816 51712
rect 65880 51648 65896 51712
rect 65960 51648 65968 51712
rect 65648 50624 65968 51648
rect 65648 50560 65656 50624
rect 65720 50560 65736 50624
rect 65800 50560 65816 50624
rect 65880 50560 65896 50624
rect 65960 50560 65968 50624
rect 65648 49536 65968 50560
rect 65648 49472 65656 49536
rect 65720 49472 65736 49536
rect 65800 49472 65816 49536
rect 65880 49472 65896 49536
rect 65960 49472 65968 49536
rect 65648 48448 65968 49472
rect 65648 48384 65656 48448
rect 65720 48384 65736 48448
rect 65800 48384 65816 48448
rect 65880 48384 65896 48448
rect 65960 48384 65968 48448
rect 65648 47360 65968 48384
rect 65648 47296 65656 47360
rect 65720 47296 65736 47360
rect 65800 47296 65816 47360
rect 65880 47296 65896 47360
rect 65960 47296 65968 47360
rect 65648 46272 65968 47296
rect 65648 46208 65656 46272
rect 65720 46208 65736 46272
rect 65800 46208 65816 46272
rect 65880 46208 65896 46272
rect 65960 46208 65968 46272
rect 65648 45184 65968 46208
rect 65648 45120 65656 45184
rect 65720 45120 65736 45184
rect 65800 45120 65816 45184
rect 65880 45120 65896 45184
rect 65960 45120 65968 45184
rect 65648 44096 65968 45120
rect 65648 44032 65656 44096
rect 65720 44032 65736 44096
rect 65800 44032 65816 44096
rect 65880 44032 65896 44096
rect 65960 44032 65968 44096
rect 65648 43008 65968 44032
rect 65648 42944 65656 43008
rect 65720 42944 65736 43008
rect 65800 42944 65816 43008
rect 65880 42944 65896 43008
rect 65960 42944 65968 43008
rect 65648 41920 65968 42944
rect 65648 41856 65656 41920
rect 65720 41856 65736 41920
rect 65800 41856 65816 41920
rect 65880 41856 65896 41920
rect 65960 41856 65968 41920
rect 65648 40832 65968 41856
rect 65648 40768 65656 40832
rect 65720 40768 65736 40832
rect 65800 40768 65816 40832
rect 65880 40768 65896 40832
rect 65960 40768 65968 40832
rect 65648 39744 65968 40768
rect 65648 39680 65656 39744
rect 65720 39680 65736 39744
rect 65800 39680 65816 39744
rect 65880 39680 65896 39744
rect 65960 39680 65968 39744
rect 65648 38656 65968 39680
rect 65648 38592 65656 38656
rect 65720 38592 65736 38656
rect 65800 38592 65816 38656
rect 65880 38592 65896 38656
rect 65960 38592 65968 38656
rect 65648 37568 65968 38592
rect 65648 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65968 37568
rect 65648 36480 65968 37504
rect 65648 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65968 36480
rect 65648 35392 65968 36416
rect 65648 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65968 35392
rect 65648 34304 65968 35328
rect 65648 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65968 34304
rect 65648 33216 65968 34240
rect 65648 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65968 33216
rect 65648 32128 65968 33152
rect 65648 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65968 32128
rect 65648 31040 65968 32064
rect 65648 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65968 31040
rect 65648 29952 65968 30976
rect 65648 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65968 29952
rect 65648 28864 65968 29888
rect 65648 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65968 28864
rect 65648 27776 65968 28800
rect 65648 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65968 27776
rect 65648 26688 65968 27712
rect 65648 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65968 26688
rect 65648 25600 65968 26624
rect 65648 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65968 25600
rect 65648 24512 65968 25536
rect 65648 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65968 24512
rect 65648 23424 65968 24448
rect 65648 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65968 23424
rect 65648 22336 65968 23360
rect 65648 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65968 22336
rect 65648 21248 65968 22272
rect 65648 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65968 21248
rect 65648 20160 65968 21184
rect 65648 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65968 20160
rect 65648 19072 65968 20096
rect 65648 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65968 19072
rect 65648 17984 65968 19008
rect 65648 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65968 17984
rect 65648 16896 65968 17920
rect 65648 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65968 16896
rect 65648 15808 65968 16832
rect 65648 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65968 15808
rect 65648 14720 65968 15744
rect 65648 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65968 14720
rect 65648 13632 65968 14656
rect 65648 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65968 13632
rect 65648 12544 65968 13568
rect 65648 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65968 12544
rect 65648 11456 65968 12480
rect 65648 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65968 11456
rect 65648 10368 65968 11392
rect 65648 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65968 10368
rect 65648 9280 65968 10304
rect 65648 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65968 9280
rect 65648 8192 65968 9216
rect 65648 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65968 8192
rect 65648 7104 65968 8128
rect 65648 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65968 7104
rect 65648 6016 65968 7040
rect 65648 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65968 6016
rect 65648 4928 65968 5952
rect 65648 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65968 4928
rect 65648 3840 65968 4864
rect 65648 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65968 3840
rect 65648 2752 65968 3776
rect 65648 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65968 2752
rect 65648 2128 65968 2688
rect 14227 2075 14293 2076
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__A0 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__A
timestamp 1649977179
transform -1 0 3312 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__A0
timestamp 1649977179
transform -1 0 2208 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__A0
timestamp 1649977179
transform 1 0 2852 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__A0
timestamp 1649977179
transform 1 0 5612 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__A0
timestamp 1649977179
transform -1 0 1748 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__A0
timestamp 1649977179
transform -1 0 1564 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__A
timestamp 1649977179
transform 1 0 6716 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__A0
timestamp 1649977179
transform 1 0 19228 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__A0
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__A0
timestamp 1649977179
transform 1 0 16008 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__A0
timestamp 1649977179
transform -1 0 3312 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__A0
timestamp 1649977179
transform 1 0 8832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__A
timestamp 1649977179
transform 1 0 5888 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0842__A
timestamp 1649977179
transform 1 0 8004 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0846__B
timestamp 1649977179
transform 1 0 7728 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0848__A
timestamp 1649977179
transform -1 0 5060 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0848__B
timestamp 1649977179
transform 1 0 5612 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__A
timestamp 1649977179
transform -1 0 3956 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__A1
timestamp 1649977179
transform 1 0 3496 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__A
timestamp 1649977179
transform -1 0 4140 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__A1
timestamp 1649977179
transform 1 0 3128 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__A
timestamp 1649977179
transform 1 0 1932 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__A1
timestamp 1649977179
transform -1 0 1564 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__A
timestamp 1649977179
transform 1 0 9384 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__A
timestamp 1649977179
transform 1 0 3128 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__A1
timestamp 1649977179
transform 1 0 2944 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__A
timestamp 1649977179
transform -1 0 6256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__A
timestamp 1649977179
transform 1 0 4324 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__A1
timestamp 1649977179
transform -1 0 3956 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__A
timestamp 1649977179
transform -1 0 11960 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__A1
timestamp 1649977179
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0875__A
timestamp 1649977179
transform -1 0 12052 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__A1
timestamp 1649977179
transform 1 0 4140 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__A
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0880__A1
timestamp 1649977179
transform 1 0 3036 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0881__A
timestamp 1649977179
transform 1 0 5152 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0883__A1
timestamp 1649977179
transform 1 0 2484 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0884__A
timestamp 1649977179
transform 1 0 9752 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__A
timestamp 1649977179
transform 1 0 2944 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__A
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__A1
timestamp 1649977179
transform 1 0 2576 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__A1
timestamp 1649977179
transform 1 0 2944 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__A1
timestamp 1649977179
transform 1 0 1564 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0905__A
timestamp 1649977179
transform 1 0 2852 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__A1
timestamp 1649977179
transform 1 0 2852 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__A1
timestamp 1649977179
transform -1 0 2852 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__A1
timestamp 1649977179
transform -1 0 3312 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__A1
timestamp 1649977179
transform 1 0 2944 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__A1
timestamp 1649977179
transform -1 0 2944 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__A
timestamp 1649977179
transform -1 0 6624 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__A1
timestamp 1649977179
transform 1 0 3036 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__A
timestamp 1649977179
transform -1 0 5796 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0932__A1
timestamp 1649977179
transform -1 0 3312 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__A1
timestamp 1649977179
transform 1 0 3128 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__A1
timestamp 1649977179
transform -1 0 4784 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0941__A1
timestamp 1649977179
transform -1 0 5888 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__A1
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__A1
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0949__A1
timestamp 1649977179
transform 1 0 5704 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__A1
timestamp 1649977179
transform 1 0 9476 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__C1
timestamp 1649977179
transform -1 0 4692 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__A1
timestamp 1649977179
transform -1 0 7268 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__C1
timestamp 1649977179
transform 1 0 5060 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__C1
timestamp 1649977179
transform 1 0 8280 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__A
timestamp 1649977179
transform 1 0 15548 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__B
timestamp 1649977179
transform -1 0 7176 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__A
timestamp 1649977179
transform 1 0 5704 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__B
timestamp 1649977179
transform 1 0 8832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__A1
timestamp 1649977179
transform 1 0 6900 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__C1
timestamp 1649977179
transform 1 0 7084 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__A1
timestamp 1649977179
transform 1 0 6256 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__C1
timestamp 1649977179
transform -1 0 6256 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__A1
timestamp 1649977179
transform 1 0 9384 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__A1
timestamp 1649977179
transform 1 0 7636 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A1
timestamp 1649977179
transform -1 0 7360 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__A1
timestamp 1649977179
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__A1
timestamp 1649977179
transform -1 0 9936 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__A1
timestamp 1649977179
transform 1 0 9292 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__A1
timestamp 1649977179
transform 1 0 9936 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__B
timestamp 1649977179
transform -1 0 5428 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__A
timestamp 1649977179
transform 1 0 8280 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__B
timestamp 1649977179
transform 1 0 10120 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__A1
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__A
timestamp 1649977179
transform 1 0 14260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__A
timestamp 1649977179
transform 1 0 13064 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__A1
timestamp 1649977179
transform 1 0 9016 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1003__A1
timestamp 1649977179
transform 1 0 11132 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__A1
timestamp 1649977179
transform -1 0 9752 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__A1
timestamp 1649977179
transform 1 0 11316 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__A
timestamp 1649977179
transform 1 0 13432 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__A1
timestamp 1649977179
transform 1 0 11316 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__A1
timestamp 1649977179
transform -1 0 14628 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1018__A1
timestamp 1649977179
transform 1 0 13340 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__A1
timestamp 1649977179
transform -1 0 12696 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__A
timestamp 1649977179
transform -1 0 23092 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__A
timestamp 1649977179
transform 1 0 21896 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__A
timestamp 1649977179
transform 1 0 23736 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__A
timestamp 1649977179
transform -1 0 23000 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__A
timestamp 1649977179
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__A1
timestamp 1649977179
transform 1 0 24472 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__A
timestamp 1649977179
transform 1 0 22448 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__A1
timestamp 1649977179
transform -1 0 24840 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__A
timestamp 1649977179
transform 1 0 25208 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__A1
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__A
timestamp 1649977179
transform 1 0 23736 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__A1
timestamp 1649977179
transform -1 0 25944 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__A
timestamp 1649977179
transform 1 0 20516 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__A1
timestamp 1649977179
transform 1 0 26128 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__A
timestamp 1649977179
transform 1 0 23184 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__A
timestamp 1649977179
transform -1 0 23920 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__A1
timestamp 1649977179
transform 1 0 28888 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__A
timestamp 1649977179
transform -1 0 28796 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__A1
timestamp 1649977179
transform 1 0 30912 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__A
timestamp 1649977179
transform -1 0 27784 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__A1
timestamp 1649977179
transform 1 0 28888 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__A
timestamp 1649977179
transform 1 0 23736 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__A1
timestamp 1649977179
transform 1 0 26312 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__A
timestamp 1649977179
transform 1 0 25208 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1063__A1
timestamp 1649977179
transform 1 0 26220 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__A
timestamp 1649977179
transform 1 0 20148 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__A
timestamp 1649977179
transform -1 0 27140 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__A1
timestamp 1649977179
transform -1 0 23184 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__C1
timestamp 1649977179
transform -1 0 23736 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__A
timestamp 1649977179
transform 1 0 28244 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__A
timestamp 1649977179
transform 1 0 27692 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1076__A1
timestamp 1649977179
transform 1 0 36156 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1076__C1
timestamp 1649977179
transform 1 0 34040 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__A1
timestamp 1649977179
transform -1 0 34224 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__C1
timestamp 1649977179
transform -1 0 36248 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1080__A1
timestamp 1649977179
transform -1 0 32568 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1080__C1
timestamp 1649977179
transform -1 0 32016 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__A1
timestamp 1649977179
transform 1 0 34960 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__C1
timestamp 1649977179
transform -1 0 36432 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__A
timestamp 1649977179
transform 1 0 30360 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__A1
timestamp 1649977179
transform 1 0 34684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__A1
timestamp 1649977179
transform -1 0 26404 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__A1
timestamp 1649977179
transform -1 0 26496 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__A1
timestamp 1649977179
transform 1 0 25852 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__A1
timestamp 1649977179
transform 1 0 26128 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__A1
timestamp 1649977179
transform 1 0 28888 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__A1
timestamp 1649977179
transform -1 0 30544 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__A
timestamp 1649977179
transform -1 0 34224 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__A
timestamp 1649977179
transform -1 0 36340 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1107__A
timestamp 1649977179
transform -1 0 34684 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__A1
timestamp 1649977179
transform 1 0 37812 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__A1
timestamp 1649977179
transform 1 0 36616 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__A1
timestamp 1649977179
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__A1
timestamp 1649977179
transform -1 0 38180 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__A1
timestamp 1649977179
transform -1 0 38732 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__A1
timestamp 1649977179
transform -1 0 38364 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__A1
timestamp 1649977179
transform 1 0 36524 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__A1
timestamp 1649977179
transform 1 0 35972 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__A1
timestamp 1649977179
transform -1 0 32476 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1132__A1
timestamp 1649977179
transform -1 0 33948 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__A1
timestamp 1649977179
transform -1 0 32752 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__A
timestamp 1649977179
transform 1 0 34776 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__A
timestamp 1649977179
transform -1 0 34408 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__A
timestamp 1649977179
transform 1 0 34040 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__A1
timestamp 1649977179
transform 1 0 34776 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__A1
timestamp 1649977179
transform 1 0 34868 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__A1
timestamp 1649977179
transform 1 0 37260 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__A1
timestamp 1649977179
transform -1 0 38916 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1151__A1
timestamp 1649977179
transform -1 0 37444 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__A1
timestamp 1649977179
transform 1 0 37352 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__A1
timestamp 1649977179
transform -1 0 39192 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__A
timestamp 1649977179
transform -1 0 32292 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1161__A1
timestamp 1649977179
transform -1 0 35236 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__A1
timestamp 1649977179
transform -1 0 34868 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1165__A1
timestamp 1649977179
transform 1 0 33028 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__A1
timestamp 1649977179
transform 1 0 32660 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__A
timestamp 1649977179
transform -1 0 28428 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1172__A
timestamp 1649977179
transform 1 0 30268 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__A1
timestamp 1649977179
transform 1 0 34776 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__A1
timestamp 1649977179
transform 1 0 37352 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__A1
timestamp 1649977179
transform -1 0 40020 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__A1
timestamp 1649977179
transform 1 0 37260 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__A1
timestamp 1649977179
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__A1
timestamp 1649977179
transform 1 0 33672 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__A1
timestamp 1649977179
transform 1 0 31924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1193__A1
timestamp 1649977179
transform 1 0 32660 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__A1
timestamp 1649977179
transform 1 0 32936 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__A1
timestamp 1649977179
transform 1 0 30636 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1199__A1
timestamp 1649977179
transform 1 0 32016 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__A
timestamp 1649977179
transform -1 0 20608 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__A
timestamp 1649977179
transform 1 0 17572 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__A
timestamp 1649977179
transform 1 0 20332 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__A
timestamp 1649977179
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__A1
timestamp 1649977179
transform 1 0 23644 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__A
timestamp 1649977179
transform 1 0 24656 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__A1
timestamp 1649977179
transform 1 0 24472 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__A
timestamp 1649977179
transform -1 0 25116 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__A1
timestamp 1649977179
transform 1 0 26220 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1220__A
timestamp 1649977179
transform 1 0 16468 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__A1
timestamp 1649977179
transform 1 0 23092 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1223__A
timestamp 1649977179
transform 1 0 14996 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__A1
timestamp 1649977179
transform 1 0 19872 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1229__A
timestamp 1649977179
transform -1 0 12972 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1231__A1
timestamp 1649977179
transform 1 0 19044 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1232__A
timestamp 1649977179
transform 1 0 14812 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1234__A1
timestamp 1649977179
transform 1 0 17020 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1235__A
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1237__A1
timestamp 1649977179
transform 1 0 16192 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__A
timestamp 1649977179
transform 1 0 14168 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1240__A1
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1241__A
timestamp 1649977179
transform -1 0 16560 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1243__A
timestamp 1649977179
transform 1 0 20516 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1245__A1
timestamp 1649977179
transform 1 0 23736 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1252__A
timestamp 1649977179
transform 1 0 28520 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__A1
timestamp 1649977179
transform 1 0 30360 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__A1
timestamp 1649977179
transform 1 0 29808 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1261__A1
timestamp 1649977179
transform 1 0 30544 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__A1
timestamp 1649977179
transform 1 0 30360 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__A1
timestamp 1649977179
transform -1 0 31004 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__A1
timestamp 1649977179
transform -1 0 32384 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__A1
timestamp 1649977179
transform 1 0 27784 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__A1
timestamp 1649977179
transform 1 0 26220 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1277__A1
timestamp 1649977179
transform 1 0 26312 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1279__A1
timestamp 1649977179
transform 1 0 27508 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1284__A
timestamp 1649977179
transform 1 0 18032 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1289__A1
timestamp 1649977179
transform -1 0 22632 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__A1
timestamp 1649977179
transform 1 0 24564 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1294__A1
timestamp 1649977179
transform 1 0 21436 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1296__A1
timestamp 1649977179
transform 1 0 21160 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1300__A1
timestamp 1649977179
transform 1 0 22908 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1302__A1
timestamp 1649977179
transform 1 0 20424 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1304__A1
timestamp 1649977179
transform 1 0 18584 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1307__A1
timestamp 1649977179
transform 1 0 18676 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__A1
timestamp 1649977179
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1311__A1
timestamp 1649977179
transform -1 0 18768 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1316__A
timestamp 1649977179
transform -1 0 16100 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1321__A1
timestamp 1649977179
transform -1 0 19412 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1324__A
timestamp 1649977179
transform -1 0 13616 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1325__A1
timestamp 1649977179
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1327__A1
timestamp 1649977179
transform 1 0 14260 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1329__A1
timestamp 1649977179
transform -1 0 14260 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1333__A1
timestamp 1649977179
transform 1 0 15916 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1335__A1
timestamp 1649977179
transform -1 0 13708 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1337__A
timestamp 1649977179
transform -1 0 21988 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1338__A1
timestamp 1649977179
transform -1 0 13800 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1340__A1
timestamp 1649977179
transform 1 0 15916 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1342__A1
timestamp 1649977179
transform -1 0 13616 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1344__A1
timestamp 1649977179
transform -1 0 18032 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1349__A
timestamp 1649977179
transform 1 0 20424 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__A
timestamp 1649977179
transform 1 0 21160 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1355__A1
timestamp 1649977179
transform 1 0 27048 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1357__A1
timestamp 1649977179
transform 1 0 26312 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1359__A1
timestamp 1649977179
transform 1 0 26312 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1361__A1
timestamp 1649977179
transform 1 0 26220 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1365__A1
timestamp 1649977179
transform 1 0 21160 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1367__A
timestamp 1649977179
transform 1 0 17204 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1368__A1
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1370__A1
timestamp 1649977179
transform 1 0 17848 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1372__A1
timestamp 1649977179
transform 1 0 15916 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1374__A1
timestamp 1649977179
transform 1 0 17480 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1376__A1
timestamp 1649977179
transform 1 0 22172 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1380__A
timestamp 1649977179
transform -1 0 22632 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1382__A
timestamp 1649977179
transform 1 0 20792 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1385__A
timestamp 1649977179
transform 1 0 17204 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1386__A1
timestamp 1649977179
transform 1 0 17020 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1388__A1
timestamp 1649977179
transform 1 0 18584 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1390__A1
timestamp 1649977179
transform 1 0 19228 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1392__A1
timestamp 1649977179
transform 1 0 21344 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1394__A1
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1398__A
timestamp 1649977179
transform -1 0 20148 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1399__A1
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1401__A1
timestamp 1649977179
transform 1 0 26312 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1403__A1
timestamp 1649977179
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1405__A1
timestamp 1649977179
transform 1 0 21160 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1407__A1
timestamp 1649977179
transform 1 0 22724 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1409__A
timestamp 1649977179
transform 1 0 10948 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1410__A1
timestamp 1649977179
transform 1 0 19320 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1427__A2
timestamp 1649977179
transform 1 0 16468 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1428__A2
timestamp 1649977179
transform 1 0 18400 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1429__A2
timestamp 1649977179
transform 1 0 22724 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1438__A2
timestamp 1649977179
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1439__A2
timestamp 1649977179
transform -1 0 20516 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1440__A2
timestamp 1649977179
transform -1 0 24564 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1453__D
timestamp 1649977179
transform -1 0 26864 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1454__A2
timestamp 1649977179
transform 1 0 14812 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1455__A2
timestamp 1649977179
transform 1 0 17848 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1456__A2
timestamp 1649977179
transform 1 0 24288 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1458__B
timestamp 1649977179
transform -1 0 25116 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1460__A
timestamp 1649977179
transform -1 0 15180 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1462__A
timestamp 1649977179
transform -1 0 37260 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1463__A
timestamp 1649977179
transform 1 0 35236 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1473__D
timestamp 1649977179
transform -1 0 28980 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1477__A2
timestamp 1649977179
transform 1 0 17848 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1482__B
timestamp 1649977179
transform -1 0 18124 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1491__A
timestamp 1649977179
transform -1 0 16376 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1506__D
timestamp 1649977179
transform -1 0 29716 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1519__D
timestamp 1649977179
transform -1 0 28888 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1540__A2
timestamp 1649977179
transform 1 0 31464 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1540__B1
timestamp 1649977179
transform 1 0 31832 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1552__A2
timestamp 1649977179
transform 1 0 33304 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1552__B1
timestamp 1649977179
transform 1 0 33948 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1558__A2
timestamp 1649977179
transform 1 0 14352 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1564__A2
timestamp 1649977179
transform 1 0 30268 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1564__B1
timestamp 1649977179
transform 1 0 30452 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1570__A2
timestamp 1649977179
transform -1 0 17572 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1578__A
timestamp 1649977179
transform 1 0 3128 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_wb_clk_i_A
timestamp 1649977179
transform -1 0 21528 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0__f_wb_clk_i_A
timestamp 1649977179
transform 1 0 12052 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1__f_wb_clk_i_A
timestamp 1649977179
transform -1 0 29716 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_1_wb_clk_i_A
timestamp 1649977179
transform 1 0 14168 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_2_wb_clk_i_A
timestamp 1649977179
transform 1 0 11224 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_3_wb_clk_i_A
timestamp 1649977179
transform -1 0 4048 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_4_wb_clk_i_A
timestamp 1649977179
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_5_wb_clk_i_A
timestamp 1649977179
transform 1 0 9752 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_6_wb_clk_i_A
timestamp 1649977179
transform 1 0 14260 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_7_wb_clk_i_A
timestamp 1649977179
transform 1 0 18124 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_8_wb_clk_i_A
timestamp 1649977179
transform 1 0 27784 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_9_wb_clk_i_A
timestamp 1649977179
transform 1 0 29532 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_10_wb_clk_i_A
timestamp 1649977179
transform 1 0 35788 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_11_wb_clk_i_A
timestamp 1649977179
transform 1 0 35788 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_12_wb_clk_i_A
timestamp 1649977179
transform 1 0 31464 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_13_wb_clk_i_A
timestamp 1649977179
transform 1 0 28796 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_14_wb_clk_i_A
timestamp 1649977179
transform 1 0 34040 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_15_wb_clk_i_A
timestamp 1649977179
transform 1 0 39192 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_16_wb_clk_i_A
timestamp 1649977179
transform 1 0 39008 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_17_wb_clk_i_A
timestamp 1649977179
transform 1 0 31832 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_18_wb_clk_i_A
timestamp 1649977179
transform 1 0 27048 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_19_wb_clk_i_A
timestamp 1649977179
transform 1 0 27968 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_20_wb_clk_i_A
timestamp 1649977179
transform 1 0 17572 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_21_wb_clk_i_A
timestamp 1649977179
transform 1 0 16836 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_22_wb_clk_i_A
timestamp 1649977179
transform 1 0 5336 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_23_wb_clk_i_A
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_24_wb_clk_i_A
timestamp 1649977179
transform 1 0 8924 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 4784 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 4416 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 1840 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 19412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 4784 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 21988 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 20700 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 2760 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 4968 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 4416 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 9752 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 7636 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 1656 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 3864 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 15364 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 15548 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 11684 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 8464 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 13616 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 12788 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 14812 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 24564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 27140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 19964 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 19412 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 11684 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 2760 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 1656 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10
timestamp 1649977179
transform 1 0 2024 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17
timestamp 1649977179
transform 1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1649977179
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4140 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37
timestamp 1649977179
transform 1 0 4508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44
timestamp 1649977179
transform 1 0 5152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1649977179
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64
timestamp 1649977179
transform 1 0 6992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72
timestamp 1649977179
transform 1 0 7728 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1649977179
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_88
timestamp 1649977179
transform 1 0 9200 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_98
timestamp 1649977179
transform 1 0 10120 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1649977179
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_123
timestamp 1649977179
transform 1 0 12420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_133 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1649977179
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_151 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14996 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_163
timestamp 1649977179
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1649977179
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_173
timestamp 1649977179
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_189
timestamp 1649977179
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1649977179
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_199
timestamp 1649977179
transform 1 0 19412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_206
timestamp 1649977179
transform 1 0 20056 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_213
timestamp 1649977179
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1649977179
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_227
timestamp 1649977179
transform 1 0 21988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_234
timestamp 1649977179
transform 1 0 22632 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_241
timestamp 1649977179
transform 1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_248
timestamp 1649977179
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_255
timestamp 1649977179
transform 1 0 24564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_262
timestamp 1649977179
transform 1 0 25208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_269
timestamp 1649977179
transform 1 0 25852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1649977179
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_283
timestamp 1649977179
transform 1 0 27140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_290
timestamp 1649977179
transform 1 0 27784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_297
timestamp 1649977179
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1649977179
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_309
timestamp 1649977179
transform 1 0 29532 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_318
timestamp 1649977179
transform 1 0 30360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_325
timestamp 1649977179
transform 1 0 31004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_332
timestamp 1649977179
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_337
timestamp 1649977179
transform 1 0 32108 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_346
timestamp 1649977179
transform 1 0 32936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_353
timestamp 1649977179
transform 1 0 33580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_360
timestamp 1649977179
transform 1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_368
timestamp 1649977179
transform 1 0 34960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_375
timestamp 1649977179
transform 1 0 35604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_382
timestamp 1649977179
transform 1 0 36248 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_396
timestamp 1649977179
transform 1 0 37536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1649977179
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_410
timestamp 1649977179
transform 1 0 38824 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_418
timestamp 1649977179
transform 1 0 39560 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_424
timestamp 1649977179
transform 1 0 40112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_431
timestamp 1649977179
transform 1 0 40756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_438
timestamp 1649977179
transform 1 0 41400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_446
timestamp 1649977179
transform 1 0 42136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_452
timestamp 1649977179
transform 1 0 42688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_459
timestamp 1649977179
transform 1 0 43332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_466
timestamp 1649977179
transform 1 0 43976 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_474
timestamp 1649977179
transform 1 0 44712 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_480
timestamp 1649977179
transform 1 0 45264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_487
timestamp 1649977179
transform 1 0 45908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_494
timestamp 1649977179
transform 1 0 46552 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_502
timestamp 1649977179
transform 1 0 47288 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_508
timestamp 1649977179
transform 1 0 47840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_515
timestamp 1649977179
transform 1 0 48484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_522
timestamp 1649977179
transform 1 0 49128 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_530
timestamp 1649977179
transform 1 0 49864 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_536
timestamp 1649977179
transform 1 0 50416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_543
timestamp 1649977179
transform 1 0 51060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_550
timestamp 1649977179
transform 1 0 51704 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_558
timestamp 1649977179
transform 1 0 52440 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_564
timestamp 1649977179
transform 1 0 52992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_571
timestamp 1649977179
transform 1 0 53636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_578
timestamp 1649977179
transform 1 0 54280 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_586
timestamp 1649977179
transform 1 0 55016 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_592
timestamp 1649977179
transform 1 0 55568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_599
timestamp 1649977179
transform 1 0 56212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_606
timestamp 1649977179
transform 1 0 56856 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_614
timestamp 1649977179
transform 1 0 57592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_620
timestamp 1649977179
transform 1 0 58144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_627
timestamp 1649977179
transform 1 0 58788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_634
timestamp 1649977179
transform 1 0 59432 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_642
timestamp 1649977179
transform 1 0 60168 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_648
timestamp 1649977179
transform 1 0 60720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_655
timestamp 1649977179
transform 1 0 61364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_662
timestamp 1649977179
transform 1 0 62008 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_670
timestamp 1649977179
transform 1 0 62744 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_676
timestamp 1649977179
transform 1 0 63296 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_683 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 63940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_695
timestamp 1649977179
transform 1 0 65044 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_699
timestamp 1649977179
transform 1 0 65412 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_701
timestamp 1649977179
transform 1 0 65596 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_713
timestamp 1649977179
transform 1 0 66700 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_717
timestamp 1649977179
transform 1 0 67068 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_724
timestamp 1649977179
transform 1 0 67712 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_729
timestamp 1649977179
transform 1 0 68172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_10
timestamp 1649977179
transform 1 0 2024 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_32
timestamp 1649977179
transform 1 0 4048 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1649977179
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_73
timestamp 1649977179
transform 1 0 7820 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_79
timestamp 1649977179
transform 1 0 8372 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_96
timestamp 1649977179
transform 1 0 9936 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1649977179
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_126
timestamp 1649977179
transform 1 0 12696 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_138
timestamp 1649977179
transform 1 0 13800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_152
timestamp 1649977179
transform 1 0 15088 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_160
timestamp 1649977179
transform 1 0 15824 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_173
timestamp 1649977179
transform 1 0 17020 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_192
timestamp 1649977179
transform 1 0 18768 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_199
timestamp 1649977179
transform 1 0 19412 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_206
timestamp 1649977179
transform 1 0 20056 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_213
timestamp 1649977179
transform 1 0 20700 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1649977179
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_227
timestamp 1649977179
transform 1 0 21988 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_234
timestamp 1649977179
transform 1 0 22632 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_241
timestamp 1649977179
transform 1 0 23276 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_248
timestamp 1649977179
transform 1 0 23920 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_255
timestamp 1649977179
transform 1 0 24564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_262
timestamp 1649977179
transform 1 0 25208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_269
timestamp 1649977179
transform 1 0 25852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1649977179
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_283
timestamp 1649977179
transform 1 0 27140 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_290
timestamp 1649977179
transform 1 0 27784 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_297
timestamp 1649977179
transform 1 0 28428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_304
timestamp 1649977179
transform 1 0 29072 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_311
timestamp 1649977179
transform 1 0 29716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_318
timestamp 1649977179
transform 1 0 30360 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_325
timestamp 1649977179
transform 1 0 31004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_332
timestamp 1649977179
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_337
timestamp 1649977179
transform 1 0 32108 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_346
timestamp 1649977179
transform 1 0 32936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_353
timestamp 1649977179
transform 1 0 33580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_360
timestamp 1649977179
transform 1 0 34224 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_367
timestamp 1649977179
transform 1 0 34868 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_376
timestamp 1649977179
transform 1 0 35696 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1649977179
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1649977179
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_396
timestamp 1649977179
transform 1 0 37536 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_403
timestamp 1649977179
transform 1 0 38180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_410
timestamp 1649977179
transform 1 0 38824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_417
timestamp 1649977179
transform 1 0 39468 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_424
timestamp 1649977179
transform 1 0 40112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_431
timestamp 1649977179
transform 1 0 40756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_438
timestamp 1649977179
transform 1 0 41400 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_446
timestamp 1649977179
transform 1 0 42136 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_452
timestamp 1649977179
transform 1 0 42688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_459
timestamp 1649977179
transform 1 0 43332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_466
timestamp 1649977179
transform 1 0 43976 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_473
timestamp 1649977179
transform 1 0 44620 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_480
timestamp 1649977179
transform 1 0 45264 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_487
timestamp 1649977179
transform 1 0 45908 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_494
timestamp 1649977179
transform 1 0 46552 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_502
timestamp 1649977179
transform 1 0 47288 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_508
timestamp 1649977179
transform 1 0 47840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_515
timestamp 1649977179
transform 1 0 48484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_522
timestamp 1649977179
transform 1 0 49128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_529
timestamp 1649977179
transform 1 0 49772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_536
timestamp 1649977179
transform 1 0 50416 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_543
timestamp 1649977179
transform 1 0 51060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_550
timestamp 1649977179
transform 1 0 51704 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_558
timestamp 1649977179
transform 1 0 52440 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_564
timestamp 1649977179
transform 1 0 52992 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_571
timestamp 1649977179
transform 1 0 53636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_578
timestamp 1649977179
transform 1 0 54280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_585
timestamp 1649977179
transform 1 0 54924 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_592
timestamp 1649977179
transform 1 0 55568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_599
timestamp 1649977179
transform 1 0 56212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_606
timestamp 1649977179
transform 1 0 56856 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_614
timestamp 1649977179
transform 1 0 57592 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_620
timestamp 1649977179
transform 1 0 58144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_627
timestamp 1649977179
transform 1 0 58788 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_634
timestamp 1649977179
transform 1 0 59432 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_641
timestamp 1649977179
transform 1 0 60076 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_648
timestamp 1649977179
transform 1 0 60720 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_655
timestamp 1649977179
transform 1 0 61364 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_662
timestamp 1649977179
transform 1 0 62008 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_670
timestamp 1649977179
transform 1 0 62744 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_676
timestamp 1649977179
transform 1 0 63296 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_688
timestamp 1649977179
transform 1 0 64400 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_700
timestamp 1649977179
transform 1 0 65504 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_712
timestamp 1649977179
transform 1 0 66608 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_724
timestamp 1649977179
transform 1 0 67712 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_729
timestamp 1649977179
transform 1 0 68172 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7
timestamp 1649977179
transform 1 0 1748 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_17
timestamp 1649977179
transform 1 0 2668 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1649977179
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_34
timestamp 1649977179
transform 1 0 4232 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_40
timestamp 1649977179
transform 1 0 4784 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_50
timestamp 1649977179
transform 1 0 5704 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_61
timestamp 1649977179
transform 1 0 6716 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_68
timestamp 1649977179
transform 1 0 7360 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_90
timestamp 1649977179
transform 1 0 9384 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_99
timestamp 1649977179
transform 1 0 10212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_108
timestamp 1649977179
transform 1 0 11040 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_123
timestamp 1649977179
transform 1 0 12420 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_131
timestamp 1649977179
transform 1 0 13156 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1649977179
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_146
timestamp 1649977179
transform 1 0 14536 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_154
timestamp 1649977179
transform 1 0 15272 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_162
timestamp 1649977179
transform 1 0 16008 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_170
timestamp 1649977179
transform 1 0 16744 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_177
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_181
timestamp 1649977179
transform 1 0 17756 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_185
timestamp 1649977179
transform 1 0 18124 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1649977179
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_207
timestamp 1649977179
transform 1 0 20148 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_213
timestamp 1649977179
transform 1 0 20700 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_220
timestamp 1649977179
transform 1 0 21344 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_224
timestamp 1649977179
transform 1 0 21712 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_228
timestamp 1649977179
transform 1 0 22080 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_235
timestamp 1649977179
transform 1 0 22724 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_244
timestamp 1649977179
transform 1 0 23552 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1649977179
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_258
timestamp 1649977179
transform 1 0 24840 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_265
timestamp 1649977179
transform 1 0 25484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_272
timestamp 1649977179
transform 1 0 26128 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_284
timestamp 1649977179
transform 1 0 27232 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_295
timestamp 1649977179
transform 1 0 28244 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_304
timestamp 1649977179
transform 1 0 29072 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_309
timestamp 1649977179
transform 1 0 29532 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_313
timestamp 1649977179
transform 1 0 29900 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_322
timestamp 1649977179
transform 1 0 30728 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_329
timestamp 1649977179
transform 1 0 31372 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_349
timestamp 1649977179
transform 1 0 33212 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_361
timestamp 1649977179
transform 1 0 34316 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1649977179
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1649977179
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1649977179
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1649977179
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1649977179
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1649977179
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_424
timestamp 1649977179
transform 1 0 40112 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_431
timestamp 1649977179
transform 1 0 40756 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_438
timestamp 1649977179
transform 1 0 41400 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_445
timestamp 1649977179
transform 1 0 42044 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_454
timestamp 1649977179
transform 1 0 42872 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_461
timestamp 1649977179
transform 1 0 43516 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_473
timestamp 1649977179
transform 1 0 44620 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_477
timestamp 1649977179
transform 1 0 44988 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_481
timestamp 1649977179
transform 1 0 45356 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_488
timestamp 1649977179
transform 1 0 46000 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_495
timestamp 1649977179
transform 1 0 46644 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_502
timestamp 1649977179
transform 1 0 47288 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_511
timestamp 1649977179
transform 1 0 48116 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_519
timestamp 1649977179
transform 1 0 48852 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_523
timestamp 1649977179
transform 1 0 49220 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1649977179
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_533
timestamp 1649977179
transform 1 0 50140 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_538
timestamp 1649977179
transform 1 0 50600 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_545
timestamp 1649977179
transform 1 0 51244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_552
timestamp 1649977179
transform 1 0 51888 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_560
timestamp 1649977179
transform 1 0 52624 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_565
timestamp 1649977179
transform 1 0 53084 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_572
timestamp 1649977179
transform 1 0 53728 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_584
timestamp 1649977179
transform 1 0 54832 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_592
timestamp 1649977179
transform 1 0 55568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_599
timestamp 1649977179
transform 1 0 56212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_606
timestamp 1649977179
transform 1 0 56856 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_613
timestamp 1649977179
transform 1 0 57500 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_620
timestamp 1649977179
transform 1 0 58144 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_627
timestamp 1649977179
transform 1 0 58788 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_634
timestamp 1649977179
transform 1 0 59432 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_642
timestamp 1649977179
transform 1 0 60168 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_648
timestamp 1649977179
transform 1 0 60720 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_655
timestamp 1649977179
transform 1 0 61364 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_662
timestamp 1649977179
transform 1 0 62008 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_674
timestamp 1649977179
transform 1 0 63112 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_686
timestamp 1649977179
transform 1 0 64216 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_698
timestamp 1649977179
transform 1 0 65320 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_701
timestamp 1649977179
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_713
timestamp 1649977179
transform 1 0 66700 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_725
timestamp 1649977179
transform 1 0 67804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_729
timestamp 1649977179
transform 1 0 68172 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_12
timestamp 1649977179
transform 1 0 2208 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_18
timestamp 1649977179
transform 1 0 2760 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_35
timestamp 1649977179
transform 1 0 4324 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_41
timestamp 1649977179
transform 1 0 4876 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_45
timestamp 1649977179
transform 1 0 5244 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1649977179
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_62
timestamp 1649977179
transform 1 0 6808 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_75
timestamp 1649977179
transform 1 0 8004 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_83
timestamp 1649977179
transform 1 0 8740 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_88
timestamp 1649977179
transform 1 0 9200 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_97
timestamp 1649977179
transform 1 0 10028 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1649977179
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_127
timestamp 1649977179
transform 1 0 12788 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_133
timestamp 1649977179
transform 1 0 13340 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_145
timestamp 1649977179
transform 1 0 14444 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_151
timestamp 1649977179
transform 1 0 14996 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_160
timestamp 1649977179
transform 1 0 15824 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_185
timestamp 1649977179
transform 1 0 18124 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_194
timestamp 1649977179
transform 1 0 18952 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_201
timestamp 1649977179
transform 1 0 19596 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_207
timestamp 1649977179
transform 1 0 20148 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_214
timestamp 1649977179
transform 1 0 20792 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_220
timestamp 1649977179
transform 1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_228
timestamp 1649977179
transform 1 0 22080 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_235
timestamp 1649977179
transform 1 0 22724 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_239
timestamp 1649977179
transform 1 0 23092 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_248
timestamp 1649977179
transform 1 0 23920 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_268
timestamp 1649977179
transform 1 0 25760 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_276
timestamp 1649977179
transform 1 0 26496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_281
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1649977179
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_305
timestamp 1649977179
transform 1 0 29164 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_325
timestamp 1649977179
transform 1 0 31004 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_333
timestamp 1649977179
transform 1 0 31740 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_337
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_346
timestamp 1649977179
transform 1 0 32936 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_368
timestamp 1649977179
transform 1 0 34960 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_388
timestamp 1649977179
transform 1 0 36800 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1649977179
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1649977179
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1649977179
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1649977179
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1649977179
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1649977179
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1649977179
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1649977179
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1649977179
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1649977179
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1649977179
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1649977179
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1649977179
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1649977179
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1649977179
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1649977179
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1649977179
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1649977179
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1649977179
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1649977179
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1649977179
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_597
timestamp 1649977179
transform 1 0 56028 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_602
timestamp 1649977179
transform 1 0 56488 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1649977179
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1649977179
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_620
timestamp 1649977179
transform 1 0 58144 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_627
timestamp 1649977179
transform 1 0 58788 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_634
timestamp 1649977179
transform 1 0 59432 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_641
timestamp 1649977179
transform 1 0 60076 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_648
timestamp 1649977179
transform 1 0 60720 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_655
timestamp 1649977179
transform 1 0 61364 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_667
timestamp 1649977179
transform 1 0 62468 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 1649977179
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_673
timestamp 1649977179
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_685
timestamp 1649977179
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_697
timestamp 1649977179
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_709
timestamp 1649977179
transform 1 0 66332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_721
timestamp 1649977179
transform 1 0 67436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 1649977179
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_729
timestamp 1649977179
transform 1 0 68172 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_6
timestamp 1649977179
transform 1 0 1656 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_19
timestamp 1649977179
transform 1 0 2852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_32
timestamp 1649977179
transform 1 0 4048 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_52
timestamp 1649977179
transform 1 0 5888 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_62
timestamp 1649977179
transform 1 0 6808 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_70
timestamp 1649977179
transform 1 0 7544 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_76
timestamp 1649977179
transform 1 0 8096 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1649977179
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_93
timestamp 1649977179
transform 1 0 9660 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_105
timestamp 1649977179
transform 1 0 10764 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_122
timestamp 1649977179
transform 1 0 12328 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1649977179
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_152
timestamp 1649977179
transform 1 0 15088 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_172
timestamp 1649977179
transform 1 0 16928 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_179
timestamp 1649977179
transform 1 0 17572 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1649977179
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_213
timestamp 1649977179
transform 1 0 20700 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_233
timestamp 1649977179
transform 1 0 22540 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_244
timestamp 1649977179
transform 1 0 23552 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_255
timestamp 1649977179
transform 1 0 24564 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_261
timestamp 1649977179
transform 1 0 25116 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_264
timestamp 1649977179
transform 1 0 25392 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_284
timestamp 1649977179
transform 1 0 27232 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_304
timestamp 1649977179
transform 1 0 29072 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1649977179
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1649977179
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_333
timestamp 1649977179
transform 1 0 31740 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_341
timestamp 1649977179
transform 1 0 32476 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_349
timestamp 1649977179
transform 1 0 33212 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1649977179
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1649977179
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_370
timestamp 1649977179
transform 1 0 35144 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_376
timestamp 1649977179
transform 1 0 35696 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_382
timestamp 1649977179
transform 1 0 36248 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_410
timestamp 1649977179
transform 1 0 38824 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_418
timestamp 1649977179
transform 1 0 39560 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1649977179
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1649977179
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1649977179
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1649977179
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1649977179
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1649977179
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1649977179
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1649977179
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1649977179
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1649977179
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1649977179
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1649977179
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1649977179
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1649977179
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1649977179
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1649977179
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1649977179
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1649977179
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1649977179
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_601
timestamp 1649977179
transform 1 0 56396 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_609
timestamp 1649977179
transform 1 0 57132 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_613
timestamp 1649977179
transform 1 0 57500 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_620
timestamp 1649977179
transform 1 0 58144 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_627
timestamp 1649977179
transform 1 0 58788 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_634
timestamp 1649977179
transform 1 0 59432 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_642
timestamp 1649977179
transform 1 0 60168 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_648
timestamp 1649977179
transform 1 0 60720 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_660
timestamp 1649977179
transform 1 0 61824 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_672
timestamp 1649977179
transform 1 0 62928 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_684
timestamp 1649977179
transform 1 0 64032 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_696
timestamp 1649977179
transform 1 0 65136 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_701
timestamp 1649977179
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_713
timestamp 1649977179
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_725
timestamp 1649977179
transform 1 0 67804 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_8
timestamp 1649977179
transform 1 0 1840 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_21
timestamp 1649977179
transform 1 0 3036 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_24
timestamp 1649977179
transform 1 0 3312 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_30
timestamp 1649977179
transform 1 0 3864 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_36
timestamp 1649977179
transform 1 0 4416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_43
timestamp 1649977179
transform 1 0 5060 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1649977179
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_67
timestamp 1649977179
transform 1 0 7268 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_77
timestamp 1649977179
transform 1 0 8188 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_85
timestamp 1649977179
transform 1 0 8924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_98
timestamp 1649977179
transform 1 0 10120 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1649977179
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_121
timestamp 1649977179
transform 1 0 12236 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_132
timestamp 1649977179
transform 1 0 13248 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_146
timestamp 1649977179
transform 1 0 14536 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_154
timestamp 1649977179
transform 1 0 15272 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_160
timestamp 1649977179
transform 1 0 15824 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_164
timestamp 1649977179
transform 1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_173
timestamp 1649977179
transform 1 0 17020 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_180
timestamp 1649977179
transform 1 0 17664 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_186
timestamp 1649977179
transform 1 0 18216 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_190
timestamp 1649977179
transform 1 0 18584 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_199
timestamp 1649977179
transform 1 0 19412 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_206
timestamp 1649977179
transform 1 0 20056 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_220
timestamp 1649977179
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_228
timestamp 1649977179
transform 1 0 22080 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_234
timestamp 1649977179
transform 1 0 22632 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_237
timestamp 1649977179
transform 1 0 22908 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_249
timestamp 1649977179
transform 1 0 24012 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_263
timestamp 1649977179
transform 1 0 25300 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_276
timestamp 1649977179
transform 1 0 26496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_281
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_290
timestamp 1649977179
transform 1 0 27784 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_302
timestamp 1649977179
transform 1 0 28888 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_310
timestamp 1649977179
transform 1 0 29624 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_328
timestamp 1649977179
transform 1 0 31280 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_337
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_341
timestamp 1649977179
transform 1 0 32476 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_353
timestamp 1649977179
transform 1 0 33580 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_365
timestamp 1649977179
transform 1 0 34684 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_371
timestamp 1649977179
transform 1 0 35236 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1649977179
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1649977179
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_398
timestamp 1649977179
transform 1 0 37720 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_410
timestamp 1649977179
transform 1 0 38824 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_427
timestamp 1649977179
transform 1 0 40388 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_439
timestamp 1649977179
transform 1 0 41492 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1649977179
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1649977179
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1649977179
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1649977179
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1649977179
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1649977179
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1649977179
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1649977179
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1649977179
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1649977179
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1649977179
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1649977179
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1649977179
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1649977179
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1649977179
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1649977179
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1649977179
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1649977179
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1649977179
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_617
timestamp 1649977179
transform 1 0 57868 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_625
timestamp 1649977179
transform 1 0 58604 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_630
timestamp 1649977179
transform 1 0 59064 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_637
timestamp 1649977179
transform 1 0 59708 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_644
timestamp 1649977179
transform 1 0 60352 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_656
timestamp 1649977179
transform 1 0 61456 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_668
timestamp 1649977179
transform 1 0 62560 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_673
timestamp 1649977179
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_685
timestamp 1649977179
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_697
timestamp 1649977179
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_709
timestamp 1649977179
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_724
timestamp 1649977179
transform 1 0 67712 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_729
timestamp 1649977179
transform 1 0 68172 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_5
timestamp 1649977179
transform 1 0 1564 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_12
timestamp 1649977179
transform 1 0 2208 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_18
timestamp 1649977179
transform 1 0 2760 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1649977179
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_32
timestamp 1649977179
transform 1 0 4048 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_42
timestamp 1649977179
transform 1 0 4968 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_48
timestamp 1649977179
transform 1 0 5520 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_55
timestamp 1649977179
transform 1 0 6164 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_63
timestamp 1649977179
transform 1 0 6900 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_89
timestamp 1649977179
transform 1 0 9292 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_95
timestamp 1649977179
transform 1 0 9844 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_116
timestamp 1649977179
transform 1 0 11776 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp 1649977179
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_145
timestamp 1649977179
transform 1 0 14444 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_154
timestamp 1649977179
transform 1 0 15272 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_164
timestamp 1649977179
transform 1 0 16192 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_168
timestamp 1649977179
transform 1 0 16560 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_178
timestamp 1649977179
transform 1 0 17480 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_188
timestamp 1649977179
transform 1 0 18400 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_206
timestamp 1649977179
transform 1 0 20056 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_224
timestamp 1649977179
transform 1 0 21712 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_244
timestamp 1649977179
transform 1 0 23552 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_253
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_261
timestamp 1649977179
transform 1 0 25116 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_269
timestamp 1649977179
transform 1 0 25852 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_273
timestamp 1649977179
transform 1 0 26220 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_278
timestamp 1649977179
transform 1 0 26680 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_284
timestamp 1649977179
transform 1 0 27232 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_290
timestamp 1649977179
transform 1 0 27784 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_298
timestamp 1649977179
transform 1 0 28520 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_304
timestamp 1649977179
transform 1 0 29072 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_309
timestamp 1649977179
transform 1 0 29532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_320
timestamp 1649977179
transform 1 0 30544 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_326
timestamp 1649977179
transform 1 0 31096 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_336
timestamp 1649977179
transform 1 0 32016 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_360
timestamp 1649977179
transform 1 0 34224 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_375
timestamp 1649977179
transform 1 0 35604 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_381
timestamp 1649977179
transform 1 0 36156 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_387
timestamp 1649977179
transform 1 0 36708 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_399
timestamp 1649977179
transform 1 0 37812 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_405
timestamp 1649977179
transform 1 0 38364 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_417
timestamp 1649977179
transform 1 0 39468 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1649977179
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1649977179
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1649977179
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1649977179
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1649977179
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1649977179
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1649977179
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1649977179
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1649977179
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1649977179
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1649977179
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1649977179
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1649977179
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1649977179
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1649977179
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1649977179
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1649977179
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1649977179
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1649977179
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1649977179
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1649977179
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_625
timestamp 1649977179
transform 1 0 58604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_637
timestamp 1649977179
transform 1 0 59708 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 1649977179
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_645
timestamp 1649977179
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_657
timestamp 1649977179
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_669
timestamp 1649977179
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_681
timestamp 1649977179
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_693
timestamp 1649977179
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 1649977179
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_701
timestamp 1649977179
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_713
timestamp 1649977179
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_725
timestamp 1649977179
transform 1 0 67804 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_11
timestamp 1649977179
transform 1 0 2116 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_17
timestamp 1649977179
transform 1 0 2668 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_34
timestamp 1649977179
transform 1 0 4232 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_49
timestamp 1649977179
transform 1 0 5612 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_68
timestamp 1649977179
transform 1 0 7360 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_80
timestamp 1649977179
transform 1 0 8464 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_96
timestamp 1649977179
transform 1 0 9936 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_108
timestamp 1649977179
transform 1 0 11040 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_129
timestamp 1649977179
transform 1 0 12972 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_162
timestamp 1649977179
transform 1 0 16008 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_202
timestamp 1649977179
transform 1 0 19688 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_209
timestamp 1649977179
transform 1 0 20332 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_216
timestamp 1649977179
transform 1 0 20976 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_225
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_229
timestamp 1649977179
transform 1 0 22172 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_246
timestamp 1649977179
transform 1 0 23736 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_270
timestamp 1649977179
transform 1 0 25944 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_276
timestamp 1649977179
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_281
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_298
timestamp 1649977179
transform 1 0 28520 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_312
timestamp 1649977179
transform 1 0 29808 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_332
timestamp 1649977179
transform 1 0 31648 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_337
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_345
timestamp 1649977179
transform 1 0 32844 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_349
timestamp 1649977179
transform 1 0 33212 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_361
timestamp 1649977179
transform 1 0 34316 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_369
timestamp 1649977179
transform 1 0 35052 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_378
timestamp 1649977179
transform 1 0 35880 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_387
timestamp 1649977179
transform 1 0 36708 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1649977179
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_398
timestamp 1649977179
transform 1 0 37720 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_410
timestamp 1649977179
transform 1 0 38824 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_422
timestamp 1649977179
transform 1 0 39928 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_434
timestamp 1649977179
transform 1 0 41032 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_446
timestamp 1649977179
transform 1 0 42136 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1649977179
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1649977179
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1649977179
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1649977179
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1649977179
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1649977179
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1649977179
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1649977179
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1649977179
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1649977179
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1649977179
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1649977179
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1649977179
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1649977179
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1649977179
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1649977179
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1649977179
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1649977179
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_617
timestamp 1649977179
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_629
timestamp 1649977179
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_641
timestamp 1649977179
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_653
timestamp 1649977179
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 1649977179
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1649977179
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_673
timestamp 1649977179
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_685
timestamp 1649977179
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_697
timestamp 1649977179
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_709
timestamp 1649977179
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_724
timestamp 1649977179
transform 1 0 67712 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_729
timestamp 1649977179
transform 1 0 68172 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_11
timestamp 1649977179
transform 1 0 2116 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_18
timestamp 1649977179
transform 1 0 2760 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1649977179
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_66
timestamp 1649977179
transform 1 0 7176 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_70
timestamp 1649977179
transform 1 0 7544 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_96
timestamp 1649977179
transform 1 0 9936 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_109
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_121
timestamp 1649977179
transform 1 0 12236 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_125
timestamp 1649977179
transform 1 0 12604 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_129
timestamp 1649977179
transform 1 0 12972 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_136
timestamp 1649977179
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_147
timestamp 1649977179
transform 1 0 14628 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_154
timestamp 1649977179
transform 1 0 15272 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_161
timestamp 1649977179
transform 1 0 15916 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_181
timestamp 1649977179
transform 1 0 17756 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 1649977179
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_207
timestamp 1649977179
transform 1 0 20148 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_227
timestamp 1649977179
transform 1 0 21988 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_241
timestamp 1649977179
transform 1 0 23276 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_245
timestamp 1649977179
transform 1 0 23644 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_248
timestamp 1649977179
transform 1 0 23920 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_253
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_257
timestamp 1649977179
transform 1 0 24748 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_262
timestamp 1649977179
transform 1 0 25208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_271
timestamp 1649977179
transform 1 0 26036 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_283
timestamp 1649977179
transform 1 0 27140 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_295
timestamp 1649977179
transform 1 0 28244 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_301
timestamp 1649977179
transform 1 0 28796 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_304
timestamp 1649977179
transform 1 0 29072 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_314
timestamp 1649977179
transform 1 0 29992 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_326
timestamp 1649977179
transform 1 0 31096 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_334
timestamp 1649977179
transform 1 0 31832 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_352
timestamp 1649977179
transform 1 0 33488 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_368
timestamp 1649977179
transform 1 0 34960 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_388
timestamp 1649977179
transform 1 0 36800 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_399
timestamp 1649977179
transform 1 0 37812 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_408
timestamp 1649977179
transform 1 0 38640 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_437
timestamp 1649977179
transform 1 0 41308 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_449
timestamp 1649977179
transform 1 0 42412 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_461
timestamp 1649977179
transform 1 0 43516 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_473
timestamp 1649977179
transform 1 0 44620 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1649977179
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1649977179
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1649977179
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1649977179
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1649977179
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1649977179
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1649977179
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1649977179
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1649977179
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1649977179
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1649977179
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1649977179
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1649977179
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1649977179
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1649977179
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_625
timestamp 1649977179
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 1649977179
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 1649977179
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_645
timestamp 1649977179
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_657
timestamp 1649977179
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_669
timestamp 1649977179
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_681
timestamp 1649977179
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_693
timestamp 1649977179
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 1649977179
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_701
timestamp 1649977179
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_713
timestamp 1649977179
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_725
timestamp 1649977179
transform 1 0 67804 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_7
timestamp 1649977179
transform 1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_14
timestamp 1649977179
transform 1 0 2392 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_36
timestamp 1649977179
transform 1 0 4416 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_44
timestamp 1649977179
transform 1 0 5152 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_50
timestamp 1649977179
transform 1 0 5704 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_59
timestamp 1649977179
transform 1 0 6532 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_67
timestamp 1649977179
transform 1 0 7268 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_75
timestamp 1649977179
transform 1 0 8004 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_82
timestamp 1649977179
transform 1 0 8648 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_96
timestamp 1649977179
transform 1 0 9936 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_108
timestamp 1649977179
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_123
timestamp 1649977179
transform 1 0 12420 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_132
timestamp 1649977179
transform 1 0 13248 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_139
timestamp 1649977179
transform 1 0 13892 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_151
timestamp 1649977179
transform 1 0 14996 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_157
timestamp 1649977179
transform 1 0 15548 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1649977179
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_174
timestamp 1649977179
transform 1 0 17112 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_178
timestamp 1649977179
transform 1 0 17480 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_182
timestamp 1649977179
transform 1 0 17848 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_186
timestamp 1649977179
transform 1 0 18216 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_193
timestamp 1649977179
transform 1 0 18860 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_199
timestamp 1649977179
transform 1 0 19412 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1649977179
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1649977179
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1649977179
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_241
timestamp 1649977179
transform 1 0 23276 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_245
timestamp 1649977179
transform 1 0 23644 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_248
timestamp 1649977179
transform 1 0 23920 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_257
timestamp 1649977179
transform 1 0 24748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_269
timestamp 1649977179
transform 1 0 25852 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_275
timestamp 1649977179
transform 1 0 26404 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1649977179
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_281
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_292
timestamp 1649977179
transform 1 0 27968 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_303
timestamp 1649977179
transform 1 0 28980 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_327
timestamp 1649977179
transform 1 0 31188 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1649977179
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1649977179
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_349
timestamp 1649977179
transform 1 0 33212 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_358
timestamp 1649977179
transform 1 0 34040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_367
timestamp 1649977179
transform 1 0 34868 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_375
timestamp 1649977179
transform 1 0 35604 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_384
timestamp 1649977179
transform 1 0 36432 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_393
timestamp 1649977179
transform 1 0 37260 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_396
timestamp 1649977179
transform 1 0 37536 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_408
timestamp 1649977179
transform 1 0 38640 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_414
timestamp 1649977179
transform 1 0 39192 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_426
timestamp 1649977179
transform 1 0 40296 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_438
timestamp 1649977179
transform 1 0 41400 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_446
timestamp 1649977179
transform 1 0 42136 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1649977179
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1649977179
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1649977179
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1649977179
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1649977179
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1649977179
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1649977179
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1649977179
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1649977179
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1649977179
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1649977179
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1649977179
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1649977179
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1649977179
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1649977179
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_597
timestamp 1649977179
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1649977179
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1649977179
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_617
timestamp 1649977179
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_629
timestamp 1649977179
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_641
timestamp 1649977179
transform 1 0 60076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_653
timestamp 1649977179
transform 1 0 61180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_665
timestamp 1649977179
transform 1 0 62284 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_671
timestamp 1649977179
transform 1 0 62836 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_673
timestamp 1649977179
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_685
timestamp 1649977179
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_697
timestamp 1649977179
transform 1 0 65228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_709
timestamp 1649977179
transform 1 0 66332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_721
timestamp 1649977179
transform 1 0 67436 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_727
timestamp 1649977179
transform 1 0 67988 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_729
timestamp 1649977179
transform 1 0 68172 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_21
timestamp 1649977179
transform 1 0 3036 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_33
timestamp 1649977179
transform 1 0 4140 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_36
timestamp 1649977179
transform 1 0 4416 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_56
timestamp 1649977179
transform 1 0 6256 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_60
timestamp 1649977179
transform 1 0 6624 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_63
timestamp 1649977179
transform 1 0 6900 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_73
timestamp 1649977179
transform 1 0 7820 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_77
timestamp 1649977179
transform 1 0 8188 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1649977179
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_95
timestamp 1649977179
transform 1 0 9844 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_103
timestamp 1649977179
transform 1 0 10580 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_109
timestamp 1649977179
transform 1 0 11132 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_116
timestamp 1649977179
transform 1 0 11776 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 1649977179
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_145
timestamp 1649977179
transform 1 0 14444 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_162
timestamp 1649977179
transform 1 0 16008 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_170
timestamp 1649977179
transform 1 0 16744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_180
timestamp 1649977179
transform 1 0 17664 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_187
timestamp 1649977179
transform 1 0 18308 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1649977179
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_199
timestamp 1649977179
transform 1 0 19412 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_227
timestamp 1649977179
transform 1 0 21988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_239
timestamp 1649977179
transform 1 0 23092 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_247
timestamp 1649977179
transform 1 0 23828 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1649977179
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_256
timestamp 1649977179
transform 1 0 24656 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_270
timestamp 1649977179
transform 1 0 25944 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_281
timestamp 1649977179
transform 1 0 26956 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_295
timestamp 1649977179
transform 1 0 28244 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_301
timestamp 1649977179
transform 1 0 28796 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_304
timestamp 1649977179
transform 1 0 29072 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_317
timestamp 1649977179
transform 1 0 30268 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_325
timestamp 1649977179
transform 1 0 31004 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_343
timestamp 1649977179
transform 1 0 32660 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_351
timestamp 1649977179
transform 1 0 33396 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_360
timestamp 1649977179
transform 1 0 34224 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_367
timestamp 1649977179
transform 1 0 34868 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_373
timestamp 1649977179
transform 1 0 35420 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_387
timestamp 1649977179
transform 1 0 36708 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_393
timestamp 1649977179
transform 1 0 37260 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_399
timestamp 1649977179
transform 1 0 37812 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_408
timestamp 1649977179
transform 1 0 38640 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_414
timestamp 1649977179
transform 1 0 39192 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_437
timestamp 1649977179
transform 1 0 41308 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_449
timestamp 1649977179
transform 1 0 42412 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_461
timestamp 1649977179
transform 1 0 43516 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_473
timestamp 1649977179
transform 1 0 44620 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1649977179
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1649977179
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1649977179
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1649977179
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1649977179
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1649977179
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1649977179
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1649977179
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1649977179
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1649977179
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1649977179
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1649977179
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_589
timestamp 1649977179
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_601
timestamp 1649977179
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_613
timestamp 1649977179
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_625
timestamp 1649977179
transform 1 0 58604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_637
timestamp 1649977179
transform 1 0 59708 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_643
timestamp 1649977179
transform 1 0 60260 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_645
timestamp 1649977179
transform 1 0 60444 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_657
timestamp 1649977179
transform 1 0 61548 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_669
timestamp 1649977179
transform 1 0 62652 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_681
timestamp 1649977179
transform 1 0 63756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_693
timestamp 1649977179
transform 1 0 64860 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_699
timestamp 1649977179
transform 1 0 65412 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_701
timestamp 1649977179
transform 1 0 65596 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_713
timestamp 1649977179
transform 1 0 66700 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_725
timestamp 1649977179
transform 1 0 67804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_729
timestamp 1649977179
transform 1 0 68172 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_6
timestamp 1649977179
transform 1 0 1656 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_12
timestamp 1649977179
transform 1 0 2208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_32
timestamp 1649977179
transform 1 0 4048 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_11_43
timestamp 1649977179
transform 1 0 5060 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1649977179
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_59
timestamp 1649977179
transform 1 0 6532 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_63
timestamp 1649977179
transform 1 0 6900 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_70
timestamp 1649977179
transform 1 0 7544 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_80
timestamp 1649977179
transform 1 0 8464 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_86
timestamp 1649977179
transform 1 0 9016 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_94
timestamp 1649977179
transform 1 0 9752 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_101
timestamp 1649977179
transform 1 0 10396 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp 1649977179
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_115
timestamp 1649977179
transform 1 0 11684 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_128
timestamp 1649977179
transform 1 0 12880 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_146
timestamp 1649977179
transform 1 0 14536 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_154
timestamp 1649977179
transform 1 0 15272 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_158
timestamp 1649977179
transform 1 0 15640 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1649977179
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_173
timestamp 1649977179
transform 1 0 17020 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_177
timestamp 1649977179
transform 1 0 17388 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_194
timestamp 1649977179
transform 1 0 18952 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_200
timestamp 1649977179
transform 1 0 19504 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_212
timestamp 1649977179
transform 1 0 20608 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_244
timestamp 1649977179
transform 1 0 23552 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_262
timestamp 1649977179
transform 1 0 25208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_276
timestamp 1649977179
transform 1 0 26496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_291
timestamp 1649977179
transform 1 0 27876 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_302
timestamp 1649977179
transform 1 0 28888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_311
timestamp 1649977179
transform 1 0 29716 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_321
timestamp 1649977179
transform 1 0 30636 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_329
timestamp 1649977179
transform 1 0 31372 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_332
timestamp 1649977179
transform 1 0 31648 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_344
timestamp 1649977179
transform 1 0 32752 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_352
timestamp 1649977179
transform 1 0 33488 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_363
timestamp 1649977179
transform 1 0 34500 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_370
timestamp 1649977179
transform 1 0 35144 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_386
timestamp 1649977179
transform 1 0 36616 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_403
timestamp 1649977179
transform 1 0 38180 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1649977179
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1649977179
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1649977179
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1649977179
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1649977179
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1649977179
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1649977179
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1649977179
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1649977179
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1649977179
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1649977179
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1649977179
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1649977179
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1649977179
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1649977179
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1649977179
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1649977179
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_585
timestamp 1649977179
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_597
timestamp 1649977179
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1649977179
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1649977179
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_617
timestamp 1649977179
transform 1 0 57868 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_629
timestamp 1649977179
transform 1 0 58972 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_641
timestamp 1649977179
transform 1 0 60076 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_653
timestamp 1649977179
transform 1 0 61180 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_665
timestamp 1649977179
transform 1 0 62284 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_671
timestamp 1649977179
transform 1 0 62836 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_673
timestamp 1649977179
transform 1 0 63020 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_685
timestamp 1649977179
transform 1 0 64124 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_697
timestamp 1649977179
transform 1 0 65228 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_709
timestamp 1649977179
transform 1 0 66332 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_721
timestamp 1649977179
transform 1 0 67436 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_727
timestamp 1649977179
transform 1 0 67988 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_729
timestamp 1649977179
transform 1 0 68172 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_7
timestamp 1649977179
transform 1 0 1748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_16
timestamp 1649977179
transform 1 0 2576 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_22
timestamp 1649977179
transform 1 0 3128 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_34
timestamp 1649977179
transform 1 0 4232 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_40
timestamp 1649977179
transform 1 0 4784 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_48
timestamp 1649977179
transform 1 0 5520 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_71
timestamp 1649977179
transform 1 0 7636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_114
timestamp 1649977179
transform 1 0 11592 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_127
timestamp 1649977179
transform 1 0 12788 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp 1649977179
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_147
timestamp 1649977179
transform 1 0 14628 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_153
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_173
timestamp 1649977179
transform 1 0 17020 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_177
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_183
timestamp 1649977179
transform 1 0 17940 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 1649977179
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_201
timestamp 1649977179
transform 1 0 19596 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_210
timestamp 1649977179
transform 1 0 20424 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_222
timestamp 1649977179
transform 1 0 21528 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_244
timestamp 1649977179
transform 1 0 23552 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_258
timestamp 1649977179
transform 1 0 24840 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_266
timestamp 1649977179
transform 1 0 25576 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_270
timestamp 1649977179
transform 1 0 25944 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_287
timestamp 1649977179
transform 1 0 27508 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_299
timestamp 1649977179
transform 1 0 28612 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_302
timestamp 1649977179
transform 1 0 28888 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_309
timestamp 1649977179
transform 1 0 29532 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_319
timestamp 1649977179
transform 1 0 30452 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_330
timestamp 1649977179
transform 1 0 31464 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_336
timestamp 1649977179
transform 1 0 32016 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_353
timestamp 1649977179
transform 1 0 33580 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_359
timestamp 1649977179
transform 1 0 34132 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1649977179
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_365
timestamp 1649977179
transform 1 0 34684 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_368
timestamp 1649977179
transform 1 0 34960 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_382
timestamp 1649977179
transform 1 0 36248 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_393
timestamp 1649977179
transform 1 0 37260 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_402
timestamp 1649977179
transform 1 0 38088 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_411
timestamp 1649977179
transform 1 0 38916 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1649977179
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1649977179
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1649977179
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1649977179
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1649977179
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1649977179
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1649977179
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1649977179
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1649977179
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1649977179
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1649977179
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1649977179
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1649977179
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1649977179
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1649977179
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1649977179
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_569
timestamp 1649977179
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1649977179
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1649977179
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_589
timestamp 1649977179
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_601
timestamp 1649977179
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_613
timestamp 1649977179
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_625
timestamp 1649977179
transform 1 0 58604 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_637
timestamp 1649977179
transform 1 0 59708 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_643
timestamp 1649977179
transform 1 0 60260 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_645
timestamp 1649977179
transform 1 0 60444 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_657
timestamp 1649977179
transform 1 0 61548 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_669
timestamp 1649977179
transform 1 0 62652 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_681
timestamp 1649977179
transform 1 0 63756 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_693
timestamp 1649977179
transform 1 0 64860 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_699
timestamp 1649977179
transform 1 0 65412 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_701
timestamp 1649977179
transform 1 0 65596 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_713
timestamp 1649977179
transform 1 0 66700 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_725
timestamp 1649977179
transform 1 0 67804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_729
timestamp 1649977179
transform 1 0 68172 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_6
timestamp 1649977179
transform 1 0 1656 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_18
timestamp 1649977179
transform 1 0 2760 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_24
timestamp 1649977179
transform 1 0 3312 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_28
timestamp 1649977179
transform 1 0 3680 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_45
timestamp 1649977179
transform 1 0 5244 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_53
timestamp 1649977179
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_65
timestamp 1649977179
transform 1 0 7084 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_71
timestamp 1649977179
transform 1 0 7636 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_91
timestamp 1649977179
transform 1 0 9476 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_95
timestamp 1649977179
transform 1 0 9844 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_103
timestamp 1649977179
transform 1 0 10580 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_115
timestamp 1649977179
transform 1 0 11684 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_119
timestamp 1649977179
transform 1 0 12052 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_129
timestamp 1649977179
transform 1 0 12972 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_149
timestamp 1649977179
transform 1 0 14812 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_164
timestamp 1649977179
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_175
timestamp 1649977179
transform 1 0 17204 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_184
timestamp 1649977179
transform 1 0 18032 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_193
timestamp 1649977179
transform 1 0 18860 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_202
timestamp 1649977179
transform 1 0 19688 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_216
timestamp 1649977179
transform 1 0 20976 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_228
timestamp 1649977179
transform 1 0 22080 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_234
timestamp 1649977179
transform 1 0 22632 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_240
timestamp 1649977179
transform 1 0 23184 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_246
timestamp 1649977179
transform 1 0 23736 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_258
timestamp 1649977179
transform 1 0 24840 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_266
timestamp 1649977179
transform 1 0 25576 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_272
timestamp 1649977179
transform 1 0 26128 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_283
timestamp 1649977179
transform 1 0 27140 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_291
timestamp 1649977179
transform 1 0 27876 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_298
timestamp 1649977179
transform 1 0 28520 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_308
timestamp 1649977179
transform 1 0 29440 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_328
timestamp 1649977179
transform 1 0 31280 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_337
timestamp 1649977179
transform 1 0 32108 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_341
timestamp 1649977179
transform 1 0 32476 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_344
timestamp 1649977179
transform 1 0 32752 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_356
timestamp 1649977179
transform 1 0 33856 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_362
timestamp 1649977179
transform 1 0 34408 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_369
timestamp 1649977179
transform 1 0 35052 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_383
timestamp 1649977179
transform 1 0 36340 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1649977179
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_395
timestamp 1649977179
transform 1 0 37444 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_407
timestamp 1649977179
transform 1 0 38548 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_411
timestamp 1649977179
transform 1 0 38916 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_428
timestamp 1649977179
transform 1 0 40480 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_440
timestamp 1649977179
transform 1 0 41584 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1649977179
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1649977179
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1649977179
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1649977179
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1649977179
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1649977179
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1649977179
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1649977179
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1649977179
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1649977179
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1649977179
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1649977179
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1649977179
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1649977179
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_585
timestamp 1649977179
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_597
timestamp 1649977179
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1649977179
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1649977179
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_617
timestamp 1649977179
transform 1 0 57868 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_629
timestamp 1649977179
transform 1 0 58972 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_641
timestamp 1649977179
transform 1 0 60076 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_653
timestamp 1649977179
transform 1 0 61180 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_665
timestamp 1649977179
transform 1 0 62284 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_671
timestamp 1649977179
transform 1 0 62836 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_673
timestamp 1649977179
transform 1 0 63020 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_685
timestamp 1649977179
transform 1 0 64124 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_697
timestamp 1649977179
transform 1 0 65228 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_709
timestamp 1649977179
transform 1 0 66332 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_721
timestamp 1649977179
transform 1 0 67436 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_727
timestamp 1649977179
transform 1 0 67988 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_729
timestamp 1649977179
transform 1 0 68172 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_7
timestamp 1649977179
transform 1 0 1748 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_13
timestamp 1649977179
transform 1 0 2300 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_19
timestamp 1649977179
transform 1 0 2852 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_34
timestamp 1649977179
transform 1 0 4232 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_40
timestamp 1649977179
transform 1 0 4784 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_52
timestamp 1649977179
transform 1 0 5888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_60
timestamp 1649977179
transform 1 0 6624 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_68
timestamp 1649977179
transform 1 0 7360 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1649977179
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_87
timestamp 1649977179
transform 1 0 9108 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_100
timestamp 1649977179
transform 1 0 10304 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_127
timestamp 1649977179
transform 1 0 12788 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_133
timestamp 1649977179
transform 1 0 13340 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_136
timestamp 1649977179
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_143
timestamp 1649977179
transform 1 0 14260 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_149
timestamp 1649977179
transform 1 0 14812 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_155
timestamp 1649977179
transform 1 0 15364 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_167
timestamp 1649977179
transform 1 0 16468 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_180
timestamp 1649977179
transform 1 0 17664 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_192
timestamp 1649977179
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_199
timestamp 1649977179
transform 1 0 19412 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_211
timestamp 1649977179
transform 1 0 20516 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_215
timestamp 1649977179
transform 1 0 20884 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_232
timestamp 1649977179
transform 1 0 22448 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_238
timestamp 1649977179
transform 1 0 23000 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_244
timestamp 1649977179
transform 1 0 23552 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_248
timestamp 1649977179
transform 1 0 23920 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_253
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_257
timestamp 1649977179
transform 1 0 24748 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_268
timestamp 1649977179
transform 1 0 25760 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_280
timestamp 1649977179
transform 1 0 26864 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_291
timestamp 1649977179
transform 1 0 27876 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_297
timestamp 1649977179
transform 1 0 28428 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_304
timestamp 1649977179
transform 1 0 29072 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_311
timestamp 1649977179
transform 1 0 29716 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_323
timestamp 1649977179
transform 1 0 30820 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_347
timestamp 1649977179
transform 1 0 33028 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_355
timestamp 1649977179
transform 1 0 33764 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_360
timestamp 1649977179
transform 1 0 34224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_368
timestamp 1649977179
transform 1 0 34960 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_382
timestamp 1649977179
transform 1 0 36248 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_388
timestamp 1649977179
transform 1 0 36800 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_396
timestamp 1649977179
transform 1 0 37536 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_405
timestamp 1649977179
transform 1 0 38364 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_417
timestamp 1649977179
transform 1 0 39468 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1649977179
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1649977179
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1649977179
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1649977179
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1649977179
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1649977179
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1649977179
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1649977179
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1649977179
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1649977179
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1649977179
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1649977179
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1649977179
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1649977179
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_557
timestamp 1649977179
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_569
timestamp 1649977179
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1649977179
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1649977179
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1649977179
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_601
timestamp 1649977179
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_613
timestamp 1649977179
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_625
timestamp 1649977179
transform 1 0 58604 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_637
timestamp 1649977179
transform 1 0 59708 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_643
timestamp 1649977179
transform 1 0 60260 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_645
timestamp 1649977179
transform 1 0 60444 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_657
timestamp 1649977179
transform 1 0 61548 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_669
timestamp 1649977179
transform 1 0 62652 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_681
timestamp 1649977179
transform 1 0 63756 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_693
timestamp 1649977179
transform 1 0 64860 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_699
timestamp 1649977179
transform 1 0 65412 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_701
timestamp 1649977179
transform 1 0 65596 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_713
timestamp 1649977179
transform 1 0 66700 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_725
timestamp 1649977179
transform 1 0 67804 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_21
timestamp 1649977179
transform 1 0 3036 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_38
timestamp 1649977179
transform 1 0 4600 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1649977179
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_65
timestamp 1649977179
transform 1 0 7084 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_71
timestamp 1649977179
transform 1 0 7636 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_77
timestamp 1649977179
transform 1 0 8188 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_83
timestamp 1649977179
transform 1 0 8740 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_95
timestamp 1649977179
transform 1 0 9844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1649977179
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_129
timestamp 1649977179
transform 1 0 12972 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_146
timestamp 1649977179
transform 1 0 14536 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_158
timestamp 1649977179
transform 1 0 15640 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1649977179
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_177
timestamp 1649977179
transform 1 0 17388 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_185
timestamp 1649977179
transform 1 0 18124 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_209
timestamp 1649977179
transform 1 0 20332 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_218
timestamp 1649977179
transform 1 0 21160 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_15_225
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_232
timestamp 1649977179
transform 1 0 22448 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_241
timestamp 1649977179
transform 1 0 23276 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_252
timestamp 1649977179
transform 1 0 24288 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_258
timestamp 1649977179
transform 1 0 24840 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_262
timestamp 1649977179
transform 1 0 25208 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_268
timestamp 1649977179
transform 1 0 25760 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_274
timestamp 1649977179
transform 1 0 26312 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_293
timestamp 1649977179
transform 1 0 28060 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_303
timestamp 1649977179
transform 1 0 28980 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_313
timestamp 1649977179
transform 1 0 29900 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_325
timestamp 1649977179
transform 1 0 31004 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_333
timestamp 1649977179
transform 1 0 31740 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_337
timestamp 1649977179
transform 1 0 32108 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_345
timestamp 1649977179
transform 1 0 32844 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_357
timestamp 1649977179
transform 1 0 33948 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_365
timestamp 1649977179
transform 1 0 34684 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_374
timestamp 1649977179
transform 1 0 35512 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_388
timestamp 1649977179
transform 1 0 36800 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_396
timestamp 1649977179
transform 1 0 37536 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_400
timestamp 1649977179
transform 1 0 37904 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_409
timestamp 1649977179
transform 1 0 38732 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1649977179
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1649977179
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1649977179
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1649977179
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1649977179
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1649977179
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1649977179
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1649977179
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1649977179
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1649977179
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1649977179
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1649977179
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1649977179
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1649977179
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1649977179
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1649977179
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_573
timestamp 1649977179
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_585
timestamp 1649977179
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_597
timestamp 1649977179
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1649977179
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1649977179
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_617
timestamp 1649977179
transform 1 0 57868 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_629
timestamp 1649977179
transform 1 0 58972 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_641
timestamp 1649977179
transform 1 0 60076 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_653
timestamp 1649977179
transform 1 0 61180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_665
timestamp 1649977179
transform 1 0 62284 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_671
timestamp 1649977179
transform 1 0 62836 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_673
timestamp 1649977179
transform 1 0 63020 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_685
timestamp 1649977179
transform 1 0 64124 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_697
timestamp 1649977179
transform 1 0 65228 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_709
timestamp 1649977179
transform 1 0 66332 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_724
timestamp 1649977179
transform 1 0 67712 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_729
timestamp 1649977179
transform 1 0 68172 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_14
timestamp 1649977179
transform 1 0 2392 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_20
timestamp 1649977179
transform 1 0 2944 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_60
timestamp 1649977179
transform 1 0 6624 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_64
timestamp 1649977179
transform 1 0 6992 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_67
timestamp 1649977179
transform 1 0 7268 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_79
timestamp 1649977179
transform 1 0 8372 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_101
timestamp 1649977179
transform 1 0 10396 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_113
timestamp 1649977179
transform 1 0 11500 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_119
timestamp 1649977179
transform 1 0 12052 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_127
timestamp 1649977179
transform 1 0 12788 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_135
timestamp 1649977179
transform 1 0 13524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_160
timestamp 1649977179
transform 1 0 15824 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_182
timestamp 1649977179
transform 1 0 17848 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_191
timestamp 1649977179
transform 1 0 18676 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1649977179
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_201
timestamp 1649977179
transform 1 0 19596 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_210
timestamp 1649977179
transform 1 0 20424 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_216
timestamp 1649977179
transform 1 0 20976 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_222
timestamp 1649977179
transform 1 0 21528 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_228
timestamp 1649977179
transform 1 0 22080 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_234
timestamp 1649977179
transform 1 0 22632 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_242
timestamp 1649977179
transform 1 0 23368 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_248
timestamp 1649977179
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_253
timestamp 1649977179
transform 1 0 24380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_264
timestamp 1649977179
transform 1 0 25392 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_270
timestamp 1649977179
transform 1 0 25944 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_292
timestamp 1649977179
transform 1 0 27968 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_303
timestamp 1649977179
transform 1 0 28980 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1649977179
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_316
timestamp 1649977179
transform 1 0 30176 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_328
timestamp 1649977179
transform 1 0 31280 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_339
timestamp 1649977179
transform 1 0 32292 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_345
timestamp 1649977179
transform 1 0 32844 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_354
timestamp 1649977179
transform 1 0 33672 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_360
timestamp 1649977179
transform 1 0 34224 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_370
timestamp 1649977179
transform 1 0 35144 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_377
timestamp 1649977179
transform 1 0 35788 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_383
timestamp 1649977179
transform 1 0 36340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_389
timestamp 1649977179
transform 1 0 36892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_397
timestamp 1649977179
transform 1 0 37628 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_403
timestamp 1649977179
transform 1 0 38180 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_409
timestamp 1649977179
transform 1 0 38732 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_417
timestamp 1649977179
transform 1 0 39468 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1649977179
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1649977179
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1649977179
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1649977179
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1649977179
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1649977179
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1649977179
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1649977179
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1649977179
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1649977179
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1649977179
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1649977179
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1649977179
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1649977179
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_557
timestamp 1649977179
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_569
timestamp 1649977179
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1649977179
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1649977179
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_589
timestamp 1649977179
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_601
timestamp 1649977179
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_613
timestamp 1649977179
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_625
timestamp 1649977179
transform 1 0 58604 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_637
timestamp 1649977179
transform 1 0 59708 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_643
timestamp 1649977179
transform 1 0 60260 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_645
timestamp 1649977179
transform 1 0 60444 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_657
timestamp 1649977179
transform 1 0 61548 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_669
timestamp 1649977179
transform 1 0 62652 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_681
timestamp 1649977179
transform 1 0 63756 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_693
timestamp 1649977179
transform 1 0 64860 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_699
timestamp 1649977179
transform 1 0 65412 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_701
timestamp 1649977179
transform 1 0 65596 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_713
timestamp 1649977179
transform 1 0 66700 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_725
timestamp 1649977179
transform 1 0 67804 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_17
timestamp 1649977179
transform 1 0 2668 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_21
timestamp 1649977179
transform 1 0 3036 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_38
timestamp 1649977179
transform 1 0 4600 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_46
timestamp 1649977179
transform 1 0 5336 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1649977179
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_81
timestamp 1649977179
transform 1 0 8556 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_87
timestamp 1649977179
transform 1 0 9108 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_93
timestamp 1649977179
transform 1 0 9660 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_97
timestamp 1649977179
transform 1 0 10028 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_108
timestamp 1649977179
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_120
timestamp 1649977179
transform 1 0 12144 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_127
timestamp 1649977179
transform 1 0 12788 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_137
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_145
timestamp 1649977179
transform 1 0 14444 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_151
timestamp 1649977179
transform 1 0 14996 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_159
timestamp 1649977179
transform 1 0 15732 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1649977179
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_171
timestamp 1649977179
transform 1 0 16836 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_181
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_190
timestamp 1649977179
transform 1 0 18584 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_196
timestamp 1649977179
transform 1 0 19136 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_199
timestamp 1649977179
transform 1 0 19412 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_203
timestamp 1649977179
transform 1 0 19780 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1649977179
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_231
timestamp 1649977179
transform 1 0 22356 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_248
timestamp 1649977179
transform 1 0 23920 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_257
timestamp 1649977179
transform 1 0 24748 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_271
timestamp 1649977179
transform 1 0 26036 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1649977179
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_287
timestamp 1649977179
transform 1 0 27508 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_295
timestamp 1649977179
transform 1 0 28244 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_301
timestamp 1649977179
transform 1 0 28796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_312
timestamp 1649977179
transform 1 0 29808 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_332
timestamp 1649977179
transform 1 0 31648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_337
timestamp 1649977179
transform 1 0 32108 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_346
timestamp 1649977179
transform 1 0 32936 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_374
timestamp 1649977179
transform 1 0 35512 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_382
timestamp 1649977179
transform 1 0 36248 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_388
timestamp 1649977179
transform 1 0 36800 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_393
timestamp 1649977179
transform 1 0 37260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_403
timestamp 1649977179
transform 1 0 38180 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_411
timestamp 1649977179
transform 1 0 38916 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1649977179
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1649977179
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1649977179
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1649977179
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1649977179
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1649977179
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1649977179
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1649977179
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1649977179
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1649977179
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1649977179
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1649977179
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1649977179
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1649977179
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1649977179
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_561
timestamp 1649977179
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_573
timestamp 1649977179
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_585
timestamp 1649977179
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_597
timestamp 1649977179
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1649977179
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1649977179
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_617
timestamp 1649977179
transform 1 0 57868 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_629
timestamp 1649977179
transform 1 0 58972 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_641
timestamp 1649977179
transform 1 0 60076 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_653
timestamp 1649977179
transform 1 0 61180 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_665
timestamp 1649977179
transform 1 0 62284 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_671
timestamp 1649977179
transform 1 0 62836 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_673
timestamp 1649977179
transform 1 0 63020 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_685
timestamp 1649977179
transform 1 0 64124 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_697
timestamp 1649977179
transform 1 0 65228 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_709
timestamp 1649977179
transform 1 0 66332 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_724
timestamp 1649977179
transform 1 0 67712 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_729
timestamp 1649977179
transform 1 0 68172 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_17
timestamp 1649977179
transform 1 0 2668 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_23
timestamp 1649977179
transform 1 0 3220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_32
timestamp 1649977179
transform 1 0 4048 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_36
timestamp 1649977179
transform 1 0 4416 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_39
timestamp 1649977179
transform 1 0 4692 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_45
timestamp 1649977179
transform 1 0 5244 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_51
timestamp 1649977179
transform 1 0 5796 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_63
timestamp 1649977179
transform 1 0 6900 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_69
timestamp 1649977179
transform 1 0 7452 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_78
timestamp 1649977179
transform 1 0 8280 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_87
timestamp 1649977179
transform 1 0 9108 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_98
timestamp 1649977179
transform 1 0 10120 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_112
timestamp 1649977179
transform 1 0 11408 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_118
timestamp 1649977179
transform 1 0 11960 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_126
timestamp 1649977179
transform 1 0 12696 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1649977179
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_146
timestamp 1649977179
transform 1 0 14536 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_157
timestamp 1649977179
transform 1 0 15548 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_166
timestamp 1649977179
transform 1 0 16376 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_178
timestamp 1649977179
transform 1 0 17480 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_186
timestamp 1649977179
transform 1 0 18216 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_192
timestamp 1649977179
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_201
timestamp 1649977179
transform 1 0 19596 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_207
timestamp 1649977179
transform 1 0 20148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_219
timestamp 1649977179
transform 1 0 21252 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_223
timestamp 1649977179
transform 1 0 21620 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_231
timestamp 1649977179
transform 1 0 22356 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_243
timestamp 1649977179
transform 1 0 23460 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1649977179
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_255
timestamp 1649977179
transform 1 0 24564 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_264
timestamp 1649977179
transform 1 0 25392 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_288
timestamp 1649977179
transform 1 0 27600 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_298
timestamp 1649977179
transform 1 0 28520 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1649977179
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_316
timestamp 1649977179
transform 1 0 30176 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_328
timestamp 1649977179
transform 1 0 31280 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_334
timestamp 1649977179
transform 1 0 31832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_337
timestamp 1649977179
transform 1 0 32108 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_349
timestamp 1649977179
transform 1 0 33212 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_361
timestamp 1649977179
transform 1 0 34316 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_365
timestamp 1649977179
transform 1 0 34684 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_377
timestamp 1649977179
transform 1 0 35788 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_381
timestamp 1649977179
transform 1 0 36156 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_392
timestamp 1649977179
transform 1 0 37168 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_396
timestamp 1649977179
transform 1 0 37536 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_405
timestamp 1649977179
transform 1 0 38364 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_411
timestamp 1649977179
transform 1 0 38916 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1649977179
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_437
timestamp 1649977179
transform 1 0 41308 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_449
timestamp 1649977179
transform 1 0 42412 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_461
timestamp 1649977179
transform 1 0 43516 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_473
timestamp 1649977179
transform 1 0 44620 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1649977179
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1649977179
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1649977179
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1649977179
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1649977179
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1649977179
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1649977179
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1649977179
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_557
timestamp 1649977179
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_569
timestamp 1649977179
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1649977179
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1649977179
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_589
timestamp 1649977179
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_601
timestamp 1649977179
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_613
timestamp 1649977179
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_625
timestamp 1649977179
transform 1 0 58604 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_637
timestamp 1649977179
transform 1 0 59708 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_643
timestamp 1649977179
transform 1 0 60260 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_645
timestamp 1649977179
transform 1 0 60444 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_657
timestamp 1649977179
transform 1 0 61548 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_669
timestamp 1649977179
transform 1 0 62652 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_681
timestamp 1649977179
transform 1 0 63756 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_693
timestamp 1649977179
transform 1 0 64860 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_699
timestamp 1649977179
transform 1 0 65412 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_701
timestamp 1649977179
transform 1 0 65596 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_713
timestamp 1649977179
transform 1 0 66700 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_725
timestamp 1649977179
transform 1 0 67804 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_7
timestamp 1649977179
transform 1 0 1748 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_18
timestamp 1649977179
transform 1 0 2760 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_38
timestamp 1649977179
transform 1 0 4600 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_46
timestamp 1649977179
transform 1 0 5336 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_52
timestamp 1649977179
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_61
timestamp 1649977179
transform 1 0 6716 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_75
timestamp 1649977179
transform 1 0 8004 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_95
timestamp 1649977179
transform 1 0 9844 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_106
timestamp 1649977179
transform 1 0 10856 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_120
timestamp 1649977179
transform 1 0 12144 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_124
timestamp 1649977179
transform 1 0 12512 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_130
timestamp 1649977179
transform 1 0 13064 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_138
timestamp 1649977179
transform 1 0 13800 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_144
timestamp 1649977179
transform 1 0 14352 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_152
timestamp 1649977179
transform 1 0 15088 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_160
timestamp 1649977179
transform 1 0 15824 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_180
timestamp 1649977179
transform 1 0 17664 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_192
timestamp 1649977179
transform 1 0 18768 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_198
timestamp 1649977179
transform 1 0 19320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_207
timestamp 1649977179
transform 1 0 20148 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_216
timestamp 1649977179
transform 1 0 20976 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_232
timestamp 1649977179
transform 1 0 22448 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_244
timestamp 1649977179
transform 1 0 23552 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_251
timestamp 1649977179
transform 1 0 24196 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_260
timestamp 1649977179
transform 1 0 25024 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_272
timestamp 1649977179
transform 1 0 26128 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_288
timestamp 1649977179
transform 1 0 27600 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_294
timestamp 1649977179
transform 1 0 28152 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_300
timestamp 1649977179
transform 1 0 28704 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_311
timestamp 1649977179
transform 1 0 29716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_323
timestamp 1649977179
transform 1 0 30820 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1649977179
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_337
timestamp 1649977179
transform 1 0 32108 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_343
timestamp 1649977179
transform 1 0 32660 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_355
timestamp 1649977179
transform 1 0 33764 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_369
timestamp 1649977179
transform 1 0 35052 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_373
timestamp 1649977179
transform 1 0 35420 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_379
timestamp 1649977179
transform 1 0 35972 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1649977179
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_403
timestamp 1649977179
transform 1 0 38180 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_412
timestamp 1649977179
transform 1 0 39008 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_420
timestamp 1649977179
transform 1 0 39744 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_437
timestamp 1649977179
transform 1 0 41308 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_445
timestamp 1649977179
transform 1 0 42044 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1649977179
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1649977179
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1649977179
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1649977179
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1649977179
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1649977179
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1649977179
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1649977179
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1649977179
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1649977179
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1649977179
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1649977179
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_561
timestamp 1649977179
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_573
timestamp 1649977179
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_585
timestamp 1649977179
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_597
timestamp 1649977179
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1649977179
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1649977179
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_617
timestamp 1649977179
transform 1 0 57868 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_629
timestamp 1649977179
transform 1 0 58972 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_641
timestamp 1649977179
transform 1 0 60076 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_653
timestamp 1649977179
transform 1 0 61180 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_665
timestamp 1649977179
transform 1 0 62284 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_671
timestamp 1649977179
transform 1 0 62836 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_673
timestamp 1649977179
transform 1 0 63020 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_685
timestamp 1649977179
transform 1 0 64124 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_697
timestamp 1649977179
transform 1 0 65228 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_709
timestamp 1649977179
transform 1 0 66332 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_721
timestamp 1649977179
transform 1 0 67436 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_727
timestamp 1649977179
transform 1 0 67988 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_729
timestamp 1649977179
transform 1 0 68172 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_9
timestamp 1649977179
transform 1 0 1932 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_21
timestamp 1649977179
transform 1 0 3036 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_33
timestamp 1649977179
transform 1 0 4140 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_39
timestamp 1649977179
transform 1 0 4692 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_59
timestamp 1649977179
transform 1 0 6532 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_69
timestamp 1649977179
transform 1 0 7452 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_73
timestamp 1649977179
transform 1 0 7820 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_79
timestamp 1649977179
transform 1 0 8372 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_92
timestamp 1649977179
transform 1 0 9568 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_106
timestamp 1649977179
transform 1 0 10856 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_112
timestamp 1649977179
transform 1 0 11408 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_120
timestamp 1649977179
transform 1 0 12144 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_126
timestamp 1649977179
transform 1 0 12696 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_136
timestamp 1649977179
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_147
timestamp 1649977179
transform 1 0 14628 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_159
timestamp 1649977179
transform 1 0 15732 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_171
timestamp 1649977179
transform 1 0 16836 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_177
timestamp 1649977179
transform 1 0 17388 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_191
timestamp 1649977179
transform 1 0 18676 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1649977179
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_202
timestamp 1649977179
transform 1 0 19688 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_210
timestamp 1649977179
transform 1 0 20424 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_213
timestamp 1649977179
transform 1 0 20700 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_227
timestamp 1649977179
transform 1 0 21988 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_244
timestamp 1649977179
transform 1 0 23552 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_267
timestamp 1649977179
transform 1 0 25668 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_289
timestamp 1649977179
transform 1 0 27692 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_304
timestamp 1649977179
transform 1 0 29072 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_316
timestamp 1649977179
transform 1 0 30176 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_336
timestamp 1649977179
transform 1 0 32016 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_360
timestamp 1649977179
transform 1 0 34224 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_365
timestamp 1649977179
transform 1 0 34684 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_368
timestamp 1649977179
transform 1 0 34960 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_380
timestamp 1649977179
transform 1 0 36064 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_392
timestamp 1649977179
transform 1 0 37168 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_395
timestamp 1649977179
transform 1 0 37444 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_407
timestamp 1649977179
transform 1 0 38548 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_413
timestamp 1649977179
transform 1 0 39100 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_416
timestamp 1649977179
transform 1 0 39376 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_421
timestamp 1649977179
transform 1 0 39836 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1649977179
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1649977179
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1649977179
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1649977179
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1649977179
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1649977179
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1649977179
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1649977179
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1649977179
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1649977179
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_533
timestamp 1649977179
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_545
timestamp 1649977179
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_557
timestamp 1649977179
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_569
timestamp 1649977179
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1649977179
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1649977179
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_589
timestamp 1649977179
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_601
timestamp 1649977179
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_613
timestamp 1649977179
transform 1 0 57500 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_625
timestamp 1649977179
transform 1 0 58604 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_637
timestamp 1649977179
transform 1 0 59708 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_643
timestamp 1649977179
transform 1 0 60260 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_645
timestamp 1649977179
transform 1 0 60444 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_657
timestamp 1649977179
transform 1 0 61548 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_669
timestamp 1649977179
transform 1 0 62652 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_681
timestamp 1649977179
transform 1 0 63756 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_693
timestamp 1649977179
transform 1 0 64860 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_699
timestamp 1649977179
transform 1 0 65412 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_701
timestamp 1649977179
transform 1 0 65596 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_713
timestamp 1649977179
transform 1 0 66700 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_725
timestamp 1649977179
transform 1 0 67804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_729
timestamp 1649977179
transform 1 0 68172 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_13
timestamp 1649977179
transform 1 0 2300 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_33
timestamp 1649977179
transform 1 0 4140 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_47
timestamp 1649977179
transform 1 0 5428 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_62
timestamp 1649977179
transform 1 0 6808 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_71
timestamp 1649977179
transform 1 0 7636 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_75
timestamp 1649977179
transform 1 0 8004 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_86
timestamp 1649977179
transform 1 0 9016 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_106
timestamp 1649977179
transform 1 0 10856 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_121
timestamp 1649977179
transform 1 0 12236 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_129
timestamp 1649977179
transform 1 0 12972 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_134
timestamp 1649977179
transform 1 0 13432 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_142
timestamp 1649977179
transform 1 0 14168 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_150
timestamp 1649977179
transform 1 0 14904 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_156
timestamp 1649977179
transform 1 0 15456 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_162
timestamp 1649977179
transform 1 0 16008 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_174
timestamp 1649977179
transform 1 0 17112 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_182
timestamp 1649977179
transform 1 0 17848 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_200
timestamp 1649977179
transform 1 0 19504 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_220
timestamp 1649977179
transform 1 0 21344 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_225
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_233
timestamp 1649977179
transform 1 0 22540 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_239
timestamp 1649977179
transform 1 0 23092 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_243
timestamp 1649977179
transform 1 0 23460 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_250
timestamp 1649977179
transform 1 0 24104 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_256
timestamp 1649977179
transform 1 0 24656 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_265
timestamp 1649977179
transform 1 0 25484 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_271
timestamp 1649977179
transform 1 0 26036 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1649977179
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_283
timestamp 1649977179
transform 1 0 27140 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_289
timestamp 1649977179
transform 1 0 27692 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_297
timestamp 1649977179
transform 1 0 28428 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_311
timestamp 1649977179
transform 1 0 29716 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_319
timestamp 1649977179
transform 1 0 30452 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_323
timestamp 1649977179
transform 1 0 30820 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_332
timestamp 1649977179
transform 1 0 31648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_337
timestamp 1649977179
transform 1 0 32108 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_348
timestamp 1649977179
transform 1 0 33120 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_352
timestamp 1649977179
transform 1 0 33488 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_357
timestamp 1649977179
transform 1 0 33948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_361
timestamp 1649977179
transform 1 0 34316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_367
timestamp 1649977179
transform 1 0 34868 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_387
timestamp 1649977179
transform 1 0 36708 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1649977179
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_393
timestamp 1649977179
transform 1 0 37260 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_399
timestamp 1649977179
transform 1 0 37812 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_427
timestamp 1649977179
transform 1 0 40388 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_439
timestamp 1649977179
transform 1 0 41492 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1649977179
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1649977179
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1649977179
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1649977179
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1649977179
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1649977179
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1649977179
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1649977179
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1649977179
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_529
timestamp 1649977179
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1649977179
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1649977179
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1649977179
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_561
timestamp 1649977179
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_573
timestamp 1649977179
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_585
timestamp 1649977179
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_597
timestamp 1649977179
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1649977179
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1649977179
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_617
timestamp 1649977179
transform 1 0 57868 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_629
timestamp 1649977179
transform 1 0 58972 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_641
timestamp 1649977179
transform 1 0 60076 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_653
timestamp 1649977179
transform 1 0 61180 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_665
timestamp 1649977179
transform 1 0 62284 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_671
timestamp 1649977179
transform 1 0 62836 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_673
timestamp 1649977179
transform 1 0 63020 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_685
timestamp 1649977179
transform 1 0 64124 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_697
timestamp 1649977179
transform 1 0 65228 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_709
timestamp 1649977179
transform 1 0 66332 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_721
timestamp 1649977179
transform 1 0 67436 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_727
timestamp 1649977179
transform 1 0 67988 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_729
timestamp 1649977179
transform 1 0 68172 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_21
timestamp 1649977179
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_39
timestamp 1649977179
transform 1 0 4692 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_51
timestamp 1649977179
transform 1 0 5796 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_59
timestamp 1649977179
transform 1 0 6532 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_68
timestamp 1649977179
transform 1 0 7360 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_80
timestamp 1649977179
transform 1 0 8464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_90
timestamp 1649977179
transform 1 0 9384 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_96
timestamp 1649977179
transform 1 0 9936 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_102
timestamp 1649977179
transform 1 0 10488 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_119
timestamp 1649977179
transform 1 0 12052 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_129
timestamp 1649977179
transform 1 0 12972 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_135
timestamp 1649977179
transform 1 0 13524 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_144
timestamp 1649977179
transform 1 0 14352 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_148
timestamp 1649977179
transform 1 0 14720 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_156
timestamp 1649977179
transform 1 0 15456 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_168
timestamp 1649977179
transform 1 0 16560 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_179
timestamp 1649977179
transform 1 0 17572 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_191
timestamp 1649977179
transform 1 0 18676 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_205
timestamp 1649977179
transform 1 0 19964 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_209
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_217
timestamp 1649977179
transform 1 0 21068 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_225
timestamp 1649977179
transform 1 0 21804 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1649977179
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1649977179
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1649977179
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_253
timestamp 1649977179
transform 1 0 24380 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_256
timestamp 1649977179
transform 1 0 24656 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_268
timestamp 1649977179
transform 1 0 25760 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_274
timestamp 1649977179
transform 1 0 26312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_280
timestamp 1649977179
transform 1 0 26864 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_288
timestamp 1649977179
transform 1 0 27600 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_298
timestamp 1649977179
transform 1 0 28520 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_304
timestamp 1649977179
transform 1 0 29072 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_314
timestamp 1649977179
transform 1 0 29992 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_320
timestamp 1649977179
transform 1 0 30544 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_328
timestamp 1649977179
transform 1 0 31280 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_342
timestamp 1649977179
transform 1 0 32568 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_348
timestamp 1649977179
transform 1 0 33120 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_356
timestamp 1649977179
transform 1 0 33856 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_360
timestamp 1649977179
transform 1 0 34224 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_365
timestamp 1649977179
transform 1 0 34684 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_389
timestamp 1649977179
transform 1 0 36892 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_405
timestamp 1649977179
transform 1 0 38364 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_414
timestamp 1649977179
transform 1 0 39192 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1649977179
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1649977179
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1649977179
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1649977179
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1649977179
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1649977179
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1649977179
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1649977179
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1649977179
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1649977179
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1649977179
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1649977179
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_533
timestamp 1649977179
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_545
timestamp 1649977179
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_557
timestamp 1649977179
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_569
timestamp 1649977179
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1649977179
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1649977179
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_589
timestamp 1649977179
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_601
timestamp 1649977179
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_613
timestamp 1649977179
transform 1 0 57500 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_625
timestamp 1649977179
transform 1 0 58604 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_637
timestamp 1649977179
transform 1 0 59708 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_643
timestamp 1649977179
transform 1 0 60260 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_645
timestamp 1649977179
transform 1 0 60444 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_657
timestamp 1649977179
transform 1 0 61548 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_669
timestamp 1649977179
transform 1 0 62652 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_681
timestamp 1649977179
transform 1 0 63756 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_693
timestamp 1649977179
transform 1 0 64860 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_699
timestamp 1649977179
transform 1 0 65412 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_701
timestamp 1649977179
transform 1 0 65596 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_713
timestamp 1649977179
transform 1 0 66700 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_725
timestamp 1649977179
transform 1 0 67804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_729
timestamp 1649977179
transform 1 0 68172 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_12
timestamp 1649977179
transform 1 0 2208 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_24
timestamp 1649977179
transform 1 0 3312 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_36
timestamp 1649977179
transform 1 0 4416 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_42
timestamp 1649977179
transform 1 0 4968 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_50
timestamp 1649977179
transform 1 0 5704 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_101
timestamp 1649977179
transform 1 0 10396 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_109
timestamp 1649977179
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_120
timestamp 1649977179
transform 1 0 12144 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_140
timestamp 1649977179
transform 1 0 13984 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_164
timestamp 1649977179
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_185
timestamp 1649977179
transform 1 0 18124 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_197
timestamp 1649977179
transform 1 0 19228 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_209
timestamp 1649977179
transform 1 0 20332 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1649977179
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_233
timestamp 1649977179
transform 1 0 22540 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_253
timestamp 1649977179
transform 1 0 24380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_261
timestamp 1649977179
transform 1 0 25116 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1649977179
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1649977179
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_297
timestamp 1649977179
transform 1 0 28428 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_303
timestamp 1649977179
transform 1 0 28980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_317
timestamp 1649977179
transform 1 0 30268 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_324
timestamp 1649977179
transform 1 0 30912 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_332
timestamp 1649977179
transform 1 0 31648 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_342
timestamp 1649977179
transform 1 0 32568 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_346
timestamp 1649977179
transform 1 0 32936 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_363
timestamp 1649977179
transform 1 0 34500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_374
timestamp 1649977179
transform 1 0 35512 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1649977179
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1649977179
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_395
timestamp 1649977179
transform 1 0 37444 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_401
timestamp 1649977179
transform 1 0 37996 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_413
timestamp 1649977179
transform 1 0 39100 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_425
timestamp 1649977179
transform 1 0 40204 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_437
timestamp 1649977179
transform 1 0 41308 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_445
timestamp 1649977179
transform 1 0 42044 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1649977179
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1649977179
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1649977179
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1649977179
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1649977179
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1649977179
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1649977179
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_517
timestamp 1649977179
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_529
timestamp 1649977179
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_541
timestamp 1649977179
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1649977179
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1649977179
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_561
timestamp 1649977179
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_573
timestamp 1649977179
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_585
timestamp 1649977179
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_597
timestamp 1649977179
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1649977179
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1649977179
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_617
timestamp 1649977179
transform 1 0 57868 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_629
timestamp 1649977179
transform 1 0 58972 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_641
timestamp 1649977179
transform 1 0 60076 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_653
timestamp 1649977179
transform 1 0 61180 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_665
timestamp 1649977179
transform 1 0 62284 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_671
timestamp 1649977179
transform 1 0 62836 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_673
timestamp 1649977179
transform 1 0 63020 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_685
timestamp 1649977179
transform 1 0 64124 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_697
timestamp 1649977179
transform 1 0 65228 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_709
timestamp 1649977179
transform 1 0 66332 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_721
timestamp 1649977179
transform 1 0 67436 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_727
timestamp 1649977179
transform 1 0 67988 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_729
timestamp 1649977179
transform 1 0 68172 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1649977179
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_13
timestamp 1649977179
transform 1 0 2300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_25
timestamp 1649977179
transform 1 0 3404 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_45
timestamp 1649977179
transform 1 0 5244 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_59
timestamp 1649977179
transform 1 0 6532 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_66
timestamp 1649977179
transform 1 0 7176 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_80
timestamp 1649977179
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_88
timestamp 1649977179
transform 1 0 9200 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_100
timestamp 1649977179
transform 1 0 10304 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_149
timestamp 1649977179
transform 1 0 14812 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_157
timestamp 1649977179
transform 1 0 15548 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_162
timestamp 1649977179
transform 1 0 16008 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_168
timestamp 1649977179
transform 1 0 16560 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1649977179
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_207
timestamp 1649977179
transform 1 0 20148 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_231
timestamp 1649977179
transform 1 0 22356 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_243
timestamp 1649977179
transform 1 0 23460 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1649977179
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_253
timestamp 1649977179
transform 1 0 24380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_257
timestamp 1649977179
transform 1 0 24748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_263
timestamp 1649977179
transform 1 0 25300 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_272
timestamp 1649977179
transform 1 0 26128 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_24_286
timestamp 1649977179
transform 1 0 27416 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_292
timestamp 1649977179
transform 1 0 27968 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_300
timestamp 1649977179
transform 1 0 28704 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_311
timestamp 1649977179
transform 1 0 29716 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_315
timestamp 1649977179
transform 1 0 30084 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_332
timestamp 1649977179
transform 1 0 31648 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_338
timestamp 1649977179
transform 1 0 32200 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_350
timestamp 1649977179
transform 1 0 33304 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_356
timestamp 1649977179
transform 1 0 33856 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_365
timestamp 1649977179
transform 1 0 34684 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_380
timestamp 1649977179
transform 1 0 36064 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_384
timestamp 1649977179
transform 1 0 36432 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_390
timestamp 1649977179
transform 1 0 36984 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_402
timestamp 1649977179
transform 1 0 38088 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_411
timestamp 1649977179
transform 1 0 38916 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1649977179
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_437
timestamp 1649977179
transform 1 0 41308 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_449
timestamp 1649977179
transform 1 0 42412 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_461
timestamp 1649977179
transform 1 0 43516 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_473
timestamp 1649977179
transform 1 0 44620 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1649977179
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1649977179
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1649977179
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1649977179
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1649977179
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1649977179
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_533
timestamp 1649977179
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_545
timestamp 1649977179
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_557
timestamp 1649977179
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_569
timestamp 1649977179
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1649977179
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1649977179
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_589
timestamp 1649977179
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_601
timestamp 1649977179
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_613
timestamp 1649977179
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_625
timestamp 1649977179
transform 1 0 58604 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_637
timestamp 1649977179
transform 1 0 59708 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_643
timestamp 1649977179
transform 1 0 60260 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_645
timestamp 1649977179
transform 1 0 60444 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_657
timestamp 1649977179
transform 1 0 61548 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_669
timestamp 1649977179
transform 1 0 62652 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_681
timestamp 1649977179
transform 1 0 63756 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_693
timestamp 1649977179
transform 1 0 64860 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_699
timestamp 1649977179
transform 1 0 65412 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_701
timestamp 1649977179
transform 1 0 65596 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_713
timestamp 1649977179
transform 1 0 66700 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_725
timestamp 1649977179
transform 1 0 67804 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_9
timestamp 1649977179
transform 1 0 1932 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_18
timestamp 1649977179
transform 1 0 2760 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_24
timestamp 1649977179
transform 1 0 3312 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_36
timestamp 1649977179
transform 1 0 4416 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_40
timestamp 1649977179
transform 1 0 4784 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_48
timestamp 1649977179
transform 1 0 5520 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_60
timestamp 1649977179
transform 1 0 6624 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_71
timestamp 1649977179
transform 1 0 7636 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_77
timestamp 1649977179
transform 1 0 8188 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_83
timestamp 1649977179
transform 1 0 8740 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_95
timestamp 1649977179
transform 1 0 9844 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_107
timestamp 1649977179
transform 1 0 10948 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_121
timestamp 1649977179
transform 1 0 12236 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_130
timestamp 1649977179
transform 1 0 13064 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_136
timestamp 1649977179
transform 1 0 13616 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_142
timestamp 1649977179
transform 1 0 14168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_145
timestamp 1649977179
transform 1 0 14444 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_158
timestamp 1649977179
transform 1 0 15640 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1649977179
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_174
timestamp 1649977179
transform 1 0 17112 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_184
timestamp 1649977179
transform 1 0 18032 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_196
timestamp 1649977179
transform 1 0 19136 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_200
timestamp 1649977179
transform 1 0 19504 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_209
timestamp 1649977179
transform 1 0 20332 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_220
timestamp 1649977179
transform 1 0 21344 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_227
timestamp 1649977179
transform 1 0 21988 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_239
timestamp 1649977179
transform 1 0 23092 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_242
timestamp 1649977179
transform 1 0 23368 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_250
timestamp 1649977179
transform 1 0 24104 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_259
timestamp 1649977179
transform 1 0 24932 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_267
timestamp 1649977179
transform 1 0 25668 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_276
timestamp 1649977179
transform 1 0 26496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_281
timestamp 1649977179
transform 1 0 26956 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_295
timestamp 1649977179
transform 1 0 28244 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_319
timestamp 1649977179
transform 1 0 30452 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_330
timestamp 1649977179
transform 1 0 31464 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1649977179
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_347
timestamp 1649977179
transform 1 0 33028 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_355
timestamp 1649977179
transform 1 0 33764 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_364
timestamp 1649977179
transform 1 0 34592 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_379
timestamp 1649977179
transform 1 0 35972 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_385
timestamp 1649977179
transform 1 0 36524 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_388
timestamp 1649977179
transform 1 0 36800 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_393
timestamp 1649977179
transform 1 0 37260 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_397
timestamp 1649977179
transform 1 0 37628 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_406
timestamp 1649977179
transform 1 0 38456 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_430
timestamp 1649977179
transform 1 0 40664 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_442
timestamp 1649977179
transform 1 0 41768 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1649977179
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1649977179
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1649977179
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1649977179
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1649977179
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1649977179
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1649977179
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_517
timestamp 1649977179
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_529
timestamp 1649977179
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_541
timestamp 1649977179
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1649977179
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1649977179
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_561
timestamp 1649977179
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_573
timestamp 1649977179
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_585
timestamp 1649977179
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_597
timestamp 1649977179
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1649977179
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1649977179
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_617
timestamp 1649977179
transform 1 0 57868 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_629
timestamp 1649977179
transform 1 0 58972 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_641
timestamp 1649977179
transform 1 0 60076 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_653
timestamp 1649977179
transform 1 0 61180 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_665
timestamp 1649977179
transform 1 0 62284 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_671
timestamp 1649977179
transform 1 0 62836 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_673
timestamp 1649977179
transform 1 0 63020 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_685
timestamp 1649977179
transform 1 0 64124 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_697
timestamp 1649977179
transform 1 0 65228 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_709
timestamp 1649977179
transform 1 0 66332 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_724
timestamp 1649977179
transform 1 0 67712 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_729
timestamp 1649977179
transform 1 0 68172 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_9
timestamp 1649977179
transform 1 0 1932 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_18
timestamp 1649977179
transform 1 0 2760 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1649977179
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_45
timestamp 1649977179
transform 1 0 5244 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_49
timestamp 1649977179
transform 1 0 5612 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_54
timestamp 1649977179
transform 1 0 6072 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_65
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_74
timestamp 1649977179
transform 1 0 7912 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1649977179
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_107
timestamp 1649977179
transform 1 0 10948 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_113
timestamp 1649977179
transform 1 0 11500 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_121
timestamp 1649977179
transform 1 0 12236 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_132
timestamp 1649977179
transform 1 0 13248 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_157
timestamp 1649977179
transform 1 0 15548 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_163
timestamp 1649977179
transform 1 0 16100 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_175
timestamp 1649977179
transform 1 0 17204 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_183
timestamp 1649977179
transform 1 0 17940 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1649977179
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_202
timestamp 1649977179
transform 1 0 19688 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_212
timestamp 1649977179
transform 1 0 20608 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_220
timestamp 1649977179
transform 1 0 21344 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_229
timestamp 1649977179
transform 1 0 22172 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_241
timestamp 1649977179
transform 1 0 23276 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_245
timestamp 1649977179
transform 1 0 23644 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_248
timestamp 1649977179
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_269
timestamp 1649977179
transform 1 0 25852 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_275
timestamp 1649977179
transform 1 0 26404 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_299
timestamp 1649977179
transform 1 0 28612 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1649977179
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_319
timestamp 1649977179
transform 1 0 30452 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_330
timestamp 1649977179
transform 1 0 31464 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_348
timestamp 1649977179
transform 1 0 33120 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1649977179
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1649977179
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_367
timestamp 1649977179
transform 1 0 34868 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_387
timestamp 1649977179
transform 1 0 36708 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_395
timestamp 1649977179
transform 1 0 37444 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_403
timestamp 1649977179
transform 1 0 38180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_415
timestamp 1649977179
transform 1 0 39284 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1649977179
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1649977179
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1649977179
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1649977179
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1649977179
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1649977179
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1649977179
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1649977179
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1649977179
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1649977179
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_513
timestamp 1649977179
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1649977179
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1649977179
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_533
timestamp 1649977179
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_545
timestamp 1649977179
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_557
timestamp 1649977179
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_569
timestamp 1649977179
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1649977179
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1649977179
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_589
timestamp 1649977179
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_601
timestamp 1649977179
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_613
timestamp 1649977179
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_625
timestamp 1649977179
transform 1 0 58604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_637
timestamp 1649977179
transform 1 0 59708 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_643
timestamp 1649977179
transform 1 0 60260 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_645
timestamp 1649977179
transform 1 0 60444 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_657
timestamp 1649977179
transform 1 0 61548 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_669
timestamp 1649977179
transform 1 0 62652 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_681
timestamp 1649977179
transform 1 0 63756 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_693
timestamp 1649977179
transform 1 0 64860 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_699
timestamp 1649977179
transform 1 0 65412 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_701
timestamp 1649977179
transform 1 0 65596 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_713
timestamp 1649977179
transform 1 0 66700 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_725
timestamp 1649977179
transform 1 0 67804 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1649977179
transform 1 0 1748 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_13
timestamp 1649977179
transform 1 0 2300 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_25
timestamp 1649977179
transform 1 0 3404 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_37
timestamp 1649977179
transform 1 0 4508 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_40
timestamp 1649977179
transform 1 0 4784 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1649977179
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_62
timestamp 1649977179
transform 1 0 6808 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_74
timestamp 1649977179
transform 1 0 7912 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_94
timestamp 1649977179
transform 1 0 9752 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_107
timestamp 1649977179
transform 1 0 10948 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_129
timestamp 1649977179
transform 1 0 12972 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_141
timestamp 1649977179
transform 1 0 14076 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_147
timestamp 1649977179
transform 1 0 14628 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_153
timestamp 1649977179
transform 1 0 15180 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1649977179
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_174
timestamp 1649977179
transform 1 0 17112 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_180
timestamp 1649977179
transform 1 0 17664 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_192
timestamp 1649977179
transform 1 0 18768 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_200
timestamp 1649977179
transform 1 0 19504 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_208
timestamp 1649977179
transform 1 0 20240 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_218
timestamp 1649977179
transform 1 0 21160 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_225
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_245
timestamp 1649977179
transform 1 0 23644 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_257
timestamp 1649977179
transform 1 0 24748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_266
timestamp 1649977179
transform 1 0 25576 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_276
timestamp 1649977179
transform 1 0 26496 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_281
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_293
timestamp 1649977179
transform 1 0 28060 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_302
timestamp 1649977179
transform 1 0 28888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_306
timestamp 1649977179
transform 1 0 29256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_314
timestamp 1649977179
transform 1 0 29992 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_322
timestamp 1649977179
transform 1 0 30728 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_331
timestamp 1649977179
transform 1 0 31556 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1649977179
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_342
timestamp 1649977179
transform 1 0 32568 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_346
timestamp 1649977179
transform 1 0 32936 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_363
timestamp 1649977179
transform 1 0 34500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_381
timestamp 1649977179
transform 1 0 36156 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_389
timestamp 1649977179
transform 1 0 36892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_395
timestamp 1649977179
transform 1 0 37444 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_407
timestamp 1649977179
transform 1 0 38548 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_413
timestamp 1649977179
transform 1 0 39100 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_430
timestamp 1649977179
transform 1 0 40664 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_442
timestamp 1649977179
transform 1 0 41768 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1649977179
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1649977179
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1649977179
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1649977179
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1649977179
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1649977179
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1649977179
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_517
timestamp 1649977179
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_529
timestamp 1649977179
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_541
timestamp 1649977179
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1649977179
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1649977179
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_561
timestamp 1649977179
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_573
timestamp 1649977179
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_585
timestamp 1649977179
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_597
timestamp 1649977179
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1649977179
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1649977179
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_617
timestamp 1649977179
transform 1 0 57868 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_629
timestamp 1649977179
transform 1 0 58972 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_641
timestamp 1649977179
transform 1 0 60076 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_653
timestamp 1649977179
transform 1 0 61180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_665
timestamp 1649977179
transform 1 0 62284 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_671
timestamp 1649977179
transform 1 0 62836 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_673
timestamp 1649977179
transform 1 0 63020 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_685
timestamp 1649977179
transform 1 0 64124 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_697
timestamp 1649977179
transform 1 0 65228 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_709
timestamp 1649977179
transform 1 0 66332 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_724
timestamp 1649977179
transform 1 0 67712 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_729
timestamp 1649977179
transform 1 0 68172 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_15
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_18
timestamp 1649977179
transform 1 0 2760 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1649977179
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_38
timestamp 1649977179
transform 1 0 4600 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_50
timestamp 1649977179
transform 1 0 5704 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_56
timestamp 1649977179
transform 1 0 6256 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_74
timestamp 1649977179
transform 1 0 7912 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_80
timestamp 1649977179
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_89
timestamp 1649977179
transform 1 0 9292 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_98
timestamp 1649977179
transform 1 0 10120 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_110
timestamp 1649977179
transform 1 0 11224 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_113
timestamp 1649977179
transform 1 0 11500 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_125
timestamp 1649977179
transform 1 0 12604 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_132
timestamp 1649977179
transform 1 0 13248 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_145
timestamp 1649977179
transform 1 0 14444 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_162
timestamp 1649977179
transform 1 0 16008 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_176
timestamp 1649977179
transform 1 0 17296 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_184
timestamp 1649977179
transform 1 0 18032 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1649977179
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_203
timestamp 1649977179
transform 1 0 19780 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1649977179
transform 1 0 20884 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1649977179
transform 1 0 21252 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_222
timestamp 1649977179
transform 1 0 21528 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_246
timestamp 1649977179
transform 1 0 23736 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_258
timestamp 1649977179
transform 1 0 24840 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_264
timestamp 1649977179
transform 1 0 25392 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_272
timestamp 1649977179
transform 1 0 26128 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_292
timestamp 1649977179
transform 1 0 27968 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_300
timestamp 1649977179
transform 1 0 28704 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_304
timestamp 1649977179
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_309
timestamp 1649977179
transform 1 0 29532 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_320
timestamp 1649977179
transform 1 0 30544 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_329
timestamp 1649977179
transform 1 0 31372 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_345
timestamp 1649977179
transform 1 0 32844 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1649977179
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1649977179
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_365
timestamp 1649977179
transform 1 0 34684 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_368
timestamp 1649977179
transform 1 0 34960 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_380
timestamp 1649977179
transform 1 0 36064 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_389
timestamp 1649977179
transform 1 0 36892 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_395
timestamp 1649977179
transform 1 0 37444 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_407
timestamp 1649977179
transform 1 0 38548 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_416
timestamp 1649977179
transform 1 0 39376 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1649977179
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1649977179
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1649977179
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1649977179
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1649977179
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1649977179
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1649977179
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1649977179
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1649977179
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1649977179
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1649977179
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1649977179
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_533
timestamp 1649977179
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_545
timestamp 1649977179
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_557
timestamp 1649977179
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_569
timestamp 1649977179
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1649977179
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1649977179
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_589
timestamp 1649977179
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_601
timestamp 1649977179
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_613
timestamp 1649977179
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_625
timestamp 1649977179
transform 1 0 58604 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_637
timestamp 1649977179
transform 1 0 59708 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_643
timestamp 1649977179
transform 1 0 60260 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_645
timestamp 1649977179
transform 1 0 60444 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_657
timestamp 1649977179
transform 1 0 61548 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_669
timestamp 1649977179
transform 1 0 62652 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_681
timestamp 1649977179
transform 1 0 63756 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_693
timestamp 1649977179
transform 1 0 64860 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_699
timestamp 1649977179
transform 1 0 65412 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_701
timestamp 1649977179
transform 1 0 65596 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_713
timestamp 1649977179
transform 1 0 66700 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_725
timestamp 1649977179
transform 1 0 67804 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_7
timestamp 1649977179
transform 1 0 1748 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_16
timestamp 1649977179
transform 1 0 2576 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_36
timestamp 1649977179
transform 1 0 4416 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_48
timestamp 1649977179
transform 1 0 5520 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_73
timestamp 1649977179
transform 1 0 7820 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_80
timestamp 1649977179
transform 1 0 8464 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_89
timestamp 1649977179
transform 1 0 9292 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_103
timestamp 1649977179
transform 1 0 10580 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_121
timestamp 1649977179
transform 1 0 12236 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_125
timestamp 1649977179
transform 1 0 12604 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_142
timestamp 1649977179
transform 1 0 14168 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_154
timestamp 1649977179
transform 1 0 15272 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1649977179
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_181
timestamp 1649977179
transform 1 0 17756 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_187
timestamp 1649977179
transform 1 0 18308 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_198
timestamp 1649977179
transform 1 0 19320 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_204
timestamp 1649977179
transform 1 0 19872 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_213
timestamp 1649977179
transform 1 0 20700 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1649977179
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_230
timestamp 1649977179
transform 1 0 22264 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_254
timestamp 1649977179
transform 1 0 24472 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_262
timestamp 1649977179
transform 1 0 25208 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_275
timestamp 1649977179
transform 1 0 26404 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1649977179
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_281
timestamp 1649977179
transform 1 0 26956 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_291
timestamp 1649977179
transform 1 0 27876 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_297
timestamp 1649977179
transform 1 0 28428 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_306
timestamp 1649977179
transform 1 0 29256 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_313
timestamp 1649977179
transform 1 0 29900 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_319
timestamp 1649977179
transform 1 0 30452 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_328
timestamp 1649977179
transform 1 0 31280 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_340
timestamp 1649977179
transform 1 0 32384 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_354
timestamp 1649977179
transform 1 0 33672 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_363
timestamp 1649977179
transform 1 0 34500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_371
timestamp 1649977179
transform 1 0 35236 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_388
timestamp 1649977179
transform 1 0 36800 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_393
timestamp 1649977179
transform 1 0 37260 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_397
timestamp 1649977179
transform 1 0 37628 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_403
timestamp 1649977179
transform 1 0 38180 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_411
timestamp 1649977179
transform 1 0 38916 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_428
timestamp 1649977179
transform 1 0 40480 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_440
timestamp 1649977179
transform 1 0 41584 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1649977179
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1649977179
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1649977179
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1649977179
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1649977179
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1649977179
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1649977179
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_517
timestamp 1649977179
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_529
timestamp 1649977179
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_541
timestamp 1649977179
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1649977179
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1649977179
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_561
timestamp 1649977179
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_573
timestamp 1649977179
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_585
timestamp 1649977179
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_597
timestamp 1649977179
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1649977179
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1649977179
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_617
timestamp 1649977179
transform 1 0 57868 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_629
timestamp 1649977179
transform 1 0 58972 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_641
timestamp 1649977179
transform 1 0 60076 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_653
timestamp 1649977179
transform 1 0 61180 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_665
timestamp 1649977179
transform 1 0 62284 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_671
timestamp 1649977179
transform 1 0 62836 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_673
timestamp 1649977179
transform 1 0 63020 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_685
timestamp 1649977179
transform 1 0 64124 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_697
timestamp 1649977179
transform 1 0 65228 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_709
timestamp 1649977179
transform 1 0 66332 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_721
timestamp 1649977179
transform 1 0 67436 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_727
timestamp 1649977179
transform 1 0 67988 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_729
timestamp 1649977179
transform 1 0 68172 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_16
timestamp 1649977179
transform 1 0 2576 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_22
timestamp 1649977179
transform 1 0 3128 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_47
timestamp 1649977179
transform 1 0 5428 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_61
timestamp 1649977179
transform 1 0 6716 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_67
timestamp 1649977179
transform 1 0 7268 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_71
timestamp 1649977179
transform 1 0 7636 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1649977179
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_95
timestamp 1649977179
transform 1 0 9844 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_102
timestamp 1649977179
transform 1 0 10488 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_106
timestamp 1649977179
transform 1 0 10856 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_123
timestamp 1649977179
transform 1 0 12420 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_132
timestamp 1649977179
transform 1 0 13248 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_157
timestamp 1649977179
transform 1 0 15548 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_165
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_173
timestamp 1649977179
transform 1 0 17020 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_181
timestamp 1649977179
transform 1 0 17756 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_192
timestamp 1649977179
transform 1 0 18768 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_207
timestamp 1649977179
transform 1 0 20148 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_211
timestamp 1649977179
transform 1 0 20516 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_217
timestamp 1649977179
transform 1 0 21068 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_229
timestamp 1649977179
transform 1 0 22172 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_243
timestamp 1649977179
transform 1 0 23460 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1649977179
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1649977179
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_271
timestamp 1649977179
transform 1 0 26036 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_283
timestamp 1649977179
transform 1 0 27140 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_290
timestamp 1649977179
transform 1 0 27784 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_294
timestamp 1649977179
transform 1 0 28152 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_297
timestamp 1649977179
transform 1 0 28428 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1649977179
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_314
timestamp 1649977179
transform 1 0 29992 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_320
timestamp 1649977179
transform 1 0 30544 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_340
timestamp 1649977179
transform 1 0 32384 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_30_358
timestamp 1649977179
transform 1 0 34040 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_30_365
timestamp 1649977179
transform 1 0 34684 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_370
timestamp 1649977179
transform 1 0 35144 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_376
timestamp 1649977179
transform 1 0 35696 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_379
timestamp 1649977179
transform 1 0 35972 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_403
timestamp 1649977179
transform 1 0 38180 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_415
timestamp 1649977179
transform 1 0 39284 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1649977179
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_423
timestamp 1649977179
transform 1 0 40020 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_435
timestamp 1649977179
transform 1 0 41124 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_447
timestamp 1649977179
transform 1 0 42228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_459
timestamp 1649977179
transform 1 0 43332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_471
timestamp 1649977179
transform 1 0 44436 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1649977179
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1649977179
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1649977179
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1649977179
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1649977179
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1649977179
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1649977179
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1649977179
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1649977179
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_557
timestamp 1649977179
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_569
timestamp 1649977179
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1649977179
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1649977179
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_589
timestamp 1649977179
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_601
timestamp 1649977179
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_613
timestamp 1649977179
transform 1 0 57500 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_625
timestamp 1649977179
transform 1 0 58604 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_637
timestamp 1649977179
transform 1 0 59708 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_643
timestamp 1649977179
transform 1 0 60260 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_645
timestamp 1649977179
transform 1 0 60444 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_657
timestamp 1649977179
transform 1 0 61548 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_669
timestamp 1649977179
transform 1 0 62652 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_681
timestamp 1649977179
transform 1 0 63756 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_693
timestamp 1649977179
transform 1 0 64860 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_699
timestamp 1649977179
transform 1 0 65412 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_701
timestamp 1649977179
transform 1 0 65596 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_713
timestamp 1649977179
transform 1 0 66700 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_725
timestamp 1649977179
transform 1 0 67804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_729
timestamp 1649977179
transform 1 0 68172 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_7
timestamp 1649977179
transform 1 0 1748 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_19
timestamp 1649977179
transform 1 0 2852 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_41
timestamp 1649977179
transform 1 0 4876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1649977179
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_60
timestamp 1649977179
transform 1 0 6624 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_74
timestamp 1649977179
transform 1 0 7912 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_88
timestamp 1649977179
transform 1 0 9200 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_94
timestamp 1649977179
transform 1 0 9752 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_100
timestamp 1649977179
transform 1 0 10304 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_126
timestamp 1649977179
transform 1 0 12696 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_132
timestamp 1649977179
transform 1 0 13248 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_144
timestamp 1649977179
transform 1 0 14352 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_151
timestamp 1649977179
transform 1 0 14996 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_163
timestamp 1649977179
transform 1 0 16100 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_171
timestamp 1649977179
transform 1 0 16836 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_177
timestamp 1649977179
transform 1 0 17388 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_189
timestamp 1649977179
transform 1 0 18492 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_193
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_201
timestamp 1649977179
transform 1 0 19596 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_214
timestamp 1649977179
transform 1 0 20792 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1649977179
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_225
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_231
timestamp 1649977179
transform 1 0 22356 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_245
timestamp 1649977179
transform 1 0 23644 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_249
timestamp 1649977179
transform 1 0 24012 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_260
timestamp 1649977179
transform 1 0 25024 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_272
timestamp 1649977179
transform 1 0 26128 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_275
timestamp 1649977179
transform 1 0 26404 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1649977179
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_297
timestamp 1649977179
transform 1 0 28428 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_303
timestamp 1649977179
transform 1 0 28980 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_320
timestamp 1649977179
transform 1 0 30544 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_326
timestamp 1649977179
transform 1 0 31096 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_331
timestamp 1649977179
transform 1 0 31556 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1649977179
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1649977179
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_349
timestamp 1649977179
transform 1 0 33212 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_366
timestamp 1649977179
transform 1 0 34776 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_378
timestamp 1649977179
transform 1 0 35880 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_384
timestamp 1649977179
transform 1 0 36432 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_393
timestamp 1649977179
transform 1 0 37260 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_404
timestamp 1649977179
transform 1 0 38272 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_412
timestamp 1649977179
transform 1 0 39008 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1649977179
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1649977179
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1649977179
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1649977179
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1649977179
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1649977179
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1649977179
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1649977179
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1649977179
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1649977179
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_517
timestamp 1649977179
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_529
timestamp 1649977179
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_541
timestamp 1649977179
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1649977179
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1649977179
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_561
timestamp 1649977179
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_573
timestamp 1649977179
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_585
timestamp 1649977179
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_597
timestamp 1649977179
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1649977179
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1649977179
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_617
timestamp 1649977179
transform 1 0 57868 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_629
timestamp 1649977179
transform 1 0 58972 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_641
timestamp 1649977179
transform 1 0 60076 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_653
timestamp 1649977179
transform 1 0 61180 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_665
timestamp 1649977179
transform 1 0 62284 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_671
timestamp 1649977179
transform 1 0 62836 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_673
timestamp 1649977179
transform 1 0 63020 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_685
timestamp 1649977179
transform 1 0 64124 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_697
timestamp 1649977179
transform 1 0 65228 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_709
timestamp 1649977179
transform 1 0 66332 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_721
timestamp 1649977179
transform 1 0 67436 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_727
timestamp 1649977179
transform 1 0 67988 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_729
timestamp 1649977179
transform 1 0 68172 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_7
timestamp 1649977179
transform 1 0 1748 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_16
timestamp 1649977179
transform 1 0 2576 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_22
timestamp 1649977179
transform 1 0 3128 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_43
timestamp 1649977179
transform 1 0 5060 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_63
timestamp 1649977179
transform 1 0 6900 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_71
timestamp 1649977179
transform 1 0 7636 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_80
timestamp 1649977179
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_104
timestamp 1649977179
transform 1 0 10672 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_112
timestamp 1649977179
transform 1 0 11408 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1649977179
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_158
timestamp 1649977179
transform 1 0 15640 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_166
timestamp 1649977179
transform 1 0 16376 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_170
timestamp 1649977179
transform 1 0 16744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_187
timestamp 1649977179
transform 1 0 18308 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1649977179
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_204
timestamp 1649977179
transform 1 0 19872 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_216
timestamp 1649977179
transform 1 0 20976 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_236
timestamp 1649977179
transform 1 0 22816 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_248
timestamp 1649977179
transform 1 0 23920 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_256
timestamp 1649977179
transform 1 0 24656 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_268
timestamp 1649977179
transform 1 0 25760 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_274
timestamp 1649977179
transform 1 0 26312 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_283
timestamp 1649977179
transform 1 0 27140 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_289
timestamp 1649977179
transform 1 0 27692 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_292
timestamp 1649977179
transform 1 0 27968 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_304
timestamp 1649977179
transform 1 0 29072 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_312
timestamp 1649977179
transform 1 0 29808 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_316
timestamp 1649977179
transform 1 0 30176 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_322
timestamp 1649977179
transform 1 0 30728 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_334
timestamp 1649977179
transform 1 0 31832 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_340
timestamp 1649977179
transform 1 0 32384 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_352
timestamp 1649977179
transform 1 0 33488 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_360
timestamp 1649977179
transform 1 0 34224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_370
timestamp 1649977179
transform 1 0 35144 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_374
timestamp 1649977179
transform 1 0 35512 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_391
timestamp 1649977179
transform 1 0 37076 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_400
timestamp 1649977179
transform 1 0 37904 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_412
timestamp 1649977179
transform 1 0 39008 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1649977179
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1649977179
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1649977179
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1649977179
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1649977179
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1649977179
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1649977179
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1649977179
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1649977179
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1649977179
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1649977179
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1649977179
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_533
timestamp 1649977179
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_545
timestamp 1649977179
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_557
timestamp 1649977179
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_569
timestamp 1649977179
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1649977179
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1649977179
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_589
timestamp 1649977179
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_601
timestamp 1649977179
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_613
timestamp 1649977179
transform 1 0 57500 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_625
timestamp 1649977179
transform 1 0 58604 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_637
timestamp 1649977179
transform 1 0 59708 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_643
timestamp 1649977179
transform 1 0 60260 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_645
timestamp 1649977179
transform 1 0 60444 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_657
timestamp 1649977179
transform 1 0 61548 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_669
timestamp 1649977179
transform 1 0 62652 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_681
timestamp 1649977179
transform 1 0 63756 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_693
timestamp 1649977179
transform 1 0 64860 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_699
timestamp 1649977179
transform 1 0 65412 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_701
timestamp 1649977179
transform 1 0 65596 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_713
timestamp 1649977179
transform 1 0 66700 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_725
timestamp 1649977179
transform 1 0 67804 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_729
timestamp 1649977179
transform 1 0 68172 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_12
timestamp 1649977179
transform 1 0 2208 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_34
timestamp 1649977179
transform 1 0 4232 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_43
timestamp 1649977179
transform 1 0 5060 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_49
timestamp 1649977179
transform 1 0 5612 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_52
timestamp 1649977179
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_59
timestamp 1649977179
transform 1 0 6532 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_68
timestamp 1649977179
transform 1 0 7360 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_80
timestamp 1649977179
transform 1 0 8464 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_86
timestamp 1649977179
transform 1 0 9016 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_92
timestamp 1649977179
transform 1 0 9568 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_108
timestamp 1649977179
transform 1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_118
timestamp 1649977179
transform 1 0 11960 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_122
timestamp 1649977179
transform 1 0 12328 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_139
timestamp 1649977179
transform 1 0 13892 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_151
timestamp 1649977179
transform 1 0 14996 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_155
timestamp 1649977179
transform 1 0 15364 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 1649977179
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_177
timestamp 1649977179
transform 1 0 17388 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_186
timestamp 1649977179
transform 1 0 18216 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_194
timestamp 1649977179
transform 1 0 18952 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_197
timestamp 1649977179
transform 1 0 19228 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_203
timestamp 1649977179
transform 1 0 19780 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_206
timestamp 1649977179
transform 1 0 20056 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_220
timestamp 1649977179
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_227
timestamp 1649977179
transform 1 0 21988 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_237
timestamp 1649977179
transform 1 0 22908 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_248
timestamp 1649977179
transform 1 0 23920 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_260
timestamp 1649977179
transform 1 0 25024 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_271
timestamp 1649977179
transform 1 0 26036 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1649977179
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_281
timestamp 1649977179
transform 1 0 26956 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_294
timestamp 1649977179
transform 1 0 28152 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_300
timestamp 1649977179
transform 1 0 28704 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_326
timestamp 1649977179
transform 1 0 31096 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_332
timestamp 1649977179
transform 1 0 31648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_353
timestamp 1649977179
transform 1 0 33580 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_362
timestamp 1649977179
transform 1 0 34408 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_368
timestamp 1649977179
transform 1 0 34960 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_377
timestamp 1649977179
transform 1 0 35788 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_383
timestamp 1649977179
transform 1 0 36340 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1649977179
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_393
timestamp 1649977179
transform 1 0 37260 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_396
timestamp 1649977179
transform 1 0 37536 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_402
timestamp 1649977179
transform 1 0 38088 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_419
timestamp 1649977179
transform 1 0 39652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_431
timestamp 1649977179
transform 1 0 40756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_443
timestamp 1649977179
transform 1 0 41860 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1649977179
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1649977179
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1649977179
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1649977179
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1649977179
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1649977179
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1649977179
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1649977179
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_517
timestamp 1649977179
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_529
timestamp 1649977179
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_541
timestamp 1649977179
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1649977179
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1649977179
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_561
timestamp 1649977179
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_573
timestamp 1649977179
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_585
timestamp 1649977179
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_597
timestamp 1649977179
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1649977179
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1649977179
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_617
timestamp 1649977179
transform 1 0 57868 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_629
timestamp 1649977179
transform 1 0 58972 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_641
timestamp 1649977179
transform 1 0 60076 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_653
timestamp 1649977179
transform 1 0 61180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_665
timestamp 1649977179
transform 1 0 62284 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_671
timestamp 1649977179
transform 1 0 62836 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_673
timestamp 1649977179
transform 1 0 63020 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_685
timestamp 1649977179
transform 1 0 64124 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_697
timestamp 1649977179
transform 1 0 65228 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_709
timestamp 1649977179
transform 1 0 66332 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_721
timestamp 1649977179
transform 1 0 67436 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_727
timestamp 1649977179
transform 1 0 67988 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_729
timestamp 1649977179
transform 1 0 68172 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_3
timestamp 1649977179
transform 1 0 1380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_17
timestamp 1649977179
transform 1 0 2668 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_21
timestamp 1649977179
transform 1 0 3036 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_24
timestamp 1649977179
transform 1 0 3312 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_32
timestamp 1649977179
transform 1 0 4048 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_56
timestamp 1649977179
transform 1 0 6256 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_76
timestamp 1649977179
transform 1 0 8096 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_85
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_88
timestamp 1649977179
transform 1 0 9200 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_100
timestamp 1649977179
transform 1 0 10304 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_108
timestamp 1649977179
transform 1 0 11040 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_111
timestamp 1649977179
transform 1 0 11316 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_123
timestamp 1649977179
transform 1 0 12420 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_135
timestamp 1649977179
transform 1 0 13524 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1649977179
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_157
timestamp 1649977179
transform 1 0 15548 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_165
timestamp 1649977179
transform 1 0 16284 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_169
timestamp 1649977179
transform 1 0 16652 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_175
timestamp 1649977179
transform 1 0 17204 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_181
timestamp 1649977179
transform 1 0 17756 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_192
timestamp 1649977179
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_205
timestamp 1649977179
transform 1 0 19964 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_211
timestamp 1649977179
transform 1 0 20516 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_218
timestamp 1649977179
transform 1 0 21160 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_226
timestamp 1649977179
transform 1 0 21896 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_232
timestamp 1649977179
transform 1 0 22448 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_236
timestamp 1649977179
transform 1 0 22816 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_247
timestamp 1649977179
transform 1 0 23828 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1649977179
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_255
timestamp 1649977179
transform 1 0 24564 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_267
timestamp 1649977179
transform 1 0 25668 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_295
timestamp 1649977179
transform 1 0 28244 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_304
timestamp 1649977179
transform 1 0 29072 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_309
timestamp 1649977179
transform 1 0 29532 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_313
timestamp 1649977179
transform 1 0 29900 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_319
timestamp 1649977179
transform 1 0 30452 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_325
timestamp 1649977179
transform 1 0 31004 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_333
timestamp 1649977179
transform 1 0 31740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_336
timestamp 1649977179
transform 1 0 32016 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_342
timestamp 1649977179
transform 1 0 32568 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_354
timestamp 1649977179
transform 1 0 33672 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_360
timestamp 1649977179
transform 1 0 34224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_365
timestamp 1649977179
transform 1 0 34684 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_376
timestamp 1649977179
transform 1 0 35696 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_382
timestamp 1649977179
transform 1 0 36248 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_402
timestamp 1649977179
transform 1 0 38088 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_414
timestamp 1649977179
transform 1 0 39192 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1649977179
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1649977179
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1649977179
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1649977179
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1649977179
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1649977179
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1649977179
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1649977179
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1649977179
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1649977179
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1649977179
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1649977179
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_533
timestamp 1649977179
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_545
timestamp 1649977179
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_557
timestamp 1649977179
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_569
timestamp 1649977179
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1649977179
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1649977179
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_589
timestamp 1649977179
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_601
timestamp 1649977179
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_613
timestamp 1649977179
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_625
timestamp 1649977179
transform 1 0 58604 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_637
timestamp 1649977179
transform 1 0 59708 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_643
timestamp 1649977179
transform 1 0 60260 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_645
timestamp 1649977179
transform 1 0 60444 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_657
timestamp 1649977179
transform 1 0 61548 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_669
timestamp 1649977179
transform 1 0 62652 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_681
timestamp 1649977179
transform 1 0 63756 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_693
timestamp 1649977179
transform 1 0 64860 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_699
timestamp 1649977179
transform 1 0 65412 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_701
timestamp 1649977179
transform 1 0 65596 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_713
timestamp 1649977179
transform 1 0 66700 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_725
timestamp 1649977179
transform 1 0 67804 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_35_3
timestamp 1649977179
transform 1 0 1380 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_11
timestamp 1649977179
transform 1 0 2116 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_23
timestamp 1649977179
transform 1 0 3220 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_31
timestamp 1649977179
transform 1 0 3956 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_35
timestamp 1649977179
transform 1 0 4324 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_52
timestamp 1649977179
transform 1 0 5888 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_60
timestamp 1649977179
transform 1 0 6624 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_66
timestamp 1649977179
transform 1 0 7176 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_70
timestamp 1649977179
transform 1 0 7544 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_87
timestamp 1649977179
transform 1 0 9108 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_91
timestamp 1649977179
transform 1 0 9476 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_108
timestamp 1649977179
transform 1 0 11040 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_113
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_119
timestamp 1649977179
transform 1 0 12052 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_139
timestamp 1649977179
transform 1 0 13892 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_151
timestamp 1649977179
transform 1 0 14996 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_159
timestamp 1649977179
transform 1 0 15732 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1649977179
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_173
timestamp 1649977179
transform 1 0 17020 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_35_185
timestamp 1649977179
transform 1 0 18124 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_207
timestamp 1649977179
transform 1 0 20148 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp 1649977179
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_235
timestamp 1649977179
transform 1 0 22724 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_248
timestamp 1649977179
transform 1 0 23920 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_254
timestamp 1649977179
transform 1 0 24472 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_260
timestamp 1649977179
transform 1 0 25024 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_269
timestamp 1649977179
transform 1 0 25852 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_273
timestamp 1649977179
transform 1 0 26220 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 1649977179
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_289
timestamp 1649977179
transform 1 0 27692 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_297
timestamp 1649977179
transform 1 0 28428 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_301
timestamp 1649977179
transform 1 0 28796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_315
timestamp 1649977179
transform 1 0 30084 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_327
timestamp 1649977179
transform 1 0 31188 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1649977179
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_337
timestamp 1649977179
transform 1 0 32108 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_345
timestamp 1649977179
transform 1 0 32844 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_351
timestamp 1649977179
transform 1 0 33396 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_368
timestamp 1649977179
transform 1 0 34960 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_388
timestamp 1649977179
transform 1 0 36800 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1649977179
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_405
timestamp 1649977179
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_417
timestamp 1649977179
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_429
timestamp 1649977179
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1649977179
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1649977179
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1649977179
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1649977179
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1649977179
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1649977179
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1649977179
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1649977179
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1649977179
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_517
timestamp 1649977179
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_529
timestamp 1649977179
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_541
timestamp 1649977179
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1649977179
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1649977179
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_561
timestamp 1649977179
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_573
timestamp 1649977179
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_585
timestamp 1649977179
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_597
timestamp 1649977179
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1649977179
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1649977179
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_617
timestamp 1649977179
transform 1 0 57868 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_629
timestamp 1649977179
transform 1 0 58972 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_641
timestamp 1649977179
transform 1 0 60076 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_653
timestamp 1649977179
transform 1 0 61180 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_665
timestamp 1649977179
transform 1 0 62284 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_671
timestamp 1649977179
transform 1 0 62836 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_673
timestamp 1649977179
transform 1 0 63020 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_685
timestamp 1649977179
transform 1 0 64124 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_697
timestamp 1649977179
transform 1 0 65228 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_709
timestamp 1649977179
transform 1 0 66332 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_724
timestamp 1649977179
transform 1 0 67712 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_729
timestamp 1649977179
transform 1 0 68172 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_3
timestamp 1649977179
transform 1 0 1380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_11
timestamp 1649977179
transform 1 0 2116 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_17
timestamp 1649977179
transform 1 0 2668 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_23
timestamp 1649977179
transform 1 0 3220 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1649977179
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_33
timestamp 1649977179
transform 1 0 4140 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_41
timestamp 1649977179
transform 1 0 4876 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_48
timestamp 1649977179
transform 1 0 5520 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_54
timestamp 1649977179
transform 1 0 6072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_68
timestamp 1649977179
transform 1 0 7360 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_74
timestamp 1649977179
transform 1 0 7912 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1649977179
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_90
timestamp 1649977179
transform 1 0 9384 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_94
timestamp 1649977179
transform 1 0 9752 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_100
timestamp 1649977179
transform 1 0 10304 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_112
timestamp 1649977179
transform 1 0 11408 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_124
timestamp 1649977179
transform 1 0 12512 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_136
timestamp 1649977179
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_141
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_146
timestamp 1649977179
transform 1 0 14536 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_157
timestamp 1649977179
transform 1 0 15548 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_173
timestamp 1649977179
transform 1 0 17020 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_179
timestamp 1649977179
transform 1 0 17572 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_192
timestamp 1649977179
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_199
timestamp 1649977179
transform 1 0 19412 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_213
timestamp 1649977179
transform 1 0 20700 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_227
timestamp 1649977179
transform 1 0 21988 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_236
timestamp 1649977179
transform 1 0 22816 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_243
timestamp 1649977179
transform 1 0 23460 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1649977179
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_253
timestamp 1649977179
transform 1 0 24380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_261
timestamp 1649977179
transform 1 0 25116 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_269
timestamp 1649977179
transform 1 0 25852 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_283
timestamp 1649977179
transform 1 0 27140 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1649977179
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1649977179
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1649977179
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_309
timestamp 1649977179
transform 1 0 29532 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_313
timestamp 1649977179
transform 1 0 29900 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_319
timestamp 1649977179
transform 1 0 30452 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_323
timestamp 1649977179
transform 1 0 30820 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_340
timestamp 1649977179
transform 1 0 32384 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_360
timestamp 1649977179
transform 1 0 34224 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1649977179
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_379
timestamp 1649977179
transform 1 0 35972 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_403
timestamp 1649977179
transform 1 0 38180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_415
timestamp 1649977179
transform 1 0 39284 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1649977179
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1649977179
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1649977179
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1649977179
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1649977179
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1649977179
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1649977179
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1649977179
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1649977179
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1649977179
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_513
timestamp 1649977179
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1649977179
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1649977179
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_533
timestamp 1649977179
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_545
timestamp 1649977179
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_557
timestamp 1649977179
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_569
timestamp 1649977179
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1649977179
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1649977179
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_589
timestamp 1649977179
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_601
timestamp 1649977179
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_613
timestamp 1649977179
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_625
timestamp 1649977179
transform 1 0 58604 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_637
timestamp 1649977179
transform 1 0 59708 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_643
timestamp 1649977179
transform 1 0 60260 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_645
timestamp 1649977179
transform 1 0 60444 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_657
timestamp 1649977179
transform 1 0 61548 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_669
timestamp 1649977179
transform 1 0 62652 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_681
timestamp 1649977179
transform 1 0 63756 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_693
timestamp 1649977179
transform 1 0 64860 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_699
timestamp 1649977179
transform 1 0 65412 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_701
timestamp 1649977179
transform 1 0 65596 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_713
timestamp 1649977179
transform 1 0 66700 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_725
timestamp 1649977179
transform 1 0 67804 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_3
timestamp 1649977179
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_15
timestamp 1649977179
transform 1 0 2484 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_35
timestamp 1649977179
transform 1 0 4324 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_47
timestamp 1649977179
transform 1 0 5428 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1649977179
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_57
timestamp 1649977179
transform 1 0 6348 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_61
timestamp 1649977179
transform 1 0 6716 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_70
timestamp 1649977179
transform 1 0 7544 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_79
timestamp 1649977179
transform 1 0 8372 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_83
timestamp 1649977179
transform 1 0 8740 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_92
timestamp 1649977179
transform 1 0 9568 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_98
timestamp 1649977179
transform 1 0 10120 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1649977179
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1649977179
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_125
timestamp 1649977179
transform 1 0 12604 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_133
timestamp 1649977179
transform 1 0 13340 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_143
timestamp 1649977179
transform 1 0 14260 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_155
timestamp 1649977179
transform 1 0 15364 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_163
timestamp 1649977179
transform 1 0 16100 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1649977179
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_185
timestamp 1649977179
transform 1 0 18124 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_189
timestamp 1649977179
transform 1 0 18492 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_198
timestamp 1649977179
transform 1 0 19320 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_206
timestamp 1649977179
transform 1 0 20056 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1649977179
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1649977179
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_235
timestamp 1649977179
transform 1 0 22724 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_239
timestamp 1649977179
transform 1 0 23092 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_256
timestamp 1649977179
transform 1 0 24656 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_262
timestamp 1649977179
transform 1 0 25208 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_267
timestamp 1649977179
transform 1 0 25668 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_275
timestamp 1649977179
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1649977179
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_281
timestamp 1649977179
transform 1 0 26956 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_285
timestamp 1649977179
transform 1 0 27324 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_294
timestamp 1649977179
transform 1 0 28152 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_302
timestamp 1649977179
transform 1 0 28888 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_308
timestamp 1649977179
transform 1 0 29440 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_324
timestamp 1649977179
transform 1 0 30912 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_332
timestamp 1649977179
transform 1 0 31648 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_339
timestamp 1649977179
transform 1 0 32292 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_351
timestamp 1649977179
transform 1 0 33396 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_363
timestamp 1649977179
transform 1 0 34500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_375
timestamp 1649977179
transform 1 0 35604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_387
timestamp 1649977179
transform 1 0 36708 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1649977179
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1649977179
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_405
timestamp 1649977179
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_417
timestamp 1649977179
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_429
timestamp 1649977179
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1649977179
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1649977179
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1649977179
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1649977179
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1649977179
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1649977179
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1649977179
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1649977179
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1649977179
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_517
timestamp 1649977179
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_529
timestamp 1649977179
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_541
timestamp 1649977179
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1649977179
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1649977179
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_561
timestamp 1649977179
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_573
timestamp 1649977179
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_585
timestamp 1649977179
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_597
timestamp 1649977179
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1649977179
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1649977179
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_617
timestamp 1649977179
transform 1 0 57868 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_629
timestamp 1649977179
transform 1 0 58972 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_641
timestamp 1649977179
transform 1 0 60076 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_653
timestamp 1649977179
transform 1 0 61180 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_665
timestamp 1649977179
transform 1 0 62284 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_671
timestamp 1649977179
transform 1 0 62836 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_673
timestamp 1649977179
transform 1 0 63020 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_685
timestamp 1649977179
transform 1 0 64124 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_697
timestamp 1649977179
transform 1 0 65228 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_709
timestamp 1649977179
transform 1 0 66332 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_724
timestamp 1649977179
transform 1 0 67712 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_729
timestamp 1649977179
transform 1 0 68172 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1649977179
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_9
timestamp 1649977179
transform 1 0 1932 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_21
timestamp 1649977179
transform 1 0 3036 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1649977179
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_45
timestamp 1649977179
transform 1 0 5244 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_53
timestamp 1649977179
transform 1 0 5980 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_62
timestamp 1649977179
transform 1 0 6808 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_71
timestamp 1649977179
transform 1 0 7636 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_80
timestamp 1649977179
transform 1 0 8464 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_90
timestamp 1649977179
transform 1 0 9384 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_110
timestamp 1649977179
transform 1 0 11224 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_130
timestamp 1649977179
transform 1 0 13064 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1649977179
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1649977179
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_148
timestamp 1649977179
transform 1 0 14720 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_159
timestamp 1649977179
transform 1 0 15732 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_163
timestamp 1649977179
transform 1 0 16100 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_166
timestamp 1649977179
transform 1 0 16376 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_180
timestamp 1649977179
transform 1 0 17664 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_188
timestamp 1649977179
transform 1 0 18400 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_192
timestamp 1649977179
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1649977179
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_207
timestamp 1649977179
transform 1 0 20148 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_227
timestamp 1649977179
transform 1 0 21988 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_233
timestamp 1649977179
transform 1 0 22540 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_242
timestamp 1649977179
transform 1 0 23368 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_248
timestamp 1649977179
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1649977179
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_265
timestamp 1649977179
transform 1 0 25484 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_282
timestamp 1649977179
transform 1 0 27048 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_304
timestamp 1649977179
transform 1 0 29072 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_319
timestamp 1649977179
transform 1 0 30452 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_326
timestamp 1649977179
transform 1 0 31096 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_330
timestamp 1649977179
transform 1 0 31464 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_347
timestamp 1649977179
transform 1 0 33028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_359
timestamp 1649977179
transform 1 0 34132 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1649977179
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1649977179
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1649977179
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1649977179
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_401
timestamp 1649977179
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1649977179
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1649977179
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1649977179
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1649977179
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1649977179
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1649977179
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1649977179
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1649977179
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1649977179
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1649977179
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1649977179
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_513
timestamp 1649977179
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1649977179
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1649977179
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_533
timestamp 1649977179
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_545
timestamp 1649977179
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_557
timestamp 1649977179
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_569
timestamp 1649977179
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1649977179
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1649977179
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_589
timestamp 1649977179
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_601
timestamp 1649977179
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_613
timestamp 1649977179
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_625
timestamp 1649977179
transform 1 0 58604 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_637
timestamp 1649977179
transform 1 0 59708 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_643
timestamp 1649977179
transform 1 0 60260 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_645
timestamp 1649977179
transform 1 0 60444 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_657
timestamp 1649977179
transform 1 0 61548 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_669
timestamp 1649977179
transform 1 0 62652 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_681
timestamp 1649977179
transform 1 0 63756 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_693
timestamp 1649977179
transform 1 0 64860 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_699
timestamp 1649977179
transform 1 0 65412 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_701
timestamp 1649977179
transform 1 0 65596 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_713
timestamp 1649977179
transform 1 0 66700 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_725
timestamp 1649977179
transform 1 0 67804 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1649977179
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_17
timestamp 1649977179
transform 1 0 2668 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_29
timestamp 1649977179
transform 1 0 3772 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_35
timestamp 1649977179
transform 1 0 4324 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_43
timestamp 1649977179
transform 1 0 5060 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_52
timestamp 1649977179
transform 1 0 5888 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_59
timestamp 1649977179
transform 1 0 6532 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_73
timestamp 1649977179
transform 1 0 7820 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_85
timestamp 1649977179
transform 1 0 8924 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_91
timestamp 1649977179
transform 1 0 9476 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_103
timestamp 1649977179
transform 1 0 10580 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1649977179
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_113
timestamp 1649977179
transform 1 0 11500 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_121
timestamp 1649977179
transform 1 0 12236 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_128
timestamp 1649977179
transform 1 0 12880 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_140
timestamp 1649977179
transform 1 0 13984 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_148
timestamp 1649977179
transform 1 0 14720 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_157
timestamp 1649977179
transform 1 0 15548 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_163
timestamp 1649977179
transform 1 0 16100 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1649977179
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_169
timestamp 1649977179
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_173
timestamp 1649977179
transform 1 0 17020 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_182
timestamp 1649977179
transform 1 0 17848 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_190
timestamp 1649977179
transform 1 0 18584 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_193
timestamp 1649977179
transform 1 0 18860 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_202
timestamp 1649977179
transform 1 0 19688 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_214
timestamp 1649977179
transform 1 0 20792 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 1649977179
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1649977179
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_231
timestamp 1649977179
transform 1 0 22356 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_245
timestamp 1649977179
transform 1 0 23644 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_259
timestamp 1649977179
transform 1 0 24932 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1649977179
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1649977179
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_286
timestamp 1649977179
transform 1 0 27416 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_292
timestamp 1649977179
transform 1 0 27968 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_314
timestamp 1649977179
transform 1 0 29992 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_320
timestamp 1649977179
transform 1 0 30544 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1649977179
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1649977179
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1649977179
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1649977179
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1649977179
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1649977179
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1649977179
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1649977179
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1649977179
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_405
timestamp 1649977179
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_417
timestamp 1649977179
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_429
timestamp 1649977179
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1649977179
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1649977179
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1649977179
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1649977179
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1649977179
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1649977179
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1649977179
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1649977179
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_505
timestamp 1649977179
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_517
timestamp 1649977179
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_529
timestamp 1649977179
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_541
timestamp 1649977179
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1649977179
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1649977179
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_561
timestamp 1649977179
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_573
timestamp 1649977179
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_585
timestamp 1649977179
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_597
timestamp 1649977179
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1649977179
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1649977179
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_617
timestamp 1649977179
transform 1 0 57868 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_629
timestamp 1649977179
transform 1 0 58972 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_641
timestamp 1649977179
transform 1 0 60076 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_653
timestamp 1649977179
transform 1 0 61180 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_665
timestamp 1649977179
transform 1 0 62284 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_671
timestamp 1649977179
transform 1 0 62836 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_673
timestamp 1649977179
transform 1 0 63020 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_685
timestamp 1649977179
transform 1 0 64124 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_697
timestamp 1649977179
transform 1 0 65228 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_709
timestamp 1649977179
transform 1 0 66332 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_721
timestamp 1649977179
transform 1 0 67436 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_727
timestamp 1649977179
transform 1 0 67988 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_729
timestamp 1649977179
transform 1 0 68172 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1649977179
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_10
timestamp 1649977179
transform 1 0 2024 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_24
timestamp 1649977179
transform 1 0 3312 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_31
timestamp 1649977179
transform 1 0 3956 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_37
timestamp 1649977179
transform 1 0 4508 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_51
timestamp 1649977179
transform 1 0 5796 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_59
timestamp 1649977179
transform 1 0 6532 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_63
timestamp 1649977179
transform 1 0 6900 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_72
timestamp 1649977179
transform 1 0 7728 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_79
timestamp 1649977179
transform 1 0 8372 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1649977179
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_85
timestamp 1649977179
transform 1 0 8924 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_89
timestamp 1649977179
transform 1 0 9292 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_106
timestamp 1649977179
transform 1 0 10856 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_118
timestamp 1649977179
transform 1 0 11960 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_127
timestamp 1649977179
transform 1 0 12788 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_133
timestamp 1649977179
transform 1 0 13340 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_136
timestamp 1649977179
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_141
timestamp 1649977179
transform 1 0 14076 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_146
timestamp 1649977179
transform 1 0 14536 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_160
timestamp 1649977179
transform 1 0 15824 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_168
timestamp 1649977179
transform 1 0 16560 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_177
timestamp 1649977179
transform 1 0 17388 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_183
timestamp 1649977179
transform 1 0 17940 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1649977179
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1649977179
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_205
timestamp 1649977179
transform 1 0 19964 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_209
timestamp 1649977179
transform 1 0 20332 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_212
timestamp 1649977179
transform 1 0 20608 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_220
timestamp 1649977179
transform 1 0 21344 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_230
timestamp 1649977179
transform 1 0 22264 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_237
timestamp 1649977179
transform 1 0 22908 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_241
timestamp 1649977179
transform 1 0 23276 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_247
timestamp 1649977179
transform 1 0 23828 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1649977179
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_253
timestamp 1649977179
transform 1 0 24380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_258
timestamp 1649977179
transform 1 0 24840 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_264
timestamp 1649977179
transform 1 0 25392 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_285
timestamp 1649977179
transform 1 0 27324 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_297
timestamp 1649977179
transform 1 0 28428 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_305
timestamp 1649977179
transform 1 0 29164 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_309
timestamp 1649977179
transform 1 0 29532 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_317
timestamp 1649977179
transform 1 0 30268 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_322
timestamp 1649977179
transform 1 0 30728 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_334
timestamp 1649977179
transform 1 0 31832 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_40_358
timestamp 1649977179
transform 1 0 34040 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1649977179
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1649977179
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1649977179
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1649977179
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1649977179
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1649977179
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1649977179
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1649977179
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_445
timestamp 1649977179
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_457
timestamp 1649977179
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1649977179
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1649977179
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1649977179
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1649977179
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1649977179
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_513
timestamp 1649977179
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1649977179
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1649977179
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_533
timestamp 1649977179
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_545
timestamp 1649977179
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_557
timestamp 1649977179
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_569
timestamp 1649977179
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1649977179
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1649977179
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_589
timestamp 1649977179
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_601
timestamp 1649977179
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_613
timestamp 1649977179
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_625
timestamp 1649977179
transform 1 0 58604 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_637
timestamp 1649977179
transform 1 0 59708 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_643
timestamp 1649977179
transform 1 0 60260 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_645
timestamp 1649977179
transform 1 0 60444 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_657
timestamp 1649977179
transform 1 0 61548 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_669
timestamp 1649977179
transform 1 0 62652 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_681
timestamp 1649977179
transform 1 0 63756 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_693
timestamp 1649977179
transform 1 0 64860 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_699
timestamp 1649977179
transform 1 0 65412 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_701
timestamp 1649977179
transform 1 0 65596 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_713
timestamp 1649977179
transform 1 0 66700 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_725
timestamp 1649977179
transform 1 0 67804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_729
timestamp 1649977179
transform 1 0 68172 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_8
timestamp 1649977179
transform 1 0 1840 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_20
timestamp 1649977179
transform 1 0 2944 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_28
timestamp 1649977179
transform 1 0 3680 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_45
timestamp 1649977179
transform 1 0 5244 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_53
timestamp 1649977179
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_57
timestamp 1649977179
transform 1 0 6348 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_61
timestamp 1649977179
transform 1 0 6716 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_72
timestamp 1649977179
transform 1 0 7728 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_88
timestamp 1649977179
transform 1 0 9200 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_108
timestamp 1649977179
transform 1 0 11040 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_113
timestamp 1649977179
transform 1 0 11500 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_126
timestamp 1649977179
transform 1 0 12696 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_140
timestamp 1649977179
transform 1 0 13984 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_164
timestamp 1649977179
transform 1 0 16192 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1649977179
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_181
timestamp 1649977179
transform 1 0 17756 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_186
timestamp 1649977179
transform 1 0 18216 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_206
timestamp 1649977179
transform 1 0 20056 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_212
timestamp 1649977179
transform 1 0 20608 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_227
timestamp 1649977179
transform 1 0 21988 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_239
timestamp 1649977179
transform 1 0 23092 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_251
timestamp 1649977179
transform 1 0 24196 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_257
timestamp 1649977179
transform 1 0 24748 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_262
timestamp 1649977179
transform 1 0 25208 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_274
timestamp 1649977179
transform 1 0 26312 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_297
timestamp 1649977179
transform 1 0 28428 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_309
timestamp 1649977179
transform 1 0 29532 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_318
timestamp 1649977179
transform 1 0 30360 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_327
timestamp 1649977179
transform 1 0 31188 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1649977179
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1649977179
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1649977179
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1649977179
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1649977179
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1649977179
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1649977179
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1649977179
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_405
timestamp 1649977179
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_417
timestamp 1649977179
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_429
timestamp 1649977179
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1649977179
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1649977179
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1649977179
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1649977179
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1649977179
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1649977179
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1649977179
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1649977179
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1649977179
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1649977179
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1649977179
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1649977179
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1649977179
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1649977179
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1649977179
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_573
timestamp 1649977179
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_585
timestamp 1649977179
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_597
timestamp 1649977179
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1649977179
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1649977179
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_617
timestamp 1649977179
transform 1 0 57868 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_629
timestamp 1649977179
transform 1 0 58972 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_641
timestamp 1649977179
transform 1 0 60076 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_653
timestamp 1649977179
transform 1 0 61180 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_665
timestamp 1649977179
transform 1 0 62284 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_671
timestamp 1649977179
transform 1 0 62836 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_673
timestamp 1649977179
transform 1 0 63020 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_685
timestamp 1649977179
transform 1 0 64124 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_697
timestamp 1649977179
transform 1 0 65228 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_709
timestamp 1649977179
transform 1 0 66332 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_721
timestamp 1649977179
transform 1 0 67436 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_727
timestamp 1649977179
transform 1 0 67988 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_729
timestamp 1649977179
transform 1 0 68172 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_3
timestamp 1649977179
transform 1 0 1380 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_9
timestamp 1649977179
transform 1 0 1932 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_21
timestamp 1649977179
transform 1 0 3036 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1649977179
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_31
timestamp 1649977179
transform 1 0 3956 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_43
timestamp 1649977179
transform 1 0 5060 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_62
timestamp 1649977179
transform 1 0 6808 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_68
timestamp 1649977179
transform 1 0 7360 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_80
timestamp 1649977179
transform 1 0 8464 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_90
timestamp 1649977179
transform 1 0 9384 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_96
timestamp 1649977179
transform 1 0 9936 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_108
timestamp 1649977179
transform 1 0 11040 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_120
timestamp 1649977179
transform 1 0 12144 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_136
timestamp 1649977179
transform 1 0 13616 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_151
timestamp 1649977179
transform 1 0 14996 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_159
timestamp 1649977179
transform 1 0 15732 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_163
timestamp 1649977179
transform 1 0 16100 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_171
timestamp 1649977179
transform 1 0 16836 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_181
timestamp 1649977179
transform 1 0 17756 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 1649977179
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_42_197
timestamp 1649977179
transform 1 0 19228 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_208
timestamp 1649977179
transform 1 0 20240 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_228
timestamp 1649977179
transform 1 0 22080 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_248
timestamp 1649977179
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_253
timestamp 1649977179
transform 1 0 24380 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_261
timestamp 1649977179
transform 1 0 25116 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_269
timestamp 1649977179
transform 1 0 25852 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_275
timestamp 1649977179
transform 1 0 26404 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_286
timestamp 1649977179
transform 1 0 27416 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_298
timestamp 1649977179
transform 1 0 28520 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_306
timestamp 1649977179
transform 1 0 29256 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_309
timestamp 1649977179
transform 1 0 29532 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_314
timestamp 1649977179
transform 1 0 29992 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_320
timestamp 1649977179
transform 1 0 30544 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_332
timestamp 1649977179
transform 1 0 31648 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_352
timestamp 1649977179
transform 1 0 33488 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1649977179
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1649977179
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1649977179
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1649977179
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1649977179
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1649977179
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1649977179
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1649977179
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1649977179
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1649977179
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1649977179
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1649977179
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1649977179
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1649977179
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1649977179
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_513
timestamp 1649977179
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1649977179
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1649977179
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1649977179
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1649977179
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_557
timestamp 1649977179
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_569
timestamp 1649977179
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1649977179
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1649977179
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_589
timestamp 1649977179
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_601
timestamp 1649977179
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_613
timestamp 1649977179
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_625
timestamp 1649977179
transform 1 0 58604 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_637
timestamp 1649977179
transform 1 0 59708 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_643
timestamp 1649977179
transform 1 0 60260 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_645
timestamp 1649977179
transform 1 0 60444 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_657
timestamp 1649977179
transform 1 0 61548 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_669
timestamp 1649977179
transform 1 0 62652 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_681
timestamp 1649977179
transform 1 0 63756 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_693
timestamp 1649977179
transform 1 0 64860 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_699
timestamp 1649977179
transform 1 0 65412 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_701
timestamp 1649977179
transform 1 0 65596 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_713
timestamp 1649977179
transform 1 0 66700 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_725
timestamp 1649977179
transform 1 0 67804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_729
timestamp 1649977179
transform 1 0 68172 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_3
timestamp 1649977179
transform 1 0 1380 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_7
timestamp 1649977179
transform 1 0 1748 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_13
timestamp 1649977179
transform 1 0 2300 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_35
timestamp 1649977179
transform 1 0 4324 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_47
timestamp 1649977179
transform 1 0 5428 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1649977179
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_57
timestamp 1649977179
transform 1 0 6348 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_81
timestamp 1649977179
transform 1 0 8556 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_101
timestamp 1649977179
transform 1 0 10396 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_109
timestamp 1649977179
transform 1 0 11132 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_113
timestamp 1649977179
transform 1 0 11500 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_132
timestamp 1649977179
transform 1 0 13248 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_138
timestamp 1649977179
transform 1 0 13800 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_146
timestamp 1649977179
transform 1 0 14536 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_150
timestamp 1649977179
transform 1 0 14904 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1649977179
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_179
timestamp 1649977179
transform 1 0 17572 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_187
timestamp 1649977179
transform 1 0 18308 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_196
timestamp 1649977179
transform 1 0 19136 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_220
timestamp 1649977179
transform 1 0 21344 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_233
timestamp 1649977179
transform 1 0 22540 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_239
timestamp 1649977179
transform 1 0 23092 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_247
timestamp 1649977179
transform 1 0 23828 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_259
timestamp 1649977179
transform 1 0 24932 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_271
timestamp 1649977179
transform 1 0 26036 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_276
timestamp 1649977179
transform 1 0 26496 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_281
timestamp 1649977179
transform 1 0 26956 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_290
timestamp 1649977179
transform 1 0 27784 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_310
timestamp 1649977179
transform 1 0 29624 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_314
timestamp 1649977179
transform 1 0 29992 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_323
timestamp 1649977179
transform 1 0 30820 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_332
timestamp 1649977179
transform 1 0 31648 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1649977179
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1649977179
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1649977179
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1649977179
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1649977179
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1649977179
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1649977179
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1649977179
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_417
timestamp 1649977179
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1649977179
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1649977179
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1649977179
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1649977179
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1649977179
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1649977179
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1649977179
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1649977179
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1649977179
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1649977179
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1649977179
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1649977179
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1649977179
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1649977179
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1649977179
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_561
timestamp 1649977179
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_573
timestamp 1649977179
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_585
timestamp 1649977179
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_597
timestamp 1649977179
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1649977179
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1649977179
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_617
timestamp 1649977179
transform 1 0 57868 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_629
timestamp 1649977179
transform 1 0 58972 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_641
timestamp 1649977179
transform 1 0 60076 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_653
timestamp 1649977179
transform 1 0 61180 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_665
timestamp 1649977179
transform 1 0 62284 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_671
timestamp 1649977179
transform 1 0 62836 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_673
timestamp 1649977179
transform 1 0 63020 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_685
timestamp 1649977179
transform 1 0 64124 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_697
timestamp 1649977179
transform 1 0 65228 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_709
timestamp 1649977179
transform 1 0 66332 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_721
timestamp 1649977179
transform 1 0 67436 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_727
timestamp 1649977179
transform 1 0 67988 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_729
timestamp 1649977179
transform 1 0 68172 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_3
timestamp 1649977179
transform 1 0 1380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_9
timestamp 1649977179
transform 1 0 1932 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_20
timestamp 1649977179
transform 1 0 2944 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_31
timestamp 1649977179
transform 1 0 3956 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_35
timestamp 1649977179
transform 1 0 4324 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_52
timestamp 1649977179
transform 1 0 5888 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_68
timestamp 1649977179
transform 1 0 7360 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1649977179
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1649977179
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_87
timestamp 1649977179
transform 1 0 9108 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_99
timestamp 1649977179
transform 1 0 10212 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_117
timestamp 1649977179
transform 1 0 11868 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_129
timestamp 1649977179
transform 1 0 12972 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_137
timestamp 1649977179
transform 1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_148
timestamp 1649977179
transform 1 0 14720 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_152
timestamp 1649977179
transform 1 0 15088 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_161
timestamp 1649977179
transform 1 0 15916 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_169
timestamp 1649977179
transform 1 0 16652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_178
timestamp 1649977179
transform 1 0 17480 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_192
timestamp 1649977179
transform 1 0 18768 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_200
timestamp 1649977179
transform 1 0 19504 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_204
timestamp 1649977179
transform 1 0 19872 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_215
timestamp 1649977179
transform 1 0 20884 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_219
timestamp 1649977179
transform 1 0 21252 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_236
timestamp 1649977179
transform 1 0 22816 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_242
timestamp 1649977179
transform 1 0 23368 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 1649977179
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_253
timestamp 1649977179
transform 1 0 24380 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_272
timestamp 1649977179
transform 1 0 26128 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_281
timestamp 1649977179
transform 1 0 26956 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_293
timestamp 1649977179
transform 1 0 28060 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_305
timestamp 1649977179
transform 1 0 29164 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_309
timestamp 1649977179
transform 1 0 29532 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_317
timestamp 1649977179
transform 1 0 30268 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_334
timestamp 1649977179
transform 1 0 31832 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_346
timestamp 1649977179
transform 1 0 32936 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_358
timestamp 1649977179
transform 1 0 34040 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1649977179
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1649977179
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1649977179
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_401
timestamp 1649977179
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1649977179
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1649977179
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1649977179
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1649977179
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1649977179
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1649977179
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1649977179
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1649977179
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1649977179
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1649977179
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1649977179
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_513
timestamp 1649977179
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1649977179
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1649977179
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_533
timestamp 1649977179
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_545
timestamp 1649977179
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_557
timestamp 1649977179
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_569
timestamp 1649977179
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1649977179
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1649977179
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_589
timestamp 1649977179
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_601
timestamp 1649977179
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_613
timestamp 1649977179
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_625
timestamp 1649977179
transform 1 0 58604 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_637
timestamp 1649977179
transform 1 0 59708 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_643
timestamp 1649977179
transform 1 0 60260 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_645
timestamp 1649977179
transform 1 0 60444 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_657
timestamp 1649977179
transform 1 0 61548 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_669
timestamp 1649977179
transform 1 0 62652 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_681
timestamp 1649977179
transform 1 0 63756 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_693
timestamp 1649977179
transform 1 0 64860 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_699
timestamp 1649977179
transform 1 0 65412 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_701
timestamp 1649977179
transform 1 0 65596 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_713
timestamp 1649977179
transform 1 0 66700 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_725
timestamp 1649977179
transform 1 0 67804 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_45_3
timestamp 1649977179
transform 1 0 1380 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_14
timestamp 1649977179
transform 1 0 2392 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_28
timestamp 1649977179
transform 1 0 3680 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_48
timestamp 1649977179
transform 1 0 5520 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_45_57
timestamp 1649977179
transform 1 0 6348 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_66
timestamp 1649977179
transform 1 0 7176 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_86
timestamp 1649977179
transform 1 0 9016 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_95
timestamp 1649977179
transform 1 0 9844 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_107
timestamp 1649977179
transform 1 0 10948 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1649977179
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_113
timestamp 1649977179
transform 1 0 11500 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_121
timestamp 1649977179
transform 1 0 12236 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_128
timestamp 1649977179
transform 1 0 12880 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_139
timestamp 1649977179
transform 1 0 13892 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_152
timestamp 1649977179
transform 1 0 15088 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_164
timestamp 1649977179
transform 1 0 16192 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_174
timestamp 1649977179
transform 1 0 17112 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_181
timestamp 1649977179
transform 1 0 17756 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_190
timestamp 1649977179
transform 1 0 18584 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_202
timestamp 1649977179
transform 1 0 19688 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_206
timestamp 1649977179
transform 1 0 20056 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_212
timestamp 1649977179
transform 1 0 20608 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_219
timestamp 1649977179
transform 1 0 21252 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1649977179
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1649977179
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_237
timestamp 1649977179
transform 1 0 22908 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_244
timestamp 1649977179
transform 1 0 23552 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1649977179
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_273
timestamp 1649977179
transform 1 0 26220 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_276
timestamp 1649977179
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_289
timestamp 1649977179
transform 1 0 27692 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_298
timestamp 1649977179
transform 1 0 28520 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_310
timestamp 1649977179
transform 1 0 29624 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_322
timestamp 1649977179
transform 1 0 30728 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_334
timestamp 1649977179
transform 1 0 31832 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1649977179
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1649977179
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1649977179
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1649977179
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1649977179
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1649977179
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1649977179
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1649977179
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1649977179
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1649977179
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1649977179
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1649977179
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1649977179
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1649977179
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1649977179
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1649977179
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1649977179
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1649977179
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1649977179
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_517
timestamp 1649977179
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_529
timestamp 1649977179
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_541
timestamp 1649977179
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1649977179
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1649977179
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_561
timestamp 1649977179
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_573
timestamp 1649977179
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_585
timestamp 1649977179
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_597
timestamp 1649977179
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1649977179
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1649977179
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_617
timestamp 1649977179
transform 1 0 57868 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_629
timestamp 1649977179
transform 1 0 58972 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_641
timestamp 1649977179
transform 1 0 60076 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_653
timestamp 1649977179
transform 1 0 61180 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_665
timestamp 1649977179
transform 1 0 62284 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_671
timestamp 1649977179
transform 1 0 62836 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_673
timestamp 1649977179
transform 1 0 63020 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_685
timestamp 1649977179
transform 1 0 64124 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_697
timestamp 1649977179
transform 1 0 65228 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_709
timestamp 1649977179
transform 1 0 66332 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_724
timestamp 1649977179
transform 1 0 67712 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_729
timestamp 1649977179
transform 1 0 68172 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_3
timestamp 1649977179
transform 1 0 1380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_9
timestamp 1649977179
transform 1 0 1932 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_13
timestamp 1649977179
transform 1 0 2300 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_24
timestamp 1649977179
transform 1 0 3312 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_37
timestamp 1649977179
transform 1 0 4508 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_45
timestamp 1649977179
transform 1 0 5244 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_63
timestamp 1649977179
transform 1 0 6900 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_75
timestamp 1649977179
transform 1 0 8004 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1649977179
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_85
timestamp 1649977179
transform 1 0 8924 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_98
timestamp 1649977179
transform 1 0 10120 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_106
timestamp 1649977179
transform 1 0 10856 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_124
timestamp 1649977179
transform 1 0 12512 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_130
timestamp 1649977179
transform 1 0 13064 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_136
timestamp 1649977179
transform 1 0 13616 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_149
timestamp 1649977179
transform 1 0 14812 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_155
timestamp 1649977179
transform 1 0 15364 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_166
timestamp 1649977179
transform 1 0 16376 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_178
timestamp 1649977179
transform 1 0 17480 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_184
timestamp 1649977179
transform 1 0 18032 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1649977179
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_200
timestamp 1649977179
transform 1 0 19504 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_206
timestamp 1649977179
transform 1 0 20056 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_217
timestamp 1649977179
transform 1 0 21068 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_223
timestamp 1649977179
transform 1 0 21620 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_227
timestamp 1649977179
transform 1 0 21988 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_233
timestamp 1649977179
transform 1 0 22540 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_239
timestamp 1649977179
transform 1 0 23092 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_248
timestamp 1649977179
transform 1 0 23920 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_253
timestamp 1649977179
transform 1 0 24380 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_256
timestamp 1649977179
transform 1 0 24656 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_268
timestamp 1649977179
transform 1 0 25760 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_277
timestamp 1649977179
transform 1 0 26588 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_281
timestamp 1649977179
transform 1 0 26956 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_284
timestamp 1649977179
transform 1 0 27232 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_296
timestamp 1649977179
transform 1 0 28336 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1649977179
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1649977179
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1649977179
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1649977179
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1649977179
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1649977179
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1649977179
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1649977179
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1649977179
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_401
timestamp 1649977179
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1649977179
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1649977179
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1649977179
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1649977179
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1649977179
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1649977179
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1649977179
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1649977179
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1649977179
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1649977179
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1649977179
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_513
timestamp 1649977179
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1649977179
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1649977179
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_533
timestamp 1649977179
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_545
timestamp 1649977179
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_557
timestamp 1649977179
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_569
timestamp 1649977179
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1649977179
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1649977179
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_589
timestamp 1649977179
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_601
timestamp 1649977179
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_613
timestamp 1649977179
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_625
timestamp 1649977179
transform 1 0 58604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_637
timestamp 1649977179
transform 1 0 59708 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_643
timestamp 1649977179
transform 1 0 60260 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_645
timestamp 1649977179
transform 1 0 60444 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_657
timestamp 1649977179
transform 1 0 61548 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_669
timestamp 1649977179
transform 1 0 62652 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_681
timestamp 1649977179
transform 1 0 63756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_693
timestamp 1649977179
transform 1 0 64860 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_699
timestamp 1649977179
transform 1 0 65412 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_701
timestamp 1649977179
transform 1 0 65596 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_713
timestamp 1649977179
transform 1 0 66700 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_725
timestamp 1649977179
transform 1 0 67804 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_3
timestamp 1649977179
transform 1 0 1380 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_7
timestamp 1649977179
transform 1 0 1748 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_16
timestamp 1649977179
transform 1 0 2576 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_22
timestamp 1649977179
transform 1 0 3128 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_34
timestamp 1649977179
transform 1 0 4232 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_46
timestamp 1649977179
transform 1 0 5336 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_54
timestamp 1649977179
transform 1 0 6072 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_57
timestamp 1649977179
transform 1 0 6348 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_67
timestamp 1649977179
transform 1 0 7268 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_73
timestamp 1649977179
transform 1 0 7820 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_85
timestamp 1649977179
transform 1 0 8924 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_99
timestamp 1649977179
transform 1 0 10212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1649977179
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_113
timestamp 1649977179
transform 1 0 11500 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_121
timestamp 1649977179
transform 1 0 12236 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_131
timestamp 1649977179
transform 1 0 13156 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_137
timestamp 1649977179
transform 1 0 13708 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_157
timestamp 1649977179
transform 1 0 15548 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_163
timestamp 1649977179
transform 1 0 16100 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1649977179
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_171
timestamp 1649977179
transform 1 0 16836 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_191
timestamp 1649977179
transform 1 0 18676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_202
timestamp 1649977179
transform 1 0 19688 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_214
timestamp 1649977179
transform 1 0 20792 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_220
timestamp 1649977179
transform 1 0 21344 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1649977179
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_235
timestamp 1649977179
transform 1 0 22724 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_241
timestamp 1649977179
transform 1 0 23276 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_253
timestamp 1649977179
transform 1 0 24380 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_269
timestamp 1649977179
transform 1 0 25852 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_275
timestamp 1649977179
transform 1 0 26404 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1649977179
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1649977179
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1649977179
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_305
timestamp 1649977179
transform 1 0 29164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_322
timestamp 1649977179
transform 1 0 30728 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_334
timestamp 1649977179
transform 1 0 31832 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1649977179
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1649977179
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1649977179
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1649977179
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1649977179
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1649977179
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1649977179
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1649977179
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1649977179
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1649977179
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1649977179
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1649977179
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1649977179
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1649977179
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1649977179
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1649977179
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1649977179
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1649977179
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1649977179
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_517
timestamp 1649977179
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_529
timestamp 1649977179
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1649977179
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1649977179
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1649977179
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_561
timestamp 1649977179
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_573
timestamp 1649977179
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_585
timestamp 1649977179
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_597
timestamp 1649977179
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1649977179
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1649977179
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_617
timestamp 1649977179
transform 1 0 57868 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_629
timestamp 1649977179
transform 1 0 58972 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_641
timestamp 1649977179
transform 1 0 60076 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_653
timestamp 1649977179
transform 1 0 61180 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_665
timestamp 1649977179
transform 1 0 62284 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_671
timestamp 1649977179
transform 1 0 62836 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_673
timestamp 1649977179
transform 1 0 63020 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_685
timestamp 1649977179
transform 1 0 64124 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_697
timestamp 1649977179
transform 1 0 65228 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_709
timestamp 1649977179
transform 1 0 66332 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_724
timestamp 1649977179
transform 1 0 67712 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_729
timestamp 1649977179
transform 1 0 68172 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_48_3
timestamp 1649977179
transform 1 0 1380 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_11
timestamp 1649977179
transform 1 0 2116 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_19
timestamp 1649977179
transform 1 0 2852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_24
timestamp 1649977179
transform 1 0 3312 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_37
timestamp 1649977179
transform 1 0 4508 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_49
timestamp 1649977179
transform 1 0 5612 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_55
timestamp 1649977179
transform 1 0 6164 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_58
timestamp 1649977179
transform 1 0 6440 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_62
timestamp 1649977179
transform 1 0 6808 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_65
timestamp 1649977179
transform 1 0 7084 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1649977179
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1649977179
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_85
timestamp 1649977179
transform 1 0 8924 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_89
timestamp 1649977179
transform 1 0 9292 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_92
timestamp 1649977179
transform 1 0 9568 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_112
timestamp 1649977179
transform 1 0 11408 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_124
timestamp 1649977179
transform 1 0 12512 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_128
timestamp 1649977179
transform 1 0 12880 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_136
timestamp 1649977179
transform 1 0 13616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_141
timestamp 1649977179
transform 1 0 14076 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_165
timestamp 1649977179
transform 1 0 16284 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_169
timestamp 1649977179
transform 1 0 16652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_178
timestamp 1649977179
transform 1 0 17480 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_184
timestamp 1649977179
transform 1 0 18032 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_197
timestamp 1649977179
transform 1 0 19228 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_205
timestamp 1649977179
transform 1 0 19964 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_222
timestamp 1649977179
transform 1 0 21528 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_226
timestamp 1649977179
transform 1 0 21896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_243
timestamp 1649977179
transform 1 0 23460 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1649977179
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1649977179
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_265
timestamp 1649977179
transform 1 0 25484 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_284
timestamp 1649977179
transform 1 0 27232 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_304
timestamp 1649977179
transform 1 0 29072 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1649977179
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1649977179
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1649977179
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1649977179
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1649977179
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1649977179
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1649977179
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1649977179
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1649977179
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_401
timestamp 1649977179
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1649977179
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1649977179
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1649977179
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1649977179
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1649977179
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1649977179
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1649977179
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1649977179
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1649977179
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1649977179
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1649977179
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_513
timestamp 1649977179
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1649977179
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1649977179
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_533
timestamp 1649977179
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_545
timestamp 1649977179
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_557
timestamp 1649977179
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_569
timestamp 1649977179
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1649977179
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1649977179
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_589
timestamp 1649977179
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_601
timestamp 1649977179
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_613
timestamp 1649977179
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_625
timestamp 1649977179
transform 1 0 58604 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_637
timestamp 1649977179
transform 1 0 59708 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_643
timestamp 1649977179
transform 1 0 60260 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_645
timestamp 1649977179
transform 1 0 60444 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_657
timestamp 1649977179
transform 1 0 61548 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_669
timestamp 1649977179
transform 1 0 62652 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_681
timestamp 1649977179
transform 1 0 63756 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_693
timestamp 1649977179
transform 1 0 64860 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_699
timestamp 1649977179
transform 1 0 65412 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_701
timestamp 1649977179
transform 1 0 65596 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_713
timestamp 1649977179
transform 1 0 66700 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_725
timestamp 1649977179
transform 1 0 67804 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_49_3
timestamp 1649977179
transform 1 0 1380 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_11
timestamp 1649977179
transform 1 0 2116 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_22
timestamp 1649977179
transform 1 0 3128 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_28
timestamp 1649977179
transform 1 0 3680 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_48
timestamp 1649977179
transform 1 0 5520 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_57
timestamp 1649977179
transform 1 0 6348 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_66
timestamp 1649977179
transform 1 0 7176 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_88
timestamp 1649977179
transform 1 0 9200 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_100
timestamp 1649977179
transform 1 0 10304 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_129
timestamp 1649977179
transform 1 0 12972 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_141
timestamp 1649977179
transform 1 0 14076 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_145
timestamp 1649977179
transform 1 0 14444 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_156
timestamp 1649977179
transform 1 0 15456 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_164
timestamp 1649977179
transform 1 0 16192 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1649977179
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_178
timestamp 1649977179
transform 1 0 17480 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_184
timestamp 1649977179
transform 1 0 18032 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_190
timestamp 1649977179
transform 1 0 18584 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_202
timestamp 1649977179
transform 1 0 19688 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_214
timestamp 1649977179
transform 1 0 20792 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 1649977179
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1649977179
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_237
timestamp 1649977179
transform 1 0 22908 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_245
timestamp 1649977179
transform 1 0 23644 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_262
timestamp 1649977179
transform 1 0 25208 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_274
timestamp 1649977179
transform 1 0 26312 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_281
timestamp 1649977179
transform 1 0 26956 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_305
timestamp 1649977179
transform 1 0 29164 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_311
timestamp 1649977179
transform 1 0 29716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_323
timestamp 1649977179
transform 1 0 30820 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1649977179
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1649977179
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1649977179
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1649977179
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1649977179
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1649977179
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1649977179
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1649977179
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1649977179
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1649977179
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1649977179
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1649977179
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1649977179
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1649977179
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1649977179
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1649977179
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1649977179
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1649977179
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1649977179
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1649977179
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_517
timestamp 1649977179
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_529
timestamp 1649977179
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1649977179
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1649977179
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1649977179
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_561
timestamp 1649977179
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_573
timestamp 1649977179
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_585
timestamp 1649977179
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_597
timestamp 1649977179
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1649977179
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1649977179
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_617
timestamp 1649977179
transform 1 0 57868 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_629
timestamp 1649977179
transform 1 0 58972 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_641
timestamp 1649977179
transform 1 0 60076 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_653
timestamp 1649977179
transform 1 0 61180 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_665
timestamp 1649977179
transform 1 0 62284 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_671
timestamp 1649977179
transform 1 0 62836 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_673
timestamp 1649977179
transform 1 0 63020 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_685
timestamp 1649977179
transform 1 0 64124 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_697
timestamp 1649977179
transform 1 0 65228 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_709
timestamp 1649977179
transform 1 0 66332 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_721
timestamp 1649977179
transform 1 0 67436 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_727
timestamp 1649977179
transform 1 0 67988 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_729
timestamp 1649977179
transform 1 0 68172 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_5
timestamp 1649977179
transform 1 0 1564 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_17
timestamp 1649977179
transform 1 0 2668 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_25
timestamp 1649977179
transform 1 0 3404 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_34
timestamp 1649977179
transform 1 0 4232 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_46
timestamp 1649977179
transform 1 0 5336 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_50_56
timestamp 1649977179
transform 1 0 6256 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_64
timestamp 1649977179
transform 1 0 6992 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_70
timestamp 1649977179
transform 1 0 7544 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_79
timestamp 1649977179
transform 1 0 8372 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1649977179
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_85
timestamp 1649977179
transform 1 0 8924 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_91
timestamp 1649977179
transform 1 0 9476 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_108
timestamp 1649977179
transform 1 0 11040 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_116
timestamp 1649977179
transform 1 0 11776 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_124
timestamp 1649977179
transform 1 0 12512 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_136
timestamp 1649977179
transform 1 0 13616 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_143
timestamp 1649977179
transform 1 0 14260 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_155
timestamp 1649977179
transform 1 0 15364 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_169
timestamp 1649977179
transform 1 0 16652 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_180
timestamp 1649977179
transform 1 0 17664 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_192
timestamp 1649977179
transform 1 0 18768 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_205
timestamp 1649977179
transform 1 0 19964 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_211
timestamp 1649977179
transform 1 0 20516 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_223
timestamp 1649977179
transform 1 0 21620 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_234
timestamp 1649977179
transform 1 0 22632 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_246
timestamp 1649977179
transform 1 0 23736 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1649977179
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_265
timestamp 1649977179
transform 1 0 25484 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_282
timestamp 1649977179
transform 1 0 27048 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_294
timestamp 1649977179
transform 1 0 28152 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_306
timestamp 1649977179
transform 1 0 29256 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1649977179
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1649977179
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1649977179
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1649977179
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1649977179
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1649977179
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1649977179
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1649977179
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1649977179
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1649977179
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1649977179
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1649977179
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1649977179
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1649977179
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1649977179
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1649977179
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1649977179
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1649977179
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1649977179
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1649977179
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1649977179
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_513
timestamp 1649977179
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1649977179
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1649977179
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_533
timestamp 1649977179
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_545
timestamp 1649977179
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_557
timestamp 1649977179
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_569
timestamp 1649977179
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1649977179
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1649977179
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_589
timestamp 1649977179
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_601
timestamp 1649977179
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_613
timestamp 1649977179
transform 1 0 57500 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_625
timestamp 1649977179
transform 1 0 58604 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_637
timestamp 1649977179
transform 1 0 59708 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_643
timestamp 1649977179
transform 1 0 60260 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_645
timestamp 1649977179
transform 1 0 60444 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_657
timestamp 1649977179
transform 1 0 61548 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_669
timestamp 1649977179
transform 1 0 62652 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_681
timestamp 1649977179
transform 1 0 63756 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_693
timestamp 1649977179
transform 1 0 64860 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_699
timestamp 1649977179
transform 1 0 65412 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_701
timestamp 1649977179
transform 1 0 65596 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_713
timestamp 1649977179
transform 1 0 66700 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_725
timestamp 1649977179
transform 1 0 67804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_729
timestamp 1649977179
transform 1 0 68172 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_3
timestamp 1649977179
transform 1 0 1380 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_10
timestamp 1649977179
transform 1 0 2024 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_19
timestamp 1649977179
transform 1 0 2852 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_31
timestamp 1649977179
transform 1 0 3956 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_35
timestamp 1649977179
transform 1 0 4324 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_52
timestamp 1649977179
transform 1 0 5888 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1649977179
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_69
timestamp 1649977179
transform 1 0 7452 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_90
timestamp 1649977179
transform 1 0 9384 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_96
timestamp 1649977179
transform 1 0 9936 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_108
timestamp 1649977179
transform 1 0 11040 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1649977179
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_125
timestamp 1649977179
transform 1 0 12604 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_139
timestamp 1649977179
transform 1 0 13892 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_145
timestamp 1649977179
transform 1 0 14444 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_151
timestamp 1649977179
transform 1 0 14996 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_162
timestamp 1649977179
transform 1 0 16008 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1649977179
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1649977179
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_193
timestamp 1649977179
transform 1 0 18860 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_199
timestamp 1649977179
transform 1 0 19412 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_216
timestamp 1649977179
transform 1 0 20976 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_230
timestamp 1649977179
transform 1 0 22264 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_250
timestamp 1649977179
transform 1 0 24104 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_270
timestamp 1649977179
transform 1 0 25944 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_278
timestamp 1649977179
transform 1 0 26680 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1649977179
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1649977179
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1649977179
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1649977179
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1649977179
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1649977179
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1649977179
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1649977179
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1649977179
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1649977179
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1649977179
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1649977179
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1649977179
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1649977179
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1649977179
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1649977179
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1649977179
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1649977179
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1649977179
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1649977179
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1649977179
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1649977179
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1649977179
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1649977179
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1649977179
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_517
timestamp 1649977179
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_529
timestamp 1649977179
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1649977179
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1649977179
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1649977179
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_561
timestamp 1649977179
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_573
timestamp 1649977179
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_585
timestamp 1649977179
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_597
timestamp 1649977179
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1649977179
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1649977179
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_617
timestamp 1649977179
transform 1 0 57868 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_629
timestamp 1649977179
transform 1 0 58972 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_641
timestamp 1649977179
transform 1 0 60076 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_653
timestamp 1649977179
transform 1 0 61180 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_665
timestamp 1649977179
transform 1 0 62284 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_671
timestamp 1649977179
transform 1 0 62836 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_673
timestamp 1649977179
transform 1 0 63020 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_685
timestamp 1649977179
transform 1 0 64124 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_697
timestamp 1649977179
transform 1 0 65228 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_709
timestamp 1649977179
transform 1 0 66332 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_721
timestamp 1649977179
transform 1 0 67436 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_727
timestamp 1649977179
transform 1 0 67988 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_729
timestamp 1649977179
transform 1 0 68172 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1649977179
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1649977179
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1649977179
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1649977179
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1649977179
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_53
timestamp 1649977179
transform 1 0 5980 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1649977179
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1649977179
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_85
timestamp 1649977179
transform 1 0 8924 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_96
timestamp 1649977179
transform 1 0 9936 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_108
timestamp 1649977179
transform 1 0 11040 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_128
timestamp 1649977179
transform 1 0 12880 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_157
timestamp 1649977179
transform 1 0 15548 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_165
timestamp 1649977179
transform 1 0 16284 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_182
timestamp 1649977179
transform 1 0 17848 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1649977179
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_202
timestamp 1649977179
transform 1 0 19688 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_214
timestamp 1649977179
transform 1 0 20792 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_236
timestamp 1649977179
transform 1 0 22816 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_248
timestamp 1649977179
transform 1 0 23920 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1649977179
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1649977179
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1649977179
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1649977179
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1649977179
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1649977179
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1649977179
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1649977179
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1649977179
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1649977179
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1649977179
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1649977179
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1649977179
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1649977179
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1649977179
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_401
timestamp 1649977179
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1649977179
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1649977179
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1649977179
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1649977179
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1649977179
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1649977179
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1649977179
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1649977179
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1649977179
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1649977179
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1649977179
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1649977179
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1649977179
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1649977179
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_533
timestamp 1649977179
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_545
timestamp 1649977179
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_557
timestamp 1649977179
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_569
timestamp 1649977179
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1649977179
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1649977179
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_589
timestamp 1649977179
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_601
timestamp 1649977179
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_613
timestamp 1649977179
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_625
timestamp 1649977179
transform 1 0 58604 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_637
timestamp 1649977179
transform 1 0 59708 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_643
timestamp 1649977179
transform 1 0 60260 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_645
timestamp 1649977179
transform 1 0 60444 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_657
timestamp 1649977179
transform 1 0 61548 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_669
timestamp 1649977179
transform 1 0 62652 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_681
timestamp 1649977179
transform 1 0 63756 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_693
timestamp 1649977179
transform 1 0 64860 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_699
timestamp 1649977179
transform 1 0 65412 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_701
timestamp 1649977179
transform 1 0 65596 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_713
timestamp 1649977179
transform 1 0 66700 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_725
timestamp 1649977179
transform 1 0 67804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_729
timestamp 1649977179
transform 1 0 68172 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1649977179
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_15
timestamp 1649977179
transform 1 0 2484 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_35
timestamp 1649977179
transform 1 0 4324 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_47
timestamp 1649977179
transform 1 0 5428 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1649977179
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1649977179
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1649977179
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1649977179
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1649977179
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1649977179
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1649977179
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1649977179
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_125
timestamp 1649977179
transform 1 0 12604 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_132
timestamp 1649977179
transform 1 0 13248 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_144
timestamp 1649977179
transform 1 0 14352 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_53_160
timestamp 1649977179
transform 1 0 15824 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_53_171
timestamp 1649977179
transform 1 0 16836 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_182
timestamp 1649977179
transform 1 0 17848 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_194
timestamp 1649977179
transform 1 0 18952 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_206
timestamp 1649977179
transform 1 0 20056 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_218
timestamp 1649977179
transform 1 0 21160 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1649977179
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_237
timestamp 1649977179
transform 1 0 22908 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_251
timestamp 1649977179
transform 1 0 24196 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_257
timestamp 1649977179
transform 1 0 24748 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_269
timestamp 1649977179
transform 1 0 25852 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_277
timestamp 1649977179
transform 1 0 26588 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1649977179
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1649977179
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1649977179
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1649977179
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1649977179
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1649977179
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1649977179
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1649977179
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1649977179
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1649977179
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1649977179
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1649977179
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1649977179
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1649977179
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1649977179
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1649977179
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1649977179
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1649977179
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1649977179
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1649977179
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1649977179
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1649977179
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1649977179
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1649977179
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1649977179
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_517
timestamp 1649977179
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_529
timestamp 1649977179
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1649977179
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1649977179
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1649977179
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_561
timestamp 1649977179
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_573
timestamp 1649977179
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_585
timestamp 1649977179
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_597
timestamp 1649977179
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1649977179
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1649977179
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_617
timestamp 1649977179
transform 1 0 57868 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_629
timestamp 1649977179
transform 1 0 58972 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_641
timestamp 1649977179
transform 1 0 60076 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_653
timestamp 1649977179
transform 1 0 61180 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_665
timestamp 1649977179
transform 1 0 62284 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_671
timestamp 1649977179
transform 1 0 62836 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_673
timestamp 1649977179
transform 1 0 63020 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_685
timestamp 1649977179
transform 1 0 64124 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_697
timestamp 1649977179
transform 1 0 65228 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_709
timestamp 1649977179
transform 1 0 66332 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_721
timestamp 1649977179
transform 1 0 67436 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_727
timestamp 1649977179
transform 1 0 67988 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_729
timestamp 1649977179
transform 1 0 68172 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1649977179
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1649977179
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1649977179
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1649977179
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1649977179
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1649977179
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1649977179
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1649977179
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1649977179
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1649977179
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1649977179
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1649977179
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1649977179
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1649977179
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1649977179
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_141
timestamp 1649977179
transform 1 0 14076 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_149
timestamp 1649977179
transform 1 0 14812 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_157
timestamp 1649977179
transform 1 0 15548 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_169
timestamp 1649977179
transform 1 0 16652 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_181
timestamp 1649977179
transform 1 0 17756 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_193
timestamp 1649977179
transform 1 0 18860 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_199
timestamp 1649977179
transform 1 0 19412 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_216
timestamp 1649977179
transform 1 0 20976 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_228
timestamp 1649977179
transform 1 0 22080 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_234
timestamp 1649977179
transform 1 0 22632 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_238
timestamp 1649977179
transform 1 0 23000 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_244
timestamp 1649977179
transform 1 0 23552 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1649977179
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1649977179
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1649977179
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1649977179
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1649977179
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1649977179
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1649977179
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1649977179
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1649977179
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1649977179
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1649977179
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1649977179
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1649977179
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1649977179
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1649977179
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_401
timestamp 1649977179
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1649977179
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1649977179
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1649977179
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1649977179
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1649977179
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1649977179
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1649977179
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1649977179
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1649977179
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1649977179
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1649977179
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_513
timestamp 1649977179
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1649977179
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1649977179
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_533
timestamp 1649977179
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_545
timestamp 1649977179
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_557
timestamp 1649977179
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_569
timestamp 1649977179
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1649977179
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1649977179
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_589
timestamp 1649977179
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_601
timestamp 1649977179
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_613
timestamp 1649977179
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_625
timestamp 1649977179
transform 1 0 58604 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_637
timestamp 1649977179
transform 1 0 59708 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_643
timestamp 1649977179
transform 1 0 60260 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_645
timestamp 1649977179
transform 1 0 60444 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_657
timestamp 1649977179
transform 1 0 61548 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_669
timestamp 1649977179
transform 1 0 62652 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_681
timestamp 1649977179
transform 1 0 63756 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_693
timestamp 1649977179
transform 1 0 64860 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_699
timestamp 1649977179
transform 1 0 65412 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_701
timestamp 1649977179
transform 1 0 65596 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_713
timestamp 1649977179
transform 1 0 66700 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_725
timestamp 1649977179
transform 1 0 67804 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1649977179
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1649977179
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1649977179
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1649977179
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1649977179
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1649977179
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1649977179
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1649977179
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1649977179
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1649977179
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1649977179
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1649977179
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1649977179
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1649977179
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1649977179
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1649977179
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1649977179
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1649977179
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1649977179
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1649977179
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1649977179
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1649977179
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1649977179
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1649977179
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1649977179
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1649977179
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1649977179
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1649977179
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1649977179
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1649977179
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1649977179
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1649977179
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1649977179
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1649977179
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1649977179
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1649977179
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1649977179
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1649977179
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1649977179
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1649977179
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1649977179
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1649977179
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1649977179
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1649977179
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1649977179
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1649977179
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1649977179
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1649977179
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1649977179
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1649977179
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1649977179
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1649977179
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1649977179
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1649977179
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1649977179
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1649977179
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1649977179
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1649977179
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1649977179
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1649977179
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_561
timestamp 1649977179
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_573
timestamp 1649977179
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_585
timestamp 1649977179
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_597
timestamp 1649977179
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1649977179
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1649977179
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_617
timestamp 1649977179
transform 1 0 57868 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_629
timestamp 1649977179
transform 1 0 58972 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_641
timestamp 1649977179
transform 1 0 60076 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_653
timestamp 1649977179
transform 1 0 61180 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_665
timestamp 1649977179
transform 1 0 62284 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_671
timestamp 1649977179
transform 1 0 62836 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_673
timestamp 1649977179
transform 1 0 63020 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_685
timestamp 1649977179
transform 1 0 64124 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_697
timestamp 1649977179
transform 1 0 65228 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_709
timestamp 1649977179
transform 1 0 66332 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_724
timestamp 1649977179
transform 1 0 67712 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_729
timestamp 1649977179
transform 1 0 68172 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1649977179
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1649977179
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1649977179
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1649977179
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1649977179
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1649977179
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1649977179
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1649977179
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1649977179
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1649977179
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1649977179
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1649977179
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1649977179
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1649977179
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1649977179
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1649977179
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1649977179
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1649977179
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1649977179
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1649977179
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1649977179
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1649977179
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1649977179
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1649977179
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1649977179
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1649977179
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1649977179
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1649977179
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1649977179
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1649977179
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1649977179
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1649977179
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1649977179
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1649977179
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1649977179
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1649977179
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1649977179
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1649977179
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1649977179
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1649977179
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1649977179
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1649977179
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1649977179
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1649977179
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1649977179
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1649977179
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1649977179
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1649977179
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1649977179
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1649977179
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1649977179
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1649977179
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1649977179
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1649977179
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_513
timestamp 1649977179
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1649977179
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1649977179
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_533
timestamp 1649977179
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_545
timestamp 1649977179
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_557
timestamp 1649977179
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_569
timestamp 1649977179
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1649977179
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1649977179
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_589
timestamp 1649977179
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_601
timestamp 1649977179
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_613
timestamp 1649977179
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_625
timestamp 1649977179
transform 1 0 58604 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_637
timestamp 1649977179
transform 1 0 59708 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_643
timestamp 1649977179
transform 1 0 60260 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_645
timestamp 1649977179
transform 1 0 60444 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_657
timestamp 1649977179
transform 1 0 61548 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_669
timestamp 1649977179
transform 1 0 62652 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_681
timestamp 1649977179
transform 1 0 63756 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_693
timestamp 1649977179
transform 1 0 64860 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_699
timestamp 1649977179
transform 1 0 65412 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_701
timestamp 1649977179
transform 1 0 65596 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_713
timestamp 1649977179
transform 1 0 66700 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_725
timestamp 1649977179
transform 1 0 67804 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1649977179
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1649977179
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1649977179
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1649977179
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1649977179
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1649977179
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1649977179
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1649977179
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1649977179
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1649977179
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1649977179
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1649977179
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1649977179
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1649977179
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1649977179
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1649977179
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1649977179
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1649977179
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1649977179
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1649977179
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1649977179
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1649977179
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1649977179
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1649977179
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1649977179
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1649977179
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1649977179
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1649977179
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1649977179
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1649977179
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1649977179
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1649977179
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1649977179
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1649977179
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1649977179
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1649977179
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1649977179
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1649977179
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1649977179
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1649977179
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1649977179
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1649977179
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1649977179
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1649977179
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1649977179
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1649977179
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1649977179
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1649977179
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1649977179
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1649977179
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1649977179
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1649977179
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1649977179
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1649977179
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1649977179
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_517
timestamp 1649977179
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_529
timestamp 1649977179
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1649977179
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1649977179
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1649977179
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_561
timestamp 1649977179
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_573
timestamp 1649977179
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_585
timestamp 1649977179
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_597
timestamp 1649977179
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1649977179
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1649977179
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_617
timestamp 1649977179
transform 1 0 57868 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_629
timestamp 1649977179
transform 1 0 58972 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_641
timestamp 1649977179
transform 1 0 60076 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_653
timestamp 1649977179
transform 1 0 61180 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_665
timestamp 1649977179
transform 1 0 62284 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_671
timestamp 1649977179
transform 1 0 62836 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_673
timestamp 1649977179
transform 1 0 63020 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_685
timestamp 1649977179
transform 1 0 64124 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_697
timestamp 1649977179
transform 1 0 65228 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_709
timestamp 1649977179
transform 1 0 66332 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_724
timestamp 1649977179
transform 1 0 67712 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_729
timestamp 1649977179
transform 1 0 68172 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1649977179
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1649977179
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1649977179
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1649977179
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1649977179
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1649977179
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1649977179
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1649977179
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1649977179
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1649977179
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1649977179
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1649977179
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1649977179
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1649977179
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1649977179
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1649977179
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1649977179
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1649977179
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1649977179
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1649977179
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1649977179
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1649977179
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1649977179
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1649977179
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1649977179
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1649977179
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1649977179
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1649977179
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1649977179
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1649977179
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1649977179
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1649977179
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1649977179
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1649977179
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1649977179
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1649977179
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1649977179
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1649977179
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1649977179
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1649977179
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1649977179
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1649977179
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_401
timestamp 1649977179
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1649977179
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1649977179
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1649977179
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1649977179
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1649977179
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1649977179
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1649977179
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1649977179
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1649977179
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1649977179
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1649977179
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1649977179
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1649977179
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1649977179
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_533
timestamp 1649977179
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_545
timestamp 1649977179
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_557
timestamp 1649977179
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_569
timestamp 1649977179
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1649977179
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1649977179
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_589
timestamp 1649977179
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_601
timestamp 1649977179
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_613
timestamp 1649977179
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_625
timestamp 1649977179
transform 1 0 58604 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_637
timestamp 1649977179
transform 1 0 59708 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_643
timestamp 1649977179
transform 1 0 60260 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_645
timestamp 1649977179
transform 1 0 60444 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_657
timestamp 1649977179
transform 1 0 61548 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_669
timestamp 1649977179
transform 1 0 62652 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_681
timestamp 1649977179
transform 1 0 63756 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_693
timestamp 1649977179
transform 1 0 64860 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_699
timestamp 1649977179
transform 1 0 65412 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_701
timestamp 1649977179
transform 1 0 65596 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_713
timestamp 1649977179
transform 1 0 66700 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_725
timestamp 1649977179
transform 1 0 67804 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1649977179
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1649977179
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1649977179
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1649977179
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1649977179
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1649977179
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1649977179
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1649977179
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1649977179
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1649977179
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1649977179
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1649977179
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1649977179
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1649977179
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1649977179
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1649977179
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1649977179
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1649977179
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1649977179
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1649977179
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1649977179
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1649977179
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1649977179
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1649977179
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1649977179
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1649977179
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1649977179
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1649977179
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1649977179
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1649977179
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1649977179
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1649977179
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1649977179
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1649977179
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1649977179
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1649977179
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1649977179
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1649977179
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1649977179
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1649977179
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1649977179
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1649977179
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1649977179
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1649977179
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1649977179
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1649977179
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1649977179
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1649977179
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1649977179
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1649977179
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1649977179
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1649977179
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1649977179
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1649977179
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1649977179
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_517
timestamp 1649977179
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_529
timestamp 1649977179
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_541
timestamp 1649977179
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1649977179
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1649977179
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_561
timestamp 1649977179
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_573
timestamp 1649977179
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_585
timestamp 1649977179
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_597
timestamp 1649977179
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1649977179
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1649977179
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_617
timestamp 1649977179
transform 1 0 57868 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_629
timestamp 1649977179
transform 1 0 58972 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_641
timestamp 1649977179
transform 1 0 60076 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_653
timestamp 1649977179
transform 1 0 61180 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_665
timestamp 1649977179
transform 1 0 62284 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_671
timestamp 1649977179
transform 1 0 62836 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_673
timestamp 1649977179
transform 1 0 63020 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_685
timestamp 1649977179
transform 1 0 64124 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_697
timestamp 1649977179
transform 1 0 65228 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_709
timestamp 1649977179
transform 1 0 66332 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_721
timestamp 1649977179
transform 1 0 67436 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_727
timestamp 1649977179
transform 1 0 67988 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_729
timestamp 1649977179
transform 1 0 68172 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1649977179
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1649977179
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1649977179
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1649977179
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1649977179
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1649977179
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1649977179
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1649977179
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1649977179
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1649977179
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1649977179
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1649977179
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1649977179
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1649977179
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1649977179
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1649977179
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1649977179
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1649977179
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1649977179
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1649977179
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1649977179
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1649977179
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1649977179
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1649977179
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1649977179
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1649977179
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1649977179
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1649977179
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1649977179
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1649977179
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1649977179
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1649977179
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1649977179
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1649977179
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1649977179
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1649977179
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1649977179
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1649977179
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1649977179
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1649977179
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1649977179
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1649977179
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1649977179
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1649977179
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1649977179
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1649977179
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1649977179
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1649977179
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1649977179
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1649977179
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1649977179
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1649977179
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1649977179
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1649977179
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_513
timestamp 1649977179
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1649977179
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1649977179
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_533
timestamp 1649977179
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_545
timestamp 1649977179
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_557
timestamp 1649977179
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_569
timestamp 1649977179
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1649977179
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1649977179
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_589
timestamp 1649977179
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_601
timestamp 1649977179
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_613
timestamp 1649977179
transform 1 0 57500 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_625
timestamp 1649977179
transform 1 0 58604 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_637
timestamp 1649977179
transform 1 0 59708 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_643
timestamp 1649977179
transform 1 0 60260 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_645
timestamp 1649977179
transform 1 0 60444 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_657
timestamp 1649977179
transform 1 0 61548 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_669
timestamp 1649977179
transform 1 0 62652 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_681
timestamp 1649977179
transform 1 0 63756 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_693
timestamp 1649977179
transform 1 0 64860 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_699
timestamp 1649977179
transform 1 0 65412 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_701
timestamp 1649977179
transform 1 0 65596 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_713
timestamp 1649977179
transform 1 0 66700 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_725
timestamp 1649977179
transform 1 0 67804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_729
timestamp 1649977179
transform 1 0 68172 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1649977179
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1649977179
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1649977179
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1649977179
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1649977179
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1649977179
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1649977179
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1649977179
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1649977179
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1649977179
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1649977179
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1649977179
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1649977179
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1649977179
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1649977179
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1649977179
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1649977179
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1649977179
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1649977179
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1649977179
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1649977179
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1649977179
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1649977179
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1649977179
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1649977179
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1649977179
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1649977179
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1649977179
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1649977179
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1649977179
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1649977179
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1649977179
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1649977179
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1649977179
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1649977179
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1649977179
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1649977179
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1649977179
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1649977179
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1649977179
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1649977179
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1649977179
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1649977179
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1649977179
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1649977179
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1649977179
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1649977179
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1649977179
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1649977179
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1649977179
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1649977179
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1649977179
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1649977179
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1649977179
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1649977179
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_517
timestamp 1649977179
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_529
timestamp 1649977179
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_541
timestamp 1649977179
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1649977179
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1649977179
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_561
timestamp 1649977179
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_573
timestamp 1649977179
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_585
timestamp 1649977179
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_597
timestamp 1649977179
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1649977179
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1649977179
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_617
timestamp 1649977179
transform 1 0 57868 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_629
timestamp 1649977179
transform 1 0 58972 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_641
timestamp 1649977179
transform 1 0 60076 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_653
timestamp 1649977179
transform 1 0 61180 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_665
timestamp 1649977179
transform 1 0 62284 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_671
timestamp 1649977179
transform 1 0 62836 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_673
timestamp 1649977179
transform 1 0 63020 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_685
timestamp 1649977179
transform 1 0 64124 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_697
timestamp 1649977179
transform 1 0 65228 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_709
timestamp 1649977179
transform 1 0 66332 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_721
timestamp 1649977179
transform 1 0 67436 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_727
timestamp 1649977179
transform 1 0 67988 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_729
timestamp 1649977179
transform 1 0 68172 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1649977179
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1649977179
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1649977179
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1649977179
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1649977179
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1649977179
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1649977179
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1649977179
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1649977179
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1649977179
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1649977179
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1649977179
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1649977179
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1649977179
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1649977179
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1649977179
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1649977179
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1649977179
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1649977179
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1649977179
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1649977179
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1649977179
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1649977179
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1649977179
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1649977179
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1649977179
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1649977179
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1649977179
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1649977179
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1649977179
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1649977179
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1649977179
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1649977179
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1649977179
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1649977179
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1649977179
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1649977179
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1649977179
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1649977179
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1649977179
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1649977179
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1649977179
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_401
timestamp 1649977179
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1649977179
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1649977179
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1649977179
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1649977179
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1649977179
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1649977179
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1649977179
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1649977179
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1649977179
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1649977179
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1649977179
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1649977179
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1649977179
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1649977179
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_533
timestamp 1649977179
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_545
timestamp 1649977179
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_557
timestamp 1649977179
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_569
timestamp 1649977179
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1649977179
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1649977179
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_589
timestamp 1649977179
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_601
timestamp 1649977179
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_613
timestamp 1649977179
transform 1 0 57500 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_625
timestamp 1649977179
transform 1 0 58604 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_637
timestamp 1649977179
transform 1 0 59708 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_643
timestamp 1649977179
transform 1 0 60260 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_645
timestamp 1649977179
transform 1 0 60444 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_657
timestamp 1649977179
transform 1 0 61548 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_669
timestamp 1649977179
transform 1 0 62652 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_681
timestamp 1649977179
transform 1 0 63756 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_693
timestamp 1649977179
transform 1 0 64860 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_699
timestamp 1649977179
transform 1 0 65412 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_701
timestamp 1649977179
transform 1 0 65596 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_713
timestamp 1649977179
transform 1 0 66700 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_725
timestamp 1649977179
transform 1 0 67804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_729
timestamp 1649977179
transform 1 0 68172 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1649977179
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1649977179
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1649977179
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1649977179
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1649977179
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1649977179
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1649977179
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1649977179
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1649977179
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1649977179
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1649977179
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1649977179
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1649977179
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1649977179
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1649977179
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1649977179
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1649977179
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1649977179
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1649977179
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1649977179
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1649977179
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1649977179
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1649977179
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1649977179
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1649977179
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1649977179
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1649977179
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1649977179
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1649977179
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1649977179
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1649977179
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1649977179
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1649977179
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1649977179
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1649977179
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1649977179
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1649977179
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1649977179
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1649977179
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1649977179
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1649977179
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1649977179
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1649977179
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1649977179
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1649977179
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1649977179
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1649977179
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1649977179
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1649977179
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1649977179
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1649977179
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1649977179
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1649977179
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1649977179
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1649977179
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_517
timestamp 1649977179
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_529
timestamp 1649977179
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_541
timestamp 1649977179
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1649977179
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1649977179
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_561
timestamp 1649977179
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_573
timestamp 1649977179
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_585
timestamp 1649977179
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_597
timestamp 1649977179
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 1649977179
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1649977179
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_617
timestamp 1649977179
transform 1 0 57868 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_629
timestamp 1649977179
transform 1 0 58972 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_641
timestamp 1649977179
transform 1 0 60076 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_653
timestamp 1649977179
transform 1 0 61180 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_665
timestamp 1649977179
transform 1 0 62284 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_671
timestamp 1649977179
transform 1 0 62836 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_673
timestamp 1649977179
transform 1 0 63020 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_685
timestamp 1649977179
transform 1 0 64124 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_697
timestamp 1649977179
transform 1 0 65228 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_709
timestamp 1649977179
transform 1 0 66332 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_721
timestamp 1649977179
transform 1 0 67436 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_727
timestamp 1649977179
transform 1 0 67988 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_729
timestamp 1649977179
transform 1 0 68172 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1649977179
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1649977179
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1649977179
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1649977179
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1649977179
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1649977179
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1649977179
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1649977179
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1649977179
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1649977179
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1649977179
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1649977179
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1649977179
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1649977179
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1649977179
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1649977179
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1649977179
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1649977179
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1649977179
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1649977179
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1649977179
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1649977179
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1649977179
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_221
timestamp 1649977179
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_233
timestamp 1649977179
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1649977179
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1649977179
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1649977179
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1649977179
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_277
timestamp 1649977179
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_289
timestamp 1649977179
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1649977179
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1649977179
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1649977179
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1649977179
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_333
timestamp 1649977179
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_345
timestamp 1649977179
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1649977179
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1649977179
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1649977179
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1649977179
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_389
timestamp 1649977179
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_401
timestamp 1649977179
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1649977179
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1649977179
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1649977179
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1649977179
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1649977179
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1649977179
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1649977179
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1649977179
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1649977179
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1649977179
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1649977179
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_513
timestamp 1649977179
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1649977179
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1649977179
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_533
timestamp 1649977179
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_545
timestamp 1649977179
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_557
timestamp 1649977179
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_569
timestamp 1649977179
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_581
timestamp 1649977179
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1649977179
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_589
timestamp 1649977179
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_601
timestamp 1649977179
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_613
timestamp 1649977179
transform 1 0 57500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_625
timestamp 1649977179
transform 1 0 58604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_637
timestamp 1649977179
transform 1 0 59708 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_643
timestamp 1649977179
transform 1 0 60260 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_645
timestamp 1649977179
transform 1 0 60444 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_657
timestamp 1649977179
transform 1 0 61548 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_669
timestamp 1649977179
transform 1 0 62652 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_681
timestamp 1649977179
transform 1 0 63756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_693
timestamp 1649977179
transform 1 0 64860 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_699
timestamp 1649977179
transform 1 0 65412 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_701
timestamp 1649977179
transform 1 0 65596 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_713
timestamp 1649977179
transform 1 0 66700 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_725
timestamp 1649977179
transform 1 0 67804 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1649977179
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1649977179
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1649977179
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1649977179
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1649977179
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1649977179
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1649977179
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1649977179
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1649977179
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1649977179
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1649977179
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1649977179
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1649977179
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1649977179
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1649977179
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1649977179
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1649977179
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1649977179
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1649977179
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1649977179
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1649977179
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1649977179
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1649977179
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1649977179
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1649977179
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1649977179
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_249
timestamp 1649977179
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_261
timestamp 1649977179
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1649977179
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1649977179
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1649977179
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_293
timestamp 1649977179
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_305
timestamp 1649977179
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_317
timestamp 1649977179
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1649977179
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1649977179
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_337
timestamp 1649977179
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_349
timestamp 1649977179
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_361
timestamp 1649977179
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_373
timestamp 1649977179
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1649977179
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1649977179
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1649977179
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1649977179
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1649977179
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1649977179
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1649977179
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1649977179
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1649977179
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1649977179
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1649977179
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1649977179
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1649977179
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1649977179
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1649977179
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_517
timestamp 1649977179
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_529
timestamp 1649977179
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_541
timestamp 1649977179
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1649977179
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1649977179
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_561
timestamp 1649977179
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_573
timestamp 1649977179
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_585
timestamp 1649977179
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_597
timestamp 1649977179
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_609
timestamp 1649977179
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1649977179
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_617
timestamp 1649977179
transform 1 0 57868 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_629
timestamp 1649977179
transform 1 0 58972 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_641
timestamp 1649977179
transform 1 0 60076 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_653
timestamp 1649977179
transform 1 0 61180 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_665
timestamp 1649977179
transform 1 0 62284 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_671
timestamp 1649977179
transform 1 0 62836 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_673
timestamp 1649977179
transform 1 0 63020 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_685
timestamp 1649977179
transform 1 0 64124 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_697
timestamp 1649977179
transform 1 0 65228 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_709
timestamp 1649977179
transform 1 0 66332 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_724
timestamp 1649977179
transform 1 0 67712 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_729
timestamp 1649977179
transform 1 0 68172 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1649977179
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1649977179
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1649977179
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1649977179
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1649977179
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1649977179
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1649977179
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1649977179
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1649977179
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1649977179
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1649977179
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1649977179
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1649977179
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1649977179
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1649977179
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1649977179
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1649977179
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1649977179
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1649977179
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1649977179
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1649977179
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1649977179
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1649977179
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1649977179
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_233
timestamp 1649977179
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1649977179
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1649977179
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1649977179
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_265
timestamp 1649977179
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_277
timestamp 1649977179
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_289
timestamp 1649977179
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1649977179
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1649977179
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1649977179
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_321
timestamp 1649977179
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_333
timestamp 1649977179
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_345
timestamp 1649977179
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1649977179
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1649977179
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1649977179
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1649977179
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1649977179
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1649977179
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1649977179
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1649977179
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1649977179
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1649977179
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1649977179
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1649977179
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1649977179
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1649977179
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1649977179
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1649977179
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1649977179
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_513
timestamp 1649977179
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1649977179
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1649977179
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_533
timestamp 1649977179
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_545
timestamp 1649977179
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_557
timestamp 1649977179
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_569
timestamp 1649977179
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_581
timestamp 1649977179
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1649977179
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_589
timestamp 1649977179
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_601
timestamp 1649977179
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_613
timestamp 1649977179
transform 1 0 57500 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_625
timestamp 1649977179
transform 1 0 58604 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_637
timestamp 1649977179
transform 1 0 59708 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_643
timestamp 1649977179
transform 1 0 60260 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_645
timestamp 1649977179
transform 1 0 60444 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_657
timestamp 1649977179
transform 1 0 61548 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_669
timestamp 1649977179
transform 1 0 62652 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_681
timestamp 1649977179
transform 1 0 63756 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_693
timestamp 1649977179
transform 1 0 64860 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_699
timestamp 1649977179
transform 1 0 65412 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_701
timestamp 1649977179
transform 1 0 65596 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_713
timestamp 1649977179
transform 1 0 66700 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_725
timestamp 1649977179
transform 1 0 67804 0 1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1649977179
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1649977179
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1649977179
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1649977179
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1649977179
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1649977179
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1649977179
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1649977179
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1649977179
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1649977179
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1649977179
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1649977179
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1649977179
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1649977179
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1649977179
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1649977179
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1649977179
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1649977179
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1649977179
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1649977179
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1649977179
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1649977179
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1649977179
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1649977179
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1649977179
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1649977179
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_249
timestamp 1649977179
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_261
timestamp 1649977179
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1649977179
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1649977179
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1649977179
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_293
timestamp 1649977179
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_305
timestamp 1649977179
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_317
timestamp 1649977179
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1649977179
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1649977179
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1649977179
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_349
timestamp 1649977179
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_361
timestamp 1649977179
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_373
timestamp 1649977179
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1649977179
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1649977179
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1649977179
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1649977179
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1649977179
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1649977179
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1649977179
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1649977179
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1649977179
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1649977179
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1649977179
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1649977179
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1649977179
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1649977179
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_505
timestamp 1649977179
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_517
timestamp 1649977179
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_529
timestamp 1649977179
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_541
timestamp 1649977179
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1649977179
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1649977179
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_561
timestamp 1649977179
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_573
timestamp 1649977179
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_585
timestamp 1649977179
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_597
timestamp 1649977179
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_609
timestamp 1649977179
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1649977179
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_617
timestamp 1649977179
transform 1 0 57868 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_629
timestamp 1649977179
transform 1 0 58972 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_641
timestamp 1649977179
transform 1 0 60076 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_653
timestamp 1649977179
transform 1 0 61180 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_665
timestamp 1649977179
transform 1 0 62284 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_671
timestamp 1649977179
transform 1 0 62836 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_673
timestamp 1649977179
transform 1 0 63020 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_685
timestamp 1649977179
transform 1 0 64124 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_697
timestamp 1649977179
transform 1 0 65228 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_709
timestamp 1649977179
transform 1 0 66332 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_724
timestamp 1649977179
transform 1 0 67712 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_729
timestamp 1649977179
transform 1 0 68172 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1649977179
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1649977179
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1649977179
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1649977179
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1649977179
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1649977179
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1649977179
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1649977179
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1649977179
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1649977179
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1649977179
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1649977179
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1649977179
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1649977179
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1649977179
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1649977179
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1649977179
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1649977179
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1649977179
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1649977179
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1649977179
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1649977179
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1649977179
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1649977179
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1649977179
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1649977179
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1649977179
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1649977179
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1649977179
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_277
timestamp 1649977179
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_289
timestamp 1649977179
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1649977179
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1649977179
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1649977179
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_321
timestamp 1649977179
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_333
timestamp 1649977179
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_345
timestamp 1649977179
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1649977179
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1649977179
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1649977179
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1649977179
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1649977179
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_401
timestamp 1649977179
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1649977179
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1649977179
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1649977179
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1649977179
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1649977179
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1649977179
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1649977179
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1649977179
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1649977179
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1649977179
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1649977179
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_513
timestamp 1649977179
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_525
timestamp 1649977179
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_531
timestamp 1649977179
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_533
timestamp 1649977179
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_545
timestamp 1649977179
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_557
timestamp 1649977179
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_569
timestamp 1649977179
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_581
timestamp 1649977179
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_587
timestamp 1649977179
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_589
timestamp 1649977179
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_601
timestamp 1649977179
transform 1 0 56396 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_613
timestamp 1649977179
transform 1 0 57500 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_625
timestamp 1649977179
transform 1 0 58604 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_637
timestamp 1649977179
transform 1 0 59708 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_643
timestamp 1649977179
transform 1 0 60260 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_645
timestamp 1649977179
transform 1 0 60444 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_657
timestamp 1649977179
transform 1 0 61548 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_669
timestamp 1649977179
transform 1 0 62652 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_681
timestamp 1649977179
transform 1 0 63756 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_693
timestamp 1649977179
transform 1 0 64860 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_699
timestamp 1649977179
transform 1 0 65412 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_701
timestamp 1649977179
transform 1 0 65596 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_713
timestamp 1649977179
transform 1 0 66700 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_725
timestamp 1649977179
transform 1 0 67804 0 1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1649977179
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1649977179
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1649977179
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1649977179
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1649977179
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1649977179
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1649977179
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1649977179
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1649977179
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1649977179
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1649977179
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1649977179
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1649977179
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1649977179
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1649977179
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1649977179
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1649977179
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1649977179
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1649977179
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1649977179
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1649977179
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1649977179
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1649977179
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1649977179
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1649977179
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1649977179
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1649977179
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_261
timestamp 1649977179
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1649977179
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1649977179
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_281
timestamp 1649977179
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_293
timestamp 1649977179
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_305
timestamp 1649977179
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_317
timestamp 1649977179
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1649977179
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1649977179
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1649977179
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1649977179
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1649977179
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1649977179
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1649977179
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1649977179
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1649977179
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1649977179
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1649977179
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1649977179
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1649977179
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1649977179
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1649977179
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1649977179
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1649977179
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1649977179
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1649977179
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1649977179
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_505
timestamp 1649977179
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_517
timestamp 1649977179
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_529
timestamp 1649977179
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_541
timestamp 1649977179
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 1649977179
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1649977179
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_561
timestamp 1649977179
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_573
timestamp 1649977179
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_585
timestamp 1649977179
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_597
timestamp 1649977179
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_609
timestamp 1649977179
transform 1 0 57132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_615
timestamp 1649977179
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_617
timestamp 1649977179
transform 1 0 57868 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_629
timestamp 1649977179
transform 1 0 58972 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_641
timestamp 1649977179
transform 1 0 60076 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_653
timestamp 1649977179
transform 1 0 61180 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_665
timestamp 1649977179
transform 1 0 62284 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_671
timestamp 1649977179
transform 1 0 62836 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_673
timestamp 1649977179
transform 1 0 63020 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_685
timestamp 1649977179
transform 1 0 64124 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_697
timestamp 1649977179
transform 1 0 65228 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_709
timestamp 1649977179
transform 1 0 66332 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_721
timestamp 1649977179
transform 1 0 67436 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_727
timestamp 1649977179
transform 1 0 67988 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_729
timestamp 1649977179
transform 1 0 68172 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1649977179
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1649977179
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1649977179
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1649977179
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1649977179
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1649977179
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1649977179
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1649977179
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1649977179
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1649977179
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1649977179
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1649977179
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1649977179
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1649977179
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1649977179
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1649977179
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1649977179
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1649977179
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1649977179
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1649977179
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1649977179
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1649977179
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1649977179
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1649977179
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1649977179
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1649977179
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1649977179
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1649977179
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_265
timestamp 1649977179
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_277
timestamp 1649977179
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_289
timestamp 1649977179
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1649977179
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1649977179
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1649977179
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_321
timestamp 1649977179
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_333
timestamp 1649977179
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_345
timestamp 1649977179
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1649977179
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1649977179
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1649977179
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1649977179
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1649977179
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1649977179
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1649977179
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1649977179
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1649977179
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1649977179
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1649977179
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1649977179
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1649977179
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1649977179
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1649977179
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1649977179
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1649977179
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_513
timestamp 1649977179
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_525
timestamp 1649977179
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_531
timestamp 1649977179
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_533
timestamp 1649977179
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_545
timestamp 1649977179
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_557
timestamp 1649977179
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_569
timestamp 1649977179
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_581
timestamp 1649977179
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_587
timestamp 1649977179
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_589
timestamp 1649977179
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_601
timestamp 1649977179
transform 1 0 56396 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_613
timestamp 1649977179
transform 1 0 57500 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_625
timestamp 1649977179
transform 1 0 58604 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_637
timestamp 1649977179
transform 1 0 59708 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_643
timestamp 1649977179
transform 1 0 60260 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_645
timestamp 1649977179
transform 1 0 60444 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_657
timestamp 1649977179
transform 1 0 61548 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_669
timestamp 1649977179
transform 1 0 62652 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_681
timestamp 1649977179
transform 1 0 63756 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_693
timestamp 1649977179
transform 1 0 64860 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_699
timestamp 1649977179
transform 1 0 65412 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_701
timestamp 1649977179
transform 1 0 65596 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_713
timestamp 1649977179
transform 1 0 66700 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_725
timestamp 1649977179
transform 1 0 67804 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_729
timestamp 1649977179
transform 1 0 68172 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1649977179
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1649977179
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1649977179
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1649977179
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1649977179
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1649977179
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1649977179
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1649977179
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1649977179
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1649977179
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1649977179
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1649977179
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1649977179
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1649977179
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1649977179
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1649977179
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1649977179
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1649977179
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1649977179
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1649977179
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1649977179
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1649977179
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1649977179
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1649977179
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1649977179
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1649977179
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_249
timestamp 1649977179
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_261
timestamp 1649977179
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1649977179
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1649977179
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_281
timestamp 1649977179
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_293
timestamp 1649977179
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_305
timestamp 1649977179
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_317
timestamp 1649977179
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1649977179
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1649977179
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1649977179
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1649977179
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1649977179
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1649977179
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1649977179
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1649977179
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1649977179
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1649977179
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1649977179
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1649977179
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1649977179
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1649977179
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1649977179
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1649977179
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1649977179
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1649977179
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1649977179
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1649977179
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_505
timestamp 1649977179
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_517
timestamp 1649977179
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_529
timestamp 1649977179
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_541
timestamp 1649977179
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_553
timestamp 1649977179
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_559
timestamp 1649977179
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_561
timestamp 1649977179
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_573
timestamp 1649977179
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_585
timestamp 1649977179
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_597
timestamp 1649977179
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_609
timestamp 1649977179
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_615
timestamp 1649977179
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_617
timestamp 1649977179
transform 1 0 57868 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_629
timestamp 1649977179
transform 1 0 58972 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_641
timestamp 1649977179
transform 1 0 60076 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_653
timestamp 1649977179
transform 1 0 61180 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_665
timestamp 1649977179
transform 1 0 62284 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_671
timestamp 1649977179
transform 1 0 62836 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_673
timestamp 1649977179
transform 1 0 63020 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_685
timestamp 1649977179
transform 1 0 64124 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_697
timestamp 1649977179
transform 1 0 65228 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_709
timestamp 1649977179
transform 1 0 66332 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_721
timestamp 1649977179
transform 1 0 67436 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_727
timestamp 1649977179
transform 1 0 67988 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_729
timestamp 1649977179
transform 1 0 68172 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1649977179
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1649977179
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1649977179
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1649977179
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1649977179
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1649977179
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1649977179
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1649977179
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1649977179
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1649977179
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1649977179
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1649977179
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1649977179
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1649977179
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1649977179
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1649977179
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1649977179
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1649977179
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1649977179
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1649977179
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1649977179
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1649977179
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1649977179
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1649977179
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1649977179
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1649977179
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1649977179
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1649977179
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_265
timestamp 1649977179
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_277
timestamp 1649977179
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_289
timestamp 1649977179
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1649977179
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1649977179
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1649977179
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_321
timestamp 1649977179
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_333
timestamp 1649977179
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_345
timestamp 1649977179
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1649977179
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1649977179
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1649977179
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_377
timestamp 1649977179
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_389
timestamp 1649977179
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_401
timestamp 1649977179
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1649977179
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1649977179
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1649977179
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1649977179
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1649977179
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1649977179
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1649977179
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1649977179
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1649977179
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1649977179
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1649977179
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_513
timestamp 1649977179
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_525
timestamp 1649977179
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_531
timestamp 1649977179
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_533
timestamp 1649977179
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_545
timestamp 1649977179
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_557
timestamp 1649977179
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_569
timestamp 1649977179
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_581
timestamp 1649977179
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_587
timestamp 1649977179
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_589
timestamp 1649977179
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_601
timestamp 1649977179
transform 1 0 56396 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_613
timestamp 1649977179
transform 1 0 57500 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_625
timestamp 1649977179
transform 1 0 58604 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_637
timestamp 1649977179
transform 1 0 59708 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_643
timestamp 1649977179
transform 1 0 60260 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_645
timestamp 1649977179
transform 1 0 60444 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_657
timestamp 1649977179
transform 1 0 61548 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_669
timestamp 1649977179
transform 1 0 62652 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_681
timestamp 1649977179
transform 1 0 63756 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_693
timestamp 1649977179
transform 1 0 64860 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_699
timestamp 1649977179
transform 1 0 65412 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_701
timestamp 1649977179
transform 1 0 65596 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_713
timestamp 1649977179
transform 1 0 66700 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_725
timestamp 1649977179
transform 1 0 67804 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_729
timestamp 1649977179
transform 1 0 68172 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1649977179
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1649977179
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1649977179
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1649977179
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1649977179
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1649977179
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1649977179
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1649977179
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1649977179
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1649977179
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1649977179
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1649977179
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1649977179
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1649977179
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1649977179
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1649977179
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1649977179
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1649977179
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1649977179
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1649977179
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1649977179
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1649977179
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1649977179
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1649977179
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1649977179
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1649977179
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1649977179
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_261
timestamp 1649977179
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1649977179
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1649977179
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_281
timestamp 1649977179
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_293
timestamp 1649977179
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_305
timestamp 1649977179
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_317
timestamp 1649977179
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1649977179
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1649977179
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1649977179
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_349
timestamp 1649977179
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_361
timestamp 1649977179
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_373
timestamp 1649977179
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1649977179
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1649977179
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1649977179
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1649977179
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1649977179
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1649977179
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1649977179
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1649977179
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1649977179
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1649977179
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1649977179
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1649977179
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1649977179
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1649977179
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_505
timestamp 1649977179
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_517
timestamp 1649977179
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_529
timestamp 1649977179
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_541
timestamp 1649977179
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_553
timestamp 1649977179
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_559
timestamp 1649977179
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_561
timestamp 1649977179
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_573
timestamp 1649977179
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_585
timestamp 1649977179
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_597
timestamp 1649977179
transform 1 0 56028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_609
timestamp 1649977179
transform 1 0 57132 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_615
timestamp 1649977179
transform 1 0 57684 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_617
timestamp 1649977179
transform 1 0 57868 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_629
timestamp 1649977179
transform 1 0 58972 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_641
timestamp 1649977179
transform 1 0 60076 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_653
timestamp 1649977179
transform 1 0 61180 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_665
timestamp 1649977179
transform 1 0 62284 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_671
timestamp 1649977179
transform 1 0 62836 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_673
timestamp 1649977179
transform 1 0 63020 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_685
timestamp 1649977179
transform 1 0 64124 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_697
timestamp 1649977179
transform 1 0 65228 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_709
timestamp 1649977179
transform 1 0 66332 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_721
timestamp 1649977179
transform 1 0 67436 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_727
timestamp 1649977179
transform 1 0 67988 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_729
timestamp 1649977179
transform 1 0 68172 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1649977179
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1649977179
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1649977179
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1649977179
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1649977179
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1649977179
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1649977179
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1649977179
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1649977179
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1649977179
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1649977179
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1649977179
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1649977179
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1649977179
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1649977179
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1649977179
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1649977179
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1649977179
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1649977179
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1649977179
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1649977179
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1649977179
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1649977179
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1649977179
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1649977179
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1649977179
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1649977179
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1649977179
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_265
timestamp 1649977179
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_277
timestamp 1649977179
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_289
timestamp 1649977179
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1649977179
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1649977179
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1649977179
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1649977179
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_333
timestamp 1649977179
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_345
timestamp 1649977179
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1649977179
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1649977179
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_365
timestamp 1649977179
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_377
timestamp 1649977179
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_389
timestamp 1649977179
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_401
timestamp 1649977179
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1649977179
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1649977179
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1649977179
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1649977179
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1649977179
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1649977179
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1649977179
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1649977179
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1649977179
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1649977179
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1649977179
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_513
timestamp 1649977179
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_525
timestamp 1649977179
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_531
timestamp 1649977179
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_533
timestamp 1649977179
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_545
timestamp 1649977179
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_557
timestamp 1649977179
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_569
timestamp 1649977179
transform 1 0 53452 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_581
timestamp 1649977179
transform 1 0 54556 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_587
timestamp 1649977179
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_589
timestamp 1649977179
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_601
timestamp 1649977179
transform 1 0 56396 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_613
timestamp 1649977179
transform 1 0 57500 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_625
timestamp 1649977179
transform 1 0 58604 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_637
timestamp 1649977179
transform 1 0 59708 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_643
timestamp 1649977179
transform 1 0 60260 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_645
timestamp 1649977179
transform 1 0 60444 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_657
timestamp 1649977179
transform 1 0 61548 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_669
timestamp 1649977179
transform 1 0 62652 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_681
timestamp 1649977179
transform 1 0 63756 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_693
timestamp 1649977179
transform 1 0 64860 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_699
timestamp 1649977179
transform 1 0 65412 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_701
timestamp 1649977179
transform 1 0 65596 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_713
timestamp 1649977179
transform 1 0 66700 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_725
timestamp 1649977179
transform 1 0 67804 0 1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1649977179
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1649977179
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1649977179
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1649977179
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1649977179
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1649977179
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1649977179
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1649977179
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1649977179
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1649977179
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1649977179
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1649977179
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1649977179
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1649977179
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1649977179
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1649977179
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1649977179
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1649977179
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1649977179
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1649977179
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1649977179
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1649977179
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1649977179
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1649977179
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1649977179
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1649977179
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1649977179
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_261
timestamp 1649977179
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1649977179
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1649977179
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1649977179
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_293
timestamp 1649977179
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_305
timestamp 1649977179
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_317
timestamp 1649977179
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1649977179
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1649977179
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1649977179
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_349
timestamp 1649977179
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_361
timestamp 1649977179
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_373
timestamp 1649977179
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1649977179
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1649977179
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1649977179
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1649977179
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1649977179
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1649977179
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1649977179
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1649977179
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1649977179
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1649977179
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1649977179
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1649977179
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1649977179
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1649977179
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_505
timestamp 1649977179
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_517
timestamp 1649977179
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_529
timestamp 1649977179
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_541
timestamp 1649977179
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_553
timestamp 1649977179
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_559
timestamp 1649977179
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_561
timestamp 1649977179
transform 1 0 52716 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_573
timestamp 1649977179
transform 1 0 53820 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_585
timestamp 1649977179
transform 1 0 54924 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_597
timestamp 1649977179
transform 1 0 56028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_609
timestamp 1649977179
transform 1 0 57132 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_615
timestamp 1649977179
transform 1 0 57684 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_617
timestamp 1649977179
transform 1 0 57868 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_629
timestamp 1649977179
transform 1 0 58972 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_641
timestamp 1649977179
transform 1 0 60076 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_653
timestamp 1649977179
transform 1 0 61180 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_665
timestamp 1649977179
transform 1 0 62284 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_671
timestamp 1649977179
transform 1 0 62836 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_673
timestamp 1649977179
transform 1 0 63020 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_685
timestamp 1649977179
transform 1 0 64124 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_697
timestamp 1649977179
transform 1 0 65228 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_709
timestamp 1649977179
transform 1 0 66332 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_724
timestamp 1649977179
transform 1 0 67712 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_729
timestamp 1649977179
transform 1 0 68172 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1649977179
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1649977179
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1649977179
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1649977179
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1649977179
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1649977179
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1649977179
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1649977179
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1649977179
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1649977179
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1649977179
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1649977179
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1649977179
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1649977179
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1649977179
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1649977179
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1649977179
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1649977179
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1649977179
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1649977179
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1649977179
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1649977179
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1649977179
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1649977179
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1649977179
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1649977179
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1649977179
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1649977179
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1649977179
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_277
timestamp 1649977179
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_289
timestamp 1649977179
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1649977179
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1649977179
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1649977179
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_321
timestamp 1649977179
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_333
timestamp 1649977179
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_345
timestamp 1649977179
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1649977179
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1649977179
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1649977179
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1649977179
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_389
timestamp 1649977179
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_401
timestamp 1649977179
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1649977179
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1649977179
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1649977179
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1649977179
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1649977179
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1649977179
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1649977179
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1649977179
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1649977179
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1649977179
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1649977179
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_513
timestamp 1649977179
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_525
timestamp 1649977179
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_531
timestamp 1649977179
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_533
timestamp 1649977179
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_545
timestamp 1649977179
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_557
timestamp 1649977179
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_569
timestamp 1649977179
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_581
timestamp 1649977179
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_587
timestamp 1649977179
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_589
timestamp 1649977179
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_601
timestamp 1649977179
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_613
timestamp 1649977179
transform 1 0 57500 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_625
timestamp 1649977179
transform 1 0 58604 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_637
timestamp 1649977179
transform 1 0 59708 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_643
timestamp 1649977179
transform 1 0 60260 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_645
timestamp 1649977179
transform 1 0 60444 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_657
timestamp 1649977179
transform 1 0 61548 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_669
timestamp 1649977179
transform 1 0 62652 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_681
timestamp 1649977179
transform 1 0 63756 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_693
timestamp 1649977179
transform 1 0 64860 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_699
timestamp 1649977179
transform 1 0 65412 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_701
timestamp 1649977179
transform 1 0 65596 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_713
timestamp 1649977179
transform 1 0 66700 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_725
timestamp 1649977179
transform 1 0 67804 0 1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1649977179
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1649977179
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1649977179
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1649977179
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1649977179
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1649977179
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1649977179
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1649977179
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1649977179
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1649977179
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1649977179
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1649977179
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1649977179
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1649977179
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1649977179
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1649977179
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1649977179
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1649977179
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1649977179
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1649977179
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1649977179
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1649977179
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1649977179
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1649977179
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1649977179
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1649977179
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_249
timestamp 1649977179
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_261
timestamp 1649977179
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1649977179
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1649977179
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1649977179
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1649977179
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1649977179
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1649977179
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1649977179
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1649977179
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1649977179
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1649977179
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1649977179
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_373
timestamp 1649977179
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1649977179
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1649977179
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1649977179
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_405
timestamp 1649977179
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_417
timestamp 1649977179
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_429
timestamp 1649977179
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1649977179
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1649977179
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1649977179
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1649977179
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1649977179
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1649977179
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1649977179
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1649977179
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_505
timestamp 1649977179
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_517
timestamp 1649977179
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_529
timestamp 1649977179
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_541
timestamp 1649977179
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_553
timestamp 1649977179
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_559
timestamp 1649977179
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_561
timestamp 1649977179
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_573
timestamp 1649977179
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_585
timestamp 1649977179
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_597
timestamp 1649977179
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_609
timestamp 1649977179
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_615
timestamp 1649977179
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_617
timestamp 1649977179
transform 1 0 57868 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_629
timestamp 1649977179
transform 1 0 58972 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_641
timestamp 1649977179
transform 1 0 60076 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_653
timestamp 1649977179
transform 1 0 61180 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_665
timestamp 1649977179
transform 1 0 62284 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_671
timestamp 1649977179
transform 1 0 62836 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_673
timestamp 1649977179
transform 1 0 63020 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_685
timestamp 1649977179
transform 1 0 64124 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_697
timestamp 1649977179
transform 1 0 65228 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_709
timestamp 1649977179
transform 1 0 66332 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_724
timestamp 1649977179
transform 1 0 67712 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_729
timestamp 1649977179
transform 1 0 68172 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1649977179
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1649977179
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1649977179
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1649977179
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1649977179
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1649977179
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1649977179
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1649977179
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1649977179
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1649977179
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1649977179
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1649977179
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1649977179
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1649977179
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1649977179
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1649977179
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1649977179
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1649977179
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1649977179
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1649977179
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1649977179
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1649977179
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1649977179
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1649977179
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1649977179
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1649977179
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1649977179
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1649977179
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1649977179
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_277
timestamp 1649977179
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_289
timestamp 1649977179
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1649977179
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1649977179
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1649977179
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1649977179
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1649977179
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1649977179
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1649977179
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1649977179
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 1649977179
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_377
timestamp 1649977179
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_389
timestamp 1649977179
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_401
timestamp 1649977179
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1649977179
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1649977179
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1649977179
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1649977179
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1649977179
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1649977179
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1649977179
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1649977179
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1649977179
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1649977179
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1649977179
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_513
timestamp 1649977179
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_525
timestamp 1649977179
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_531
timestamp 1649977179
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_533
timestamp 1649977179
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_545
timestamp 1649977179
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_557
timestamp 1649977179
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_569
timestamp 1649977179
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_581
timestamp 1649977179
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_587
timestamp 1649977179
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_589
timestamp 1649977179
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_601
timestamp 1649977179
transform 1 0 56396 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_613
timestamp 1649977179
transform 1 0 57500 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_625
timestamp 1649977179
transform 1 0 58604 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_637
timestamp 1649977179
transform 1 0 59708 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_643
timestamp 1649977179
transform 1 0 60260 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_645
timestamp 1649977179
transform 1 0 60444 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_657
timestamp 1649977179
transform 1 0 61548 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_669
timestamp 1649977179
transform 1 0 62652 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_681
timestamp 1649977179
transform 1 0 63756 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_693
timestamp 1649977179
transform 1 0 64860 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_699
timestamp 1649977179
transform 1 0 65412 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_701
timestamp 1649977179
transform 1 0 65596 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_713
timestamp 1649977179
transform 1 0 66700 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_725
timestamp 1649977179
transform 1 0 67804 0 1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1649977179
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1649977179
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1649977179
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1649977179
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1649977179
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1649977179
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1649977179
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1649977179
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1649977179
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1649977179
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1649977179
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1649977179
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1649977179
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1649977179
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1649977179
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1649977179
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1649977179
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1649977179
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1649977179
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1649977179
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1649977179
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1649977179
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1649977179
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1649977179
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1649977179
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1649977179
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1649977179
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 1649977179
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1649977179
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1649977179
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1649977179
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1649977179
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_305
timestamp 1649977179
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_317
timestamp 1649977179
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1649977179
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1649977179
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_337
timestamp 1649977179
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_349
timestamp 1649977179
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1649977179
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_373
timestamp 1649977179
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1649977179
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1649977179
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_393
timestamp 1649977179
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_405
timestamp 1649977179
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_417
timestamp 1649977179
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_429
timestamp 1649977179
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1649977179
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1649977179
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1649977179
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1649977179
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1649977179
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1649977179
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1649977179
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1649977179
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_505
timestamp 1649977179
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_517
timestamp 1649977179
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_529
timestamp 1649977179
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_541
timestamp 1649977179
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_553
timestamp 1649977179
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_559
timestamp 1649977179
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_561
timestamp 1649977179
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_573
timestamp 1649977179
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_585
timestamp 1649977179
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_597
timestamp 1649977179
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_609
timestamp 1649977179
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_615
timestamp 1649977179
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_617
timestamp 1649977179
transform 1 0 57868 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_629
timestamp 1649977179
transform 1 0 58972 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_641
timestamp 1649977179
transform 1 0 60076 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_653
timestamp 1649977179
transform 1 0 61180 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_665
timestamp 1649977179
transform 1 0 62284 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_671
timestamp 1649977179
transform 1 0 62836 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_673
timestamp 1649977179
transform 1 0 63020 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_685
timestamp 1649977179
transform 1 0 64124 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_697
timestamp 1649977179
transform 1 0 65228 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_709
timestamp 1649977179
transform 1 0 66332 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_721
timestamp 1649977179
transform 1 0 67436 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_727
timestamp 1649977179
transform 1 0 67988 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_729
timestamp 1649977179
transform 1 0 68172 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1649977179
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1649977179
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1649977179
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1649977179
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1649977179
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1649977179
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1649977179
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1649977179
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1649977179
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1649977179
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1649977179
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1649977179
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1649977179
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1649977179
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1649977179
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1649977179
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1649977179
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1649977179
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_177
timestamp 1649977179
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1649977179
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1649977179
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1649977179
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1649977179
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1649977179
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1649977179
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1649977179
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1649977179
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_253
timestamp 1649977179
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_265
timestamp 1649977179
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_277
timestamp 1649977179
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_289
timestamp 1649977179
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1649977179
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1649977179
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_309
timestamp 1649977179
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_321
timestamp 1649977179
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_333
timestamp 1649977179
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_345
timestamp 1649977179
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1649977179
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1649977179
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_365
timestamp 1649977179
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_377
timestamp 1649977179
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_389
timestamp 1649977179
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_401
timestamp 1649977179
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 1649977179
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1649977179
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1649977179
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1649977179
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1649977179
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1649977179
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1649977179
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1649977179
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1649977179
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1649977179
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_501
timestamp 1649977179
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_513
timestamp 1649977179
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_525
timestamp 1649977179
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 1649977179
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_533
timestamp 1649977179
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_545
timestamp 1649977179
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_557
timestamp 1649977179
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_569
timestamp 1649977179
transform 1 0 53452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_581
timestamp 1649977179
transform 1 0 54556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_587
timestamp 1649977179
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_589
timestamp 1649977179
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_601
timestamp 1649977179
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_613
timestamp 1649977179
transform 1 0 57500 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_625
timestamp 1649977179
transform 1 0 58604 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_637
timestamp 1649977179
transform 1 0 59708 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_643
timestamp 1649977179
transform 1 0 60260 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_645
timestamp 1649977179
transform 1 0 60444 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_657
timestamp 1649977179
transform 1 0 61548 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_669
timestamp 1649977179
transform 1 0 62652 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_681
timestamp 1649977179
transform 1 0 63756 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_693
timestamp 1649977179
transform 1 0 64860 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_699
timestamp 1649977179
transform 1 0 65412 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_701
timestamp 1649977179
transform 1 0 65596 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_713
timestamp 1649977179
transform 1 0 66700 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_725
timestamp 1649977179
transform 1 0 67804 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_729
timestamp 1649977179
transform 1 0 68172 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1649977179
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1649977179
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1649977179
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1649977179
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1649977179
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1649977179
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1649977179
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1649977179
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1649977179
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1649977179
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1649977179
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1649977179
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1649977179
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1649977179
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1649977179
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1649977179
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1649977179
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1649977179
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1649977179
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1649977179
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1649977179
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1649977179
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1649977179
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1649977179
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1649977179
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1649977179
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1649977179
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_261
timestamp 1649977179
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1649977179
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1649977179
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1649977179
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_293
timestamp 1649977179
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_305
timestamp 1649977179
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_317
timestamp 1649977179
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1649977179
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1649977179
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_337
timestamp 1649977179
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_349
timestamp 1649977179
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_361
timestamp 1649977179
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_373
timestamp 1649977179
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1649977179
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1649977179
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1649977179
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1649977179
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1649977179
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1649977179
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1649977179
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1649977179
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1649977179
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1649977179
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1649977179
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1649977179
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1649977179
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1649977179
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_505
timestamp 1649977179
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_517
timestamp 1649977179
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_529
timestamp 1649977179
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_541
timestamp 1649977179
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_553
timestamp 1649977179
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_559
timestamp 1649977179
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_561
timestamp 1649977179
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_573
timestamp 1649977179
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_585
timestamp 1649977179
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_597
timestamp 1649977179
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_609
timestamp 1649977179
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_615
timestamp 1649977179
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_617
timestamp 1649977179
transform 1 0 57868 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_629
timestamp 1649977179
transform 1 0 58972 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_641
timestamp 1649977179
transform 1 0 60076 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_653
timestamp 1649977179
transform 1 0 61180 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_665
timestamp 1649977179
transform 1 0 62284 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_671
timestamp 1649977179
transform 1 0 62836 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_673
timestamp 1649977179
transform 1 0 63020 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_685
timestamp 1649977179
transform 1 0 64124 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_697
timestamp 1649977179
transform 1 0 65228 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_709
timestamp 1649977179
transform 1 0 66332 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_721
timestamp 1649977179
transform 1 0 67436 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_727
timestamp 1649977179
transform 1 0 67988 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_729
timestamp 1649977179
transform 1 0 68172 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1649977179
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1649977179
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1649977179
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1649977179
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1649977179
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1649977179
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1649977179
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1649977179
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1649977179
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1649977179
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1649977179
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 1649977179
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 1649977179
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1649977179
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1649977179
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1649977179
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1649977179
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1649977179
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1649977179
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1649977179
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1649977179
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1649977179
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1649977179
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1649977179
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1649977179
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1649977179
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1649977179
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_253
timestamp 1649977179
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_265
timestamp 1649977179
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_277
timestamp 1649977179
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_289
timestamp 1649977179
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1649977179
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1649977179
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_309
timestamp 1649977179
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_321
timestamp 1649977179
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_333
timestamp 1649977179
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_345
timestamp 1649977179
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1649977179
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1649977179
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1649977179
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1649977179
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_389
timestamp 1649977179
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_401
timestamp 1649977179
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1649977179
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1649977179
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1649977179
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1649977179
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 1649977179
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_457
timestamp 1649977179
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1649977179
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1649977179
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1649977179
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_489
timestamp 1649977179
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_501
timestamp 1649977179
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_513
timestamp 1649977179
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_525
timestamp 1649977179
transform 1 0 49404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_531
timestamp 1649977179
transform 1 0 49956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_533
timestamp 1649977179
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_545
timestamp 1649977179
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_557
timestamp 1649977179
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_569
timestamp 1649977179
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_581
timestamp 1649977179
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_587
timestamp 1649977179
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_589
timestamp 1649977179
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_601
timestamp 1649977179
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_613
timestamp 1649977179
transform 1 0 57500 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_625
timestamp 1649977179
transform 1 0 58604 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_637
timestamp 1649977179
transform 1 0 59708 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_643
timestamp 1649977179
transform 1 0 60260 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_645
timestamp 1649977179
transform 1 0 60444 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_657
timestamp 1649977179
transform 1 0 61548 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_669
timestamp 1649977179
transform 1 0 62652 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_681
timestamp 1649977179
transform 1 0 63756 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_693
timestamp 1649977179
transform 1 0 64860 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_699
timestamp 1649977179
transform 1 0 65412 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_701
timestamp 1649977179
transform 1 0 65596 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_713
timestamp 1649977179
transform 1 0 66700 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_725
timestamp 1649977179
transform 1 0 67804 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_729
timestamp 1649977179
transform 1 0 68172 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1649977179
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1649977179
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1649977179
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1649977179
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1649977179
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1649977179
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1649977179
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1649977179
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1649977179
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1649977179
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1649977179
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1649977179
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1649977179
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1649977179
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1649977179
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1649977179
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1649977179
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1649977179
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1649977179
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1649977179
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1649977179
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1649977179
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1649977179
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1649977179
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1649977179
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1649977179
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_249
timestamp 1649977179
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_261
timestamp 1649977179
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_273
timestamp 1649977179
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1649977179
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_281
timestamp 1649977179
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_293
timestamp 1649977179
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_305
timestamp 1649977179
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_317
timestamp 1649977179
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1649977179
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1649977179
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_337
timestamp 1649977179
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_349
timestamp 1649977179
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_361
timestamp 1649977179
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_373
timestamp 1649977179
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_385
timestamp 1649977179
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1649977179
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_393
timestamp 1649977179
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_405
timestamp 1649977179
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_417
timestamp 1649977179
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_429
timestamp 1649977179
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_441
timestamp 1649977179
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1649977179
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_449
timestamp 1649977179
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_461
timestamp 1649977179
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_473
timestamp 1649977179
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_485
timestamp 1649977179
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_497
timestamp 1649977179
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1649977179
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_505
timestamp 1649977179
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_517
timestamp 1649977179
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_529
timestamp 1649977179
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_541
timestamp 1649977179
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_553
timestamp 1649977179
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_559
timestamp 1649977179
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_561
timestamp 1649977179
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_573
timestamp 1649977179
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_585
timestamp 1649977179
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_597
timestamp 1649977179
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_609
timestamp 1649977179
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_615
timestamp 1649977179
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_617
timestamp 1649977179
transform 1 0 57868 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_629
timestamp 1649977179
transform 1 0 58972 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_641
timestamp 1649977179
transform 1 0 60076 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_653
timestamp 1649977179
transform 1 0 61180 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_665
timestamp 1649977179
transform 1 0 62284 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_671
timestamp 1649977179
transform 1 0 62836 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_673
timestamp 1649977179
transform 1 0 63020 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_685
timestamp 1649977179
transform 1 0 64124 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_697
timestamp 1649977179
transform 1 0 65228 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_709
timestamp 1649977179
transform 1 0 66332 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_721
timestamp 1649977179
transform 1 0 67436 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_727
timestamp 1649977179
transform 1 0 67988 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_729
timestamp 1649977179
transform 1 0 68172 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1649977179
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1649977179
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1649977179
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1649977179
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1649977179
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1649977179
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1649977179
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1649977179
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1649977179
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1649977179
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1649977179
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1649977179
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1649977179
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1649977179
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1649977179
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1649977179
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1649977179
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1649977179
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1649977179
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1649977179
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1649977179
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1649977179
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1649977179
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1649977179
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1649977179
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1649977179
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1649977179
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_253
timestamp 1649977179
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_265
timestamp 1649977179
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_277
timestamp 1649977179
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_289
timestamp 1649977179
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1649977179
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1649977179
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_309
timestamp 1649977179
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_321
timestamp 1649977179
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_333
timestamp 1649977179
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_345
timestamp 1649977179
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_357
timestamp 1649977179
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1649977179
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_365
timestamp 1649977179
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_377
timestamp 1649977179
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_389
timestamp 1649977179
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_401
timestamp 1649977179
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_413
timestamp 1649977179
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1649977179
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1649977179
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1649977179
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_445
timestamp 1649977179
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_457
timestamp 1649977179
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1649977179
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1649977179
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_477
timestamp 1649977179
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_489
timestamp 1649977179
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_501
timestamp 1649977179
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_513
timestamp 1649977179
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_525
timestamp 1649977179
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_531
timestamp 1649977179
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_533
timestamp 1649977179
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_545
timestamp 1649977179
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_557
timestamp 1649977179
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_569
timestamp 1649977179
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_581
timestamp 1649977179
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_587
timestamp 1649977179
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_589
timestamp 1649977179
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_601
timestamp 1649977179
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_613
timestamp 1649977179
transform 1 0 57500 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_625
timestamp 1649977179
transform 1 0 58604 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_637
timestamp 1649977179
transform 1 0 59708 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_643
timestamp 1649977179
transform 1 0 60260 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_645
timestamp 1649977179
transform 1 0 60444 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_657
timestamp 1649977179
transform 1 0 61548 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_669
timestamp 1649977179
transform 1 0 62652 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_681
timestamp 1649977179
transform 1 0 63756 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_693
timestamp 1649977179
transform 1 0 64860 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_699
timestamp 1649977179
transform 1 0 65412 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_701
timestamp 1649977179
transform 1 0 65596 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_713
timestamp 1649977179
transform 1 0 66700 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_725
timestamp 1649977179
transform 1 0 67804 0 1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1649977179
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1649977179
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1649977179
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1649977179
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1649977179
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1649977179
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1649977179
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1649977179
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1649977179
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1649977179
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1649977179
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1649977179
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1649977179
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1649977179
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1649977179
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1649977179
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1649977179
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1649977179
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1649977179
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1649977179
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1649977179
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1649977179
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1649977179
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1649977179
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1649977179
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1649977179
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1649977179
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_261
timestamp 1649977179
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1649977179
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1649977179
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_281
timestamp 1649977179
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_293
timestamp 1649977179
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_305
timestamp 1649977179
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_317
timestamp 1649977179
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 1649977179
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1649977179
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_337
timestamp 1649977179
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_349
timestamp 1649977179
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_361
timestamp 1649977179
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_373
timestamp 1649977179
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1649977179
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1649977179
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_393
timestamp 1649977179
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_405
timestamp 1649977179
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_417
timestamp 1649977179
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_429
timestamp 1649977179
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1649977179
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1649977179
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_449
timestamp 1649977179
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_461
timestamp 1649977179
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_473
timestamp 1649977179
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_485
timestamp 1649977179
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1649977179
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1649977179
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1649977179
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_517
timestamp 1649977179
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_529
timestamp 1649977179
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_541
timestamp 1649977179
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_553
timestamp 1649977179
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_559
timestamp 1649977179
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_561
timestamp 1649977179
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_573
timestamp 1649977179
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_585
timestamp 1649977179
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_597
timestamp 1649977179
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_609
timestamp 1649977179
transform 1 0 57132 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_615
timestamp 1649977179
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_617
timestamp 1649977179
transform 1 0 57868 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_629
timestamp 1649977179
transform 1 0 58972 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_641
timestamp 1649977179
transform 1 0 60076 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_653
timestamp 1649977179
transform 1 0 61180 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_665
timestamp 1649977179
transform 1 0 62284 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_671
timestamp 1649977179
transform 1 0 62836 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_673
timestamp 1649977179
transform 1 0 63020 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_685
timestamp 1649977179
transform 1 0 64124 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_697
timestamp 1649977179
transform 1 0 65228 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_709
timestamp 1649977179
transform 1 0 66332 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_724
timestamp 1649977179
transform 1 0 67712 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_729
timestamp 1649977179
transform 1 0 68172 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1649977179
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1649977179
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1649977179
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1649977179
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1649977179
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1649977179
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1649977179
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1649977179
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1649977179
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1649977179
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1649977179
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1649977179
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1649977179
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1649977179
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1649977179
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1649977179
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1649977179
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1649977179
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1649977179
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1649977179
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1649977179
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1649977179
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1649977179
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1649977179
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1649977179
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1649977179
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1649977179
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_253
timestamp 1649977179
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_265
timestamp 1649977179
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_277
timestamp 1649977179
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_289
timestamp 1649977179
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1649977179
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1649977179
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_309
timestamp 1649977179
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_321
timestamp 1649977179
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_333
timestamp 1649977179
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_345
timestamp 1649977179
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_357
timestamp 1649977179
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1649977179
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_365
timestamp 1649977179
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_377
timestamp 1649977179
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_389
timestamp 1649977179
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_401
timestamp 1649977179
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 1649977179
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1649977179
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1649977179
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1649977179
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1649977179
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1649977179
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1649977179
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1649977179
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1649977179
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1649977179
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1649977179
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_513
timestamp 1649977179
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_525
timestamp 1649977179
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_531
timestamp 1649977179
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_533
timestamp 1649977179
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_545
timestamp 1649977179
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_557
timestamp 1649977179
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_569
timestamp 1649977179
transform 1 0 53452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_581
timestamp 1649977179
transform 1 0 54556 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_587
timestamp 1649977179
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_589
timestamp 1649977179
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_601
timestamp 1649977179
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_613
timestamp 1649977179
transform 1 0 57500 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_625
timestamp 1649977179
transform 1 0 58604 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_637
timestamp 1649977179
transform 1 0 59708 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_643
timestamp 1649977179
transform 1 0 60260 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_645
timestamp 1649977179
transform 1 0 60444 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_657
timestamp 1649977179
transform 1 0 61548 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_669
timestamp 1649977179
transform 1 0 62652 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_681
timestamp 1649977179
transform 1 0 63756 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_693
timestamp 1649977179
transform 1 0 64860 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_699
timestamp 1649977179
transform 1 0 65412 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_701
timestamp 1649977179
transform 1 0 65596 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_713
timestamp 1649977179
transform 1 0 66700 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_725
timestamp 1649977179
transform 1 0 67804 0 1 48960
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1649977179
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1649977179
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1649977179
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1649977179
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1649977179
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1649977179
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1649977179
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1649977179
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1649977179
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1649977179
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1649977179
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1649977179
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1649977179
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1649977179
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1649977179
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1649977179
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1649977179
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1649977179
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1649977179
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1649977179
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1649977179
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1649977179
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1649977179
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1649977179
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1649977179
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1649977179
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1649977179
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_261
timestamp 1649977179
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_273
timestamp 1649977179
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1649977179
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_281
timestamp 1649977179
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_293
timestamp 1649977179
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_305
timestamp 1649977179
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_317
timestamp 1649977179
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1649977179
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1649977179
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_337
timestamp 1649977179
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_349
timestamp 1649977179
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_361
timestamp 1649977179
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_373
timestamp 1649977179
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1649977179
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1649977179
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1649977179
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1649977179
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1649977179
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1649977179
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1649977179
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1649977179
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_449
timestamp 1649977179
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_461
timestamp 1649977179
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_473
timestamp 1649977179
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_485
timestamp 1649977179
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1649977179
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1649977179
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1649977179
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_517
timestamp 1649977179
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_529
timestamp 1649977179
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_541
timestamp 1649977179
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_553
timestamp 1649977179
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_559
timestamp 1649977179
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_561
timestamp 1649977179
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_573
timestamp 1649977179
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_585
timestamp 1649977179
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_597
timestamp 1649977179
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_609
timestamp 1649977179
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_615
timestamp 1649977179
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_617
timestamp 1649977179
transform 1 0 57868 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_629
timestamp 1649977179
transform 1 0 58972 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_641
timestamp 1649977179
transform 1 0 60076 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_653
timestamp 1649977179
transform 1 0 61180 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_665
timestamp 1649977179
transform 1 0 62284 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_671
timestamp 1649977179
transform 1 0 62836 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_673
timestamp 1649977179
transform 1 0 63020 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_685
timestamp 1649977179
transform 1 0 64124 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_697
timestamp 1649977179
transform 1 0 65228 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_709
timestamp 1649977179
transform 1 0 66332 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_724
timestamp 1649977179
transform 1 0 67712 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_729
timestamp 1649977179
transform 1 0 68172 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1649977179
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1649977179
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1649977179
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1649977179
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1649977179
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1649977179
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1649977179
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1649977179
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1649977179
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1649977179
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1649977179
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1649977179
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1649977179
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1649977179
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1649977179
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1649977179
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1649977179
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1649977179
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1649977179
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1649977179
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1649977179
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1649977179
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1649977179
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1649977179
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1649977179
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1649977179
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1649977179
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1649977179
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_265
timestamp 1649977179
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_277
timestamp 1649977179
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_289
timestamp 1649977179
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 1649977179
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1649977179
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_309
timestamp 1649977179
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_321
timestamp 1649977179
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_333
timestamp 1649977179
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_345
timestamp 1649977179
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1649977179
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1649977179
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_365
timestamp 1649977179
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_377
timestamp 1649977179
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_389
timestamp 1649977179
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_401
timestamp 1649977179
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1649977179
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1649977179
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1649977179
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1649977179
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1649977179
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1649977179
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1649977179
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1649977179
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_477
timestamp 1649977179
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_489
timestamp 1649977179
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_501
timestamp 1649977179
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_513
timestamp 1649977179
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_525
timestamp 1649977179
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_531
timestamp 1649977179
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_533
timestamp 1649977179
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_545
timestamp 1649977179
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_557
timestamp 1649977179
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_569
timestamp 1649977179
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_581
timestamp 1649977179
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_587
timestamp 1649977179
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_589
timestamp 1649977179
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_601
timestamp 1649977179
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_613
timestamp 1649977179
transform 1 0 57500 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_625
timestamp 1649977179
transform 1 0 58604 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_637
timestamp 1649977179
transform 1 0 59708 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_643
timestamp 1649977179
transform 1 0 60260 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_645
timestamp 1649977179
transform 1 0 60444 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_657
timestamp 1649977179
transform 1 0 61548 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_669
timestamp 1649977179
transform 1 0 62652 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_681
timestamp 1649977179
transform 1 0 63756 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_693
timestamp 1649977179
transform 1 0 64860 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_699
timestamp 1649977179
transform 1 0 65412 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_701
timestamp 1649977179
transform 1 0 65596 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_713
timestamp 1649977179
transform 1 0 66700 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_725
timestamp 1649977179
transform 1 0 67804 0 1 50048
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1649977179
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1649977179
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1649977179
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1649977179
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1649977179
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1649977179
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1649977179
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1649977179
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1649977179
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1649977179
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1649977179
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1649977179
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1649977179
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1649977179
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1649977179
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1649977179
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1649977179
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1649977179
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1649977179
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1649977179
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1649977179
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1649977179
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1649977179
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1649977179
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1649977179
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1649977179
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_249
timestamp 1649977179
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_261
timestamp 1649977179
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_273
timestamp 1649977179
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1649977179
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_281
timestamp 1649977179
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_293
timestamp 1649977179
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_305
timestamp 1649977179
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_317
timestamp 1649977179
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1649977179
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1649977179
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_337
timestamp 1649977179
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_349
timestamp 1649977179
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_361
timestamp 1649977179
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_373
timestamp 1649977179
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1649977179
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1649977179
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_393
timestamp 1649977179
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_405
timestamp 1649977179
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_417
timestamp 1649977179
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_429
timestamp 1649977179
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1649977179
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1649977179
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1649977179
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1649977179
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_473
timestamp 1649977179
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_485
timestamp 1649977179
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1649977179
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1649977179
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_505
timestamp 1649977179
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_517
timestamp 1649977179
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_529
timestamp 1649977179
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_541
timestamp 1649977179
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_553
timestamp 1649977179
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_559
timestamp 1649977179
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_561
timestamp 1649977179
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_573
timestamp 1649977179
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_585
timestamp 1649977179
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_597
timestamp 1649977179
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_609
timestamp 1649977179
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_615
timestamp 1649977179
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_617
timestamp 1649977179
transform 1 0 57868 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_629
timestamp 1649977179
transform 1 0 58972 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_641
timestamp 1649977179
transform 1 0 60076 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_653
timestamp 1649977179
transform 1 0 61180 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_665
timestamp 1649977179
transform 1 0 62284 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_671
timestamp 1649977179
transform 1 0 62836 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_673
timestamp 1649977179
transform 1 0 63020 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_685
timestamp 1649977179
transform 1 0 64124 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_697
timestamp 1649977179
transform 1 0 65228 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_709
timestamp 1649977179
transform 1 0 66332 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_721
timestamp 1649977179
transform 1 0 67436 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_727
timestamp 1649977179
transform 1 0 67988 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_729
timestamp 1649977179
transform 1 0 68172 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1649977179
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1649977179
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1649977179
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1649977179
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1649977179
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1649977179
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1649977179
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1649977179
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1649977179
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1649977179
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1649977179
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1649977179
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1649977179
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1649977179
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1649977179
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1649977179
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1649977179
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1649977179
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1649977179
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1649977179
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1649977179
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1649977179
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1649977179
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1649977179
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1649977179
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1649977179
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1649977179
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_253
timestamp 1649977179
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_265
timestamp 1649977179
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_277
timestamp 1649977179
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_289
timestamp 1649977179
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_301
timestamp 1649977179
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1649977179
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_309
timestamp 1649977179
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_321
timestamp 1649977179
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_333
timestamp 1649977179
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_345
timestamp 1649977179
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1649977179
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1649977179
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_365
timestamp 1649977179
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_377
timestamp 1649977179
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_389
timestamp 1649977179
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_401
timestamp 1649977179
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1649977179
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1649977179
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1649977179
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1649977179
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_445
timestamp 1649977179
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_457
timestamp 1649977179
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1649977179
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1649977179
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_477
timestamp 1649977179
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_489
timestamp 1649977179
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_501
timestamp 1649977179
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_513
timestamp 1649977179
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_525
timestamp 1649977179
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_531
timestamp 1649977179
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_533
timestamp 1649977179
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_545
timestamp 1649977179
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_557
timestamp 1649977179
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_569
timestamp 1649977179
transform 1 0 53452 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_581
timestamp 1649977179
transform 1 0 54556 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_587
timestamp 1649977179
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_589
timestamp 1649977179
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_601
timestamp 1649977179
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_613
timestamp 1649977179
transform 1 0 57500 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_625
timestamp 1649977179
transform 1 0 58604 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_637
timestamp 1649977179
transform 1 0 59708 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_643
timestamp 1649977179
transform 1 0 60260 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_645
timestamp 1649977179
transform 1 0 60444 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_657
timestamp 1649977179
transform 1 0 61548 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_669
timestamp 1649977179
transform 1 0 62652 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_681
timestamp 1649977179
transform 1 0 63756 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_693
timestamp 1649977179
transform 1 0 64860 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_699
timestamp 1649977179
transform 1 0 65412 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_701
timestamp 1649977179
transform 1 0 65596 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_713
timestamp 1649977179
transform 1 0 66700 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_725
timestamp 1649977179
transform 1 0 67804 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_729
timestamp 1649977179
transform 1 0 68172 0 1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1649977179
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1649977179
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1649977179
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1649977179
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1649977179
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1649977179
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1649977179
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1649977179
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_81
timestamp 1649977179
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_93
timestamp 1649977179
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1649977179
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1649977179
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1649977179
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1649977179
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1649977179
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1649977179
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1649977179
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1649977179
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1649977179
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1649977179
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1649977179
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1649977179
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1649977179
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1649977179
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1649977179
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1649977179
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1649977179
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_261
timestamp 1649977179
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1649977179
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1649977179
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_281
timestamp 1649977179
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_293
timestamp 1649977179
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_305
timestamp 1649977179
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_317
timestamp 1649977179
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1649977179
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1649977179
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_337
timestamp 1649977179
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_349
timestamp 1649977179
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1649977179
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1649977179
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1649977179
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1649977179
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_393
timestamp 1649977179
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_405
timestamp 1649977179
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_417
timestamp 1649977179
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_429
timestamp 1649977179
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1649977179
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1649977179
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1649977179
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1649977179
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1649977179
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_485
timestamp 1649977179
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1649977179
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1649977179
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_505
timestamp 1649977179
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_517
timestamp 1649977179
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_529
timestamp 1649977179
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_541
timestamp 1649977179
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_553
timestamp 1649977179
transform 1 0 51980 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_559
timestamp 1649977179
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_561
timestamp 1649977179
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_573
timestamp 1649977179
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_585
timestamp 1649977179
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_597
timestamp 1649977179
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_609
timestamp 1649977179
transform 1 0 57132 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_615
timestamp 1649977179
transform 1 0 57684 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_617
timestamp 1649977179
transform 1 0 57868 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_629
timestamp 1649977179
transform 1 0 58972 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_641
timestamp 1649977179
transform 1 0 60076 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_653
timestamp 1649977179
transform 1 0 61180 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_665
timestamp 1649977179
transform 1 0 62284 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_671
timestamp 1649977179
transform 1 0 62836 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_673
timestamp 1649977179
transform 1 0 63020 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_685
timestamp 1649977179
transform 1 0 64124 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_697
timestamp 1649977179
transform 1 0 65228 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_709
timestamp 1649977179
transform 1 0 66332 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_721
timestamp 1649977179
transform 1 0 67436 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_727
timestamp 1649977179
transform 1 0 67988 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_729
timestamp 1649977179
transform 1 0 68172 0 -1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1649977179
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1649977179
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1649977179
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1649977179
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1649977179
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1649977179
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_65
timestamp 1649977179
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1649977179
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1649977179
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1649977179
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1649977179
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1649977179
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1649977179
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1649977179
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1649977179
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1649977179
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1649977179
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1649977179
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1649977179
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1649977179
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1649977179
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1649977179
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1649977179
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1649977179
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1649977179
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1649977179
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1649977179
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_253
timestamp 1649977179
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_265
timestamp 1649977179
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_277
timestamp 1649977179
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_289
timestamp 1649977179
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_301
timestamp 1649977179
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_307
timestamp 1649977179
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_309
timestamp 1649977179
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_321
timestamp 1649977179
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_333
timestamp 1649977179
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_345
timestamp 1649977179
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1649977179
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1649977179
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_365
timestamp 1649977179
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_377
timestamp 1649977179
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_389
timestamp 1649977179
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_401
timestamp 1649977179
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1649977179
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1649977179
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1649977179
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1649977179
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_445
timestamp 1649977179
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_457
timestamp 1649977179
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 1649977179
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1649977179
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_477
timestamp 1649977179
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_489
timestamp 1649977179
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_501
timestamp 1649977179
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_513
timestamp 1649977179
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_525
timestamp 1649977179
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_531
timestamp 1649977179
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_533
timestamp 1649977179
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_545
timestamp 1649977179
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_557
timestamp 1649977179
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_569
timestamp 1649977179
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_581
timestamp 1649977179
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_587
timestamp 1649977179
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_589
timestamp 1649977179
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_601
timestamp 1649977179
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_613
timestamp 1649977179
transform 1 0 57500 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_625
timestamp 1649977179
transform 1 0 58604 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_637
timestamp 1649977179
transform 1 0 59708 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_643
timestamp 1649977179
transform 1 0 60260 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_645
timestamp 1649977179
transform 1 0 60444 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_657
timestamp 1649977179
transform 1 0 61548 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_669
timestamp 1649977179
transform 1 0 62652 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_681
timestamp 1649977179
transform 1 0 63756 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_693
timestamp 1649977179
transform 1 0 64860 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_699
timestamp 1649977179
transform 1 0 65412 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_701
timestamp 1649977179
transform 1 0 65596 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_713
timestamp 1649977179
transform 1 0 66700 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_725
timestamp 1649977179
transform 1 0 67804 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_729
timestamp 1649977179
transform 1 0 68172 0 1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1649977179
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1649977179
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1649977179
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_39
timestamp 1649977179
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_51
timestamp 1649977179
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1649977179
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1649977179
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_69
timestamp 1649977179
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_81
timestamp 1649977179
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_93
timestamp 1649977179
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1649977179
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1649977179
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1649977179
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1649977179
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1649977179
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1649977179
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1649977179
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1649977179
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1649977179
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1649977179
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1649977179
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1649977179
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1649977179
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1649977179
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1649977179
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_237
timestamp 1649977179
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_249
timestamp 1649977179
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_261
timestamp 1649977179
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_273
timestamp 1649977179
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 1649977179
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_281
timestamp 1649977179
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_293
timestamp 1649977179
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_305
timestamp 1649977179
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_317
timestamp 1649977179
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_329
timestamp 1649977179
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1649977179
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_337
timestamp 1649977179
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_349
timestamp 1649977179
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_361
timestamp 1649977179
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_373
timestamp 1649977179
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1649977179
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1649977179
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_393
timestamp 1649977179
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_405
timestamp 1649977179
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_417
timestamp 1649977179
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_429
timestamp 1649977179
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_441
timestamp 1649977179
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1649977179
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_449
timestamp 1649977179
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_461
timestamp 1649977179
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_473
timestamp 1649977179
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_485
timestamp 1649977179
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 1649977179
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1649977179
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_505
timestamp 1649977179
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_517
timestamp 1649977179
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_529
timestamp 1649977179
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_541
timestamp 1649977179
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_553
timestamp 1649977179
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_559
timestamp 1649977179
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_561
timestamp 1649977179
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_573
timestamp 1649977179
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_585
timestamp 1649977179
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_597
timestamp 1649977179
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_609
timestamp 1649977179
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_615
timestamp 1649977179
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_617
timestamp 1649977179
transform 1 0 57868 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_629
timestamp 1649977179
transform 1 0 58972 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_641
timestamp 1649977179
transform 1 0 60076 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_653
timestamp 1649977179
transform 1 0 61180 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_665
timestamp 1649977179
transform 1 0 62284 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_671
timestamp 1649977179
transform 1 0 62836 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_673
timestamp 1649977179
transform 1 0 63020 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_685
timestamp 1649977179
transform 1 0 64124 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_697
timestamp 1649977179
transform 1 0 65228 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_709
timestamp 1649977179
transform 1 0 66332 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_721
timestamp 1649977179
transform 1 0 67436 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_727
timestamp 1649977179
transform 1 0 67988 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_729
timestamp 1649977179
transform 1 0 68172 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_3
timestamp 1649977179
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_15
timestamp 1649977179
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1649977179
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1649977179
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1649977179
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1649977179
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_65
timestamp 1649977179
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1649977179
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1649977179
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1649977179
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_97
timestamp 1649977179
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_109
timestamp 1649977179
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1649977179
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1649977179
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1649977179
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1649977179
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1649977179
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1649977179
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1649977179
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1649977179
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1649977179
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1649977179
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1649977179
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_221
timestamp 1649977179
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_233
timestamp 1649977179
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_245
timestamp 1649977179
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1649977179
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_253
timestamp 1649977179
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_265
timestamp 1649977179
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_277
timestamp 1649977179
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_289
timestamp 1649977179
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_301
timestamp 1649977179
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_307
timestamp 1649977179
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_309
timestamp 1649977179
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_321
timestamp 1649977179
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_333
timestamp 1649977179
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_345
timestamp 1649977179
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_357
timestamp 1649977179
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_363
timestamp 1649977179
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_365
timestamp 1649977179
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_377
timestamp 1649977179
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_389
timestamp 1649977179
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_401
timestamp 1649977179
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_413
timestamp 1649977179
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_419
timestamp 1649977179
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_421
timestamp 1649977179
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_433
timestamp 1649977179
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_445
timestamp 1649977179
transform 1 0 42044 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_457
timestamp 1649977179
transform 1 0 43148 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_469
timestamp 1649977179
transform 1 0 44252 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_475
timestamp 1649977179
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_477
timestamp 1649977179
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_489
timestamp 1649977179
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_501
timestamp 1649977179
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_513
timestamp 1649977179
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_525
timestamp 1649977179
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_531
timestamp 1649977179
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_533
timestamp 1649977179
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_545
timestamp 1649977179
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_557
timestamp 1649977179
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_569
timestamp 1649977179
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_581
timestamp 1649977179
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_587
timestamp 1649977179
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_589
timestamp 1649977179
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_601
timestamp 1649977179
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_613
timestamp 1649977179
transform 1 0 57500 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_625
timestamp 1649977179
transform 1 0 58604 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_637
timestamp 1649977179
transform 1 0 59708 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_643
timestamp 1649977179
transform 1 0 60260 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_645
timestamp 1649977179
transform 1 0 60444 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_657
timestamp 1649977179
transform 1 0 61548 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_669
timestamp 1649977179
transform 1 0 62652 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_681
timestamp 1649977179
transform 1 0 63756 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_693
timestamp 1649977179
transform 1 0 64860 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_699
timestamp 1649977179
transform 1 0 65412 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_701
timestamp 1649977179
transform 1 0 65596 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_713
timestamp 1649977179
transform 1 0 66700 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_725
timestamp 1649977179
transform 1 0 67804 0 1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_95_3
timestamp 1649977179
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_15
timestamp 1649977179
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_27
timestamp 1649977179
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_39
timestamp 1649977179
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_51
timestamp 1649977179
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1649977179
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_57
timestamp 1649977179
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_69
timestamp 1649977179
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_81
timestamp 1649977179
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_93
timestamp 1649977179
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_105
timestamp 1649977179
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1649977179
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_113
timestamp 1649977179
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_125
timestamp 1649977179
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_137
timestamp 1649977179
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_149
timestamp 1649977179
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_161
timestamp 1649977179
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1649977179
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_169
timestamp 1649977179
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_181
timestamp 1649977179
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_193
timestamp 1649977179
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_205
timestamp 1649977179
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_217
timestamp 1649977179
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1649977179
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_225
timestamp 1649977179
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_237
timestamp 1649977179
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_249
timestamp 1649977179
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_261
timestamp 1649977179
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_273
timestamp 1649977179
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_279
timestamp 1649977179
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_281
timestamp 1649977179
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_293
timestamp 1649977179
transform 1 0 28060 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_305
timestamp 1649977179
transform 1 0 29164 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_317
timestamp 1649977179
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_329
timestamp 1649977179
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_335
timestamp 1649977179
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_337
timestamp 1649977179
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_349
timestamp 1649977179
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_361
timestamp 1649977179
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_373
timestamp 1649977179
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_385
timestamp 1649977179
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 1649977179
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_393
timestamp 1649977179
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_405
timestamp 1649977179
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_417
timestamp 1649977179
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_429
timestamp 1649977179
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_441
timestamp 1649977179
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_447
timestamp 1649977179
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_449
timestamp 1649977179
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_461
timestamp 1649977179
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_473
timestamp 1649977179
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_485
timestamp 1649977179
transform 1 0 45724 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_497
timestamp 1649977179
transform 1 0 46828 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_503
timestamp 1649977179
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_505
timestamp 1649977179
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_517
timestamp 1649977179
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_529
timestamp 1649977179
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_541
timestamp 1649977179
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_553
timestamp 1649977179
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_559
timestamp 1649977179
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_561
timestamp 1649977179
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_573
timestamp 1649977179
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_585
timestamp 1649977179
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_597
timestamp 1649977179
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_609
timestamp 1649977179
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 1649977179
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_617
timestamp 1649977179
transform 1 0 57868 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_629
timestamp 1649977179
transform 1 0 58972 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_641
timestamp 1649977179
transform 1 0 60076 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_653
timestamp 1649977179
transform 1 0 61180 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_665
timestamp 1649977179
transform 1 0 62284 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_671
timestamp 1649977179
transform 1 0 62836 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_673
timestamp 1649977179
transform 1 0 63020 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_685
timestamp 1649977179
transform 1 0 64124 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_697
timestamp 1649977179
transform 1 0 65228 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_709
timestamp 1649977179
transform 1 0 66332 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_724
timestamp 1649977179
transform 1 0 67712 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_729
timestamp 1649977179
transform 1 0 68172 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_96_3
timestamp 1649977179
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_15
timestamp 1649977179
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1649977179
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1649977179
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1649977179
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_53
timestamp 1649977179
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_65
timestamp 1649977179
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1649977179
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1649977179
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_85
timestamp 1649977179
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_97
timestamp 1649977179
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_109
timestamp 1649977179
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_121
timestamp 1649977179
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 1649977179
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1649977179
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_141
timestamp 1649977179
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_153
timestamp 1649977179
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_165
timestamp 1649977179
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_177
timestamp 1649977179
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_189
timestamp 1649977179
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 1649977179
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_197
timestamp 1649977179
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_209
timestamp 1649977179
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_221
timestamp 1649977179
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_233
timestamp 1649977179
transform 1 0 22540 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_245
timestamp 1649977179
transform 1 0 23644 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_251
timestamp 1649977179
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_253
timestamp 1649977179
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_265
timestamp 1649977179
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_277
timestamp 1649977179
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_289
timestamp 1649977179
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_301
timestamp 1649977179
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_307
timestamp 1649977179
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_309
timestamp 1649977179
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_321
timestamp 1649977179
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_333
timestamp 1649977179
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_345
timestamp 1649977179
transform 1 0 32844 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_357
timestamp 1649977179
transform 1 0 33948 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_363
timestamp 1649977179
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_365
timestamp 1649977179
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_377
timestamp 1649977179
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_389
timestamp 1649977179
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_401
timestamp 1649977179
transform 1 0 37996 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_413
timestamp 1649977179
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_419
timestamp 1649977179
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_421
timestamp 1649977179
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_433
timestamp 1649977179
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_445
timestamp 1649977179
transform 1 0 42044 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_457
timestamp 1649977179
transform 1 0 43148 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_469
timestamp 1649977179
transform 1 0 44252 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_475
timestamp 1649977179
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_477
timestamp 1649977179
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_489
timestamp 1649977179
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_501
timestamp 1649977179
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_513
timestamp 1649977179
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_525
timestamp 1649977179
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_531
timestamp 1649977179
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_533
timestamp 1649977179
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_545
timestamp 1649977179
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_557
timestamp 1649977179
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_569
timestamp 1649977179
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_581
timestamp 1649977179
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_587
timestamp 1649977179
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_589
timestamp 1649977179
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_601
timestamp 1649977179
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_613
timestamp 1649977179
transform 1 0 57500 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_625
timestamp 1649977179
transform 1 0 58604 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_637
timestamp 1649977179
transform 1 0 59708 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_643
timestamp 1649977179
transform 1 0 60260 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_645
timestamp 1649977179
transform 1 0 60444 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_657
timestamp 1649977179
transform 1 0 61548 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_669
timestamp 1649977179
transform 1 0 62652 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_681
timestamp 1649977179
transform 1 0 63756 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_693
timestamp 1649977179
transform 1 0 64860 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_699
timestamp 1649977179
transform 1 0 65412 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_701
timestamp 1649977179
transform 1 0 65596 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_713
timestamp 1649977179
transform 1 0 66700 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_725
timestamp 1649977179
transform 1 0 67804 0 1 54400
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_97_3
timestamp 1649977179
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_15
timestamp 1649977179
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_27
timestamp 1649977179
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_39
timestamp 1649977179
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 1649977179
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1649977179
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_57
timestamp 1649977179
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_69
timestamp 1649977179
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_81
timestamp 1649977179
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_93
timestamp 1649977179
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_105
timestamp 1649977179
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 1649977179
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_113
timestamp 1649977179
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_125
timestamp 1649977179
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_137
timestamp 1649977179
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_149
timestamp 1649977179
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_161
timestamp 1649977179
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_167
timestamp 1649977179
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_169
timestamp 1649977179
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_181
timestamp 1649977179
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_193
timestamp 1649977179
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_205
timestamp 1649977179
transform 1 0 19964 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_217
timestamp 1649977179
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_223
timestamp 1649977179
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_225
timestamp 1649977179
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_237
timestamp 1649977179
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_249
timestamp 1649977179
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_261
timestamp 1649977179
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_273
timestamp 1649977179
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_279
timestamp 1649977179
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_281
timestamp 1649977179
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_293
timestamp 1649977179
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_305
timestamp 1649977179
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_317
timestamp 1649977179
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_329
timestamp 1649977179
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_335
timestamp 1649977179
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_337
timestamp 1649977179
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_349
timestamp 1649977179
transform 1 0 33212 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_361
timestamp 1649977179
transform 1 0 34316 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_373
timestamp 1649977179
transform 1 0 35420 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_385
timestamp 1649977179
transform 1 0 36524 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_391
timestamp 1649977179
transform 1 0 37076 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_393
timestamp 1649977179
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_405
timestamp 1649977179
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_417
timestamp 1649977179
transform 1 0 39468 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_429
timestamp 1649977179
transform 1 0 40572 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_441
timestamp 1649977179
transform 1 0 41676 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_447
timestamp 1649977179
transform 1 0 42228 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_449
timestamp 1649977179
transform 1 0 42412 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_461
timestamp 1649977179
transform 1 0 43516 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_473
timestamp 1649977179
transform 1 0 44620 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_485
timestamp 1649977179
transform 1 0 45724 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_497
timestamp 1649977179
transform 1 0 46828 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_503
timestamp 1649977179
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_505
timestamp 1649977179
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_517
timestamp 1649977179
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_529
timestamp 1649977179
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_541
timestamp 1649977179
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_553
timestamp 1649977179
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_559
timestamp 1649977179
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_561
timestamp 1649977179
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_573
timestamp 1649977179
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_585
timestamp 1649977179
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_597
timestamp 1649977179
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_609
timestamp 1649977179
transform 1 0 57132 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_615
timestamp 1649977179
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_617
timestamp 1649977179
transform 1 0 57868 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_629
timestamp 1649977179
transform 1 0 58972 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_641
timestamp 1649977179
transform 1 0 60076 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_653
timestamp 1649977179
transform 1 0 61180 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_665
timestamp 1649977179
transform 1 0 62284 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_671
timestamp 1649977179
transform 1 0 62836 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_673
timestamp 1649977179
transform 1 0 63020 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_685
timestamp 1649977179
transform 1 0 64124 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_697
timestamp 1649977179
transform 1 0 65228 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_709
timestamp 1649977179
transform 1 0 66332 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_724
timestamp 1649977179
transform 1 0 67712 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_729
timestamp 1649977179
transform 1 0 68172 0 -1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_98_3
timestamp 1649977179
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_15
timestamp 1649977179
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1649977179
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1649977179
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_41
timestamp 1649977179
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_53
timestamp 1649977179
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_65
timestamp 1649977179
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1649977179
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1649977179
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_85
timestamp 1649977179
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_97
timestamp 1649977179
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_109
timestamp 1649977179
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_121
timestamp 1649977179
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_133
timestamp 1649977179
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 1649977179
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_141
timestamp 1649977179
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_153
timestamp 1649977179
transform 1 0 15180 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_165
timestamp 1649977179
transform 1 0 16284 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_177
timestamp 1649977179
transform 1 0 17388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_189
timestamp 1649977179
transform 1 0 18492 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_195
timestamp 1649977179
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_197
timestamp 1649977179
transform 1 0 19228 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_209
timestamp 1649977179
transform 1 0 20332 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_221
timestamp 1649977179
transform 1 0 21436 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_233
timestamp 1649977179
transform 1 0 22540 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_245
timestamp 1649977179
transform 1 0 23644 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_251
timestamp 1649977179
transform 1 0 24196 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_253
timestamp 1649977179
transform 1 0 24380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_265
timestamp 1649977179
transform 1 0 25484 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_277
timestamp 1649977179
transform 1 0 26588 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_289
timestamp 1649977179
transform 1 0 27692 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_301
timestamp 1649977179
transform 1 0 28796 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_307
timestamp 1649977179
transform 1 0 29348 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_309
timestamp 1649977179
transform 1 0 29532 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_321
timestamp 1649977179
transform 1 0 30636 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_333
timestamp 1649977179
transform 1 0 31740 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_345
timestamp 1649977179
transform 1 0 32844 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_357
timestamp 1649977179
transform 1 0 33948 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_363
timestamp 1649977179
transform 1 0 34500 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_365
timestamp 1649977179
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_377
timestamp 1649977179
transform 1 0 35788 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_389
timestamp 1649977179
transform 1 0 36892 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_401
timestamp 1649977179
transform 1 0 37996 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_413
timestamp 1649977179
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_419
timestamp 1649977179
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_421
timestamp 1649977179
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_433
timestamp 1649977179
transform 1 0 40940 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_445
timestamp 1649977179
transform 1 0 42044 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_457
timestamp 1649977179
transform 1 0 43148 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_469
timestamp 1649977179
transform 1 0 44252 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_475
timestamp 1649977179
transform 1 0 44804 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_477
timestamp 1649977179
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_489
timestamp 1649977179
transform 1 0 46092 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_501
timestamp 1649977179
transform 1 0 47196 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_513
timestamp 1649977179
transform 1 0 48300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_525
timestamp 1649977179
transform 1 0 49404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_531
timestamp 1649977179
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_533
timestamp 1649977179
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_545
timestamp 1649977179
transform 1 0 51244 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_557
timestamp 1649977179
transform 1 0 52348 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_569
timestamp 1649977179
transform 1 0 53452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_581
timestamp 1649977179
transform 1 0 54556 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_587
timestamp 1649977179
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_589
timestamp 1649977179
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_601
timestamp 1649977179
transform 1 0 56396 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_613
timestamp 1649977179
transform 1 0 57500 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_625
timestamp 1649977179
transform 1 0 58604 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_637
timestamp 1649977179
transform 1 0 59708 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_643
timestamp 1649977179
transform 1 0 60260 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_645
timestamp 1649977179
transform 1 0 60444 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_657
timestamp 1649977179
transform 1 0 61548 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_669
timestamp 1649977179
transform 1 0 62652 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_681
timestamp 1649977179
transform 1 0 63756 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_693
timestamp 1649977179
transform 1 0 64860 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_699
timestamp 1649977179
transform 1 0 65412 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_701
timestamp 1649977179
transform 1 0 65596 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_713
timestamp 1649977179
transform 1 0 66700 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_725
timestamp 1649977179
transform 1 0 67804 0 1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_99_3
timestamp 1649977179
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_15
timestamp 1649977179
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_27
timestamp 1649977179
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_39
timestamp 1649977179
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 1649977179
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1649977179
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_57
timestamp 1649977179
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_69
timestamp 1649977179
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_81
timestamp 1649977179
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_93
timestamp 1649977179
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_105
timestamp 1649977179
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1649977179
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_113
timestamp 1649977179
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_125
timestamp 1649977179
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_137
timestamp 1649977179
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_149
timestamp 1649977179
transform 1 0 14812 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_161
timestamp 1649977179
transform 1 0 15916 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_167
timestamp 1649977179
transform 1 0 16468 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_169
timestamp 1649977179
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_181
timestamp 1649977179
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_193
timestamp 1649977179
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_205
timestamp 1649977179
transform 1 0 19964 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_217
timestamp 1649977179
transform 1 0 21068 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_223
timestamp 1649977179
transform 1 0 21620 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_225
timestamp 1649977179
transform 1 0 21804 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_237
timestamp 1649977179
transform 1 0 22908 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_249
timestamp 1649977179
transform 1 0 24012 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_261
timestamp 1649977179
transform 1 0 25116 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_273
timestamp 1649977179
transform 1 0 26220 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_279
timestamp 1649977179
transform 1 0 26772 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_281
timestamp 1649977179
transform 1 0 26956 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_293
timestamp 1649977179
transform 1 0 28060 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_305
timestamp 1649977179
transform 1 0 29164 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_317
timestamp 1649977179
transform 1 0 30268 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_329
timestamp 1649977179
transform 1 0 31372 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_335
timestamp 1649977179
transform 1 0 31924 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_337
timestamp 1649977179
transform 1 0 32108 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_349
timestamp 1649977179
transform 1 0 33212 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_361
timestamp 1649977179
transform 1 0 34316 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_373
timestamp 1649977179
transform 1 0 35420 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_385
timestamp 1649977179
transform 1 0 36524 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_391
timestamp 1649977179
transform 1 0 37076 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_393
timestamp 1649977179
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_405
timestamp 1649977179
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_417
timestamp 1649977179
transform 1 0 39468 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_429
timestamp 1649977179
transform 1 0 40572 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_441
timestamp 1649977179
transform 1 0 41676 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_447
timestamp 1649977179
transform 1 0 42228 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_449
timestamp 1649977179
transform 1 0 42412 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_461
timestamp 1649977179
transform 1 0 43516 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_473
timestamp 1649977179
transform 1 0 44620 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_485
timestamp 1649977179
transform 1 0 45724 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_497
timestamp 1649977179
transform 1 0 46828 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_503
timestamp 1649977179
transform 1 0 47380 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_505
timestamp 1649977179
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_517
timestamp 1649977179
transform 1 0 48668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_529
timestamp 1649977179
transform 1 0 49772 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_541
timestamp 1649977179
transform 1 0 50876 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_553
timestamp 1649977179
transform 1 0 51980 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_559
timestamp 1649977179
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_561
timestamp 1649977179
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_573
timestamp 1649977179
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_585
timestamp 1649977179
transform 1 0 54924 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_597
timestamp 1649977179
transform 1 0 56028 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_609
timestamp 1649977179
transform 1 0 57132 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_615
timestamp 1649977179
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_617
timestamp 1649977179
transform 1 0 57868 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_629
timestamp 1649977179
transform 1 0 58972 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_641
timestamp 1649977179
transform 1 0 60076 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_653
timestamp 1649977179
transform 1 0 61180 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_665
timestamp 1649977179
transform 1 0 62284 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_671
timestamp 1649977179
transform 1 0 62836 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_673
timestamp 1649977179
transform 1 0 63020 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_685
timestamp 1649977179
transform 1 0 64124 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_697
timestamp 1649977179
transform 1 0 65228 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_709
timestamp 1649977179
transform 1 0 66332 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_721
timestamp 1649977179
transform 1 0 67436 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_727
timestamp 1649977179
transform 1 0 67988 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_729
timestamp 1649977179
transform 1 0 68172 0 -1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_3
timestamp 1649977179
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_15
timestamp 1649977179
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1649977179
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_29
timestamp 1649977179
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_41
timestamp 1649977179
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_53
timestamp 1649977179
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_65
timestamp 1649977179
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 1649977179
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1649977179
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_85
timestamp 1649977179
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_97
timestamp 1649977179
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_109
timestamp 1649977179
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_121
timestamp 1649977179
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_133
timestamp 1649977179
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_139
timestamp 1649977179
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_141
timestamp 1649977179
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_153
timestamp 1649977179
transform 1 0 15180 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_165
timestamp 1649977179
transform 1 0 16284 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_177
timestamp 1649977179
transform 1 0 17388 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_189
timestamp 1649977179
transform 1 0 18492 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_195
timestamp 1649977179
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_197
timestamp 1649977179
transform 1 0 19228 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_209
timestamp 1649977179
transform 1 0 20332 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_221
timestamp 1649977179
transform 1 0 21436 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_233
timestamp 1649977179
transform 1 0 22540 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_245
timestamp 1649977179
transform 1 0 23644 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_251
timestamp 1649977179
transform 1 0 24196 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_253
timestamp 1649977179
transform 1 0 24380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_265
timestamp 1649977179
transform 1 0 25484 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_277
timestamp 1649977179
transform 1 0 26588 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_289
timestamp 1649977179
transform 1 0 27692 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_301
timestamp 1649977179
transform 1 0 28796 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_307
timestamp 1649977179
transform 1 0 29348 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_309
timestamp 1649977179
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_321
timestamp 1649977179
transform 1 0 30636 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_333
timestamp 1649977179
transform 1 0 31740 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_345
timestamp 1649977179
transform 1 0 32844 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_357
timestamp 1649977179
transform 1 0 33948 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_363
timestamp 1649977179
transform 1 0 34500 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_365
timestamp 1649977179
transform 1 0 34684 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_377
timestamp 1649977179
transform 1 0 35788 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_389
timestamp 1649977179
transform 1 0 36892 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_401
timestamp 1649977179
transform 1 0 37996 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_413
timestamp 1649977179
transform 1 0 39100 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_419
timestamp 1649977179
transform 1 0 39652 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_421
timestamp 1649977179
transform 1 0 39836 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_433
timestamp 1649977179
transform 1 0 40940 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_445
timestamp 1649977179
transform 1 0 42044 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_457
timestamp 1649977179
transform 1 0 43148 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_469
timestamp 1649977179
transform 1 0 44252 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_475
timestamp 1649977179
transform 1 0 44804 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_477
timestamp 1649977179
transform 1 0 44988 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_489
timestamp 1649977179
transform 1 0 46092 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_501
timestamp 1649977179
transform 1 0 47196 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_513
timestamp 1649977179
transform 1 0 48300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_525
timestamp 1649977179
transform 1 0 49404 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_531
timestamp 1649977179
transform 1 0 49956 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_533
timestamp 1649977179
transform 1 0 50140 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_545
timestamp 1649977179
transform 1 0 51244 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_557
timestamp 1649977179
transform 1 0 52348 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_569
timestamp 1649977179
transform 1 0 53452 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_581
timestamp 1649977179
transform 1 0 54556 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_587
timestamp 1649977179
transform 1 0 55108 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_589
timestamp 1649977179
transform 1 0 55292 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_601
timestamp 1649977179
transform 1 0 56396 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_613
timestamp 1649977179
transform 1 0 57500 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_625
timestamp 1649977179
transform 1 0 58604 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_637
timestamp 1649977179
transform 1 0 59708 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_643
timestamp 1649977179
transform 1 0 60260 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_645
timestamp 1649977179
transform 1 0 60444 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_657
timestamp 1649977179
transform 1 0 61548 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_669
timestamp 1649977179
transform 1 0 62652 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_681
timestamp 1649977179
transform 1 0 63756 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_693
timestamp 1649977179
transform 1 0 64860 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_699
timestamp 1649977179
transform 1 0 65412 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_701
timestamp 1649977179
transform 1 0 65596 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_713
timestamp 1649977179
transform 1 0 66700 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_725
timestamp 1649977179
transform 1 0 67804 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_729
timestamp 1649977179
transform 1 0 68172 0 1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_101_3
timestamp 1649977179
transform 1 0 1380 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_15
timestamp 1649977179
transform 1 0 2484 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_27
timestamp 1649977179
transform 1 0 3588 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_29
timestamp 1649977179
transform 1 0 3772 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_41
timestamp 1649977179
transform 1 0 4876 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_48
timestamp 1649977179
transform 1 0 5520 0 -1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_101_57
timestamp 1649977179
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_69
timestamp 1649977179
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_81
timestamp 1649977179
transform 1 0 8556 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_85
timestamp 1649977179
transform 1 0 8924 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_97
timestamp 1649977179
transform 1 0 10028 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_109
timestamp 1649977179
transform 1 0 11132 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_113
timestamp 1649977179
transform 1 0 11500 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_125
timestamp 1649977179
transform 1 0 12604 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_137
timestamp 1649977179
transform 1 0 13708 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_141
timestamp 1649977179
transform 1 0 14076 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_156
timestamp 1649977179
transform 1 0 15456 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_169
timestamp 1649977179
transform 1 0 16652 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_181
timestamp 1649977179
transform 1 0 17756 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_193
timestamp 1649977179
transform 1 0 18860 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_197
timestamp 1649977179
transform 1 0 19228 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_209
timestamp 1649977179
transform 1 0 20332 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_221
timestamp 1649977179
transform 1 0 21436 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_225
timestamp 1649977179
transform 1 0 21804 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_237
timestamp 1649977179
transform 1 0 22908 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_249
timestamp 1649977179
transform 1 0 24012 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_101_253
timestamp 1649977179
transform 1 0 24380 0 -1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_101_264
timestamp 1649977179
transform 1 0 25392 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_276
timestamp 1649977179
transform 1 0 26496 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_101_281
timestamp 1649977179
transform 1 0 26956 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_293
timestamp 1649977179
transform 1 0 28060 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_305
timestamp 1649977179
transform 1 0 29164 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_309
timestamp 1649977179
transform 1 0 29532 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_321
timestamp 1649977179
transform 1 0 30636 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_333
timestamp 1649977179
transform 1 0 31740 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_337
timestamp 1649977179
transform 1 0 32108 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_349
timestamp 1649977179
transform 1 0 33212 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_361
timestamp 1649977179
transform 1 0 34316 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_365
timestamp 1649977179
transform 1 0 34684 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_101_372
timestamp 1649977179
transform 1 0 35328 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_384
timestamp 1649977179
transform 1 0 36432 0 -1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_101_393
timestamp 1649977179
transform 1 0 37260 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_405
timestamp 1649977179
transform 1 0 38364 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_417
timestamp 1649977179
transform 1 0 39468 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_421
timestamp 1649977179
transform 1 0 39836 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_433
timestamp 1649977179
transform 1 0 40940 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_445
timestamp 1649977179
transform 1 0 42044 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_449
timestamp 1649977179
transform 1 0 42412 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_461
timestamp 1649977179
transform 1 0 43516 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_473
timestamp 1649977179
transform 1 0 44620 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_480
timestamp 1649977179
transform 1 0 45264 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_492
timestamp 1649977179
transform 1 0 46368 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_505
timestamp 1649977179
transform 1 0 47564 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_517
timestamp 1649977179
transform 1 0 48668 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_529
timestamp 1649977179
transform 1 0 49772 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_533
timestamp 1649977179
transform 1 0 50140 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_545
timestamp 1649977179
transform 1 0 51244 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_557
timestamp 1649977179
transform 1 0 52348 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_561
timestamp 1649977179
transform 1 0 52716 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_573
timestamp 1649977179
transform 1 0 53820 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_585
timestamp 1649977179
transform 1 0 54924 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_592
timestamp 1649977179
transform 1 0 55568 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_604
timestamp 1649977179
transform 1 0 56672 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_617
timestamp 1649977179
transform 1 0 57868 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_629
timestamp 1649977179
transform 1 0 58972 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_641
timestamp 1649977179
transform 1 0 60076 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_645
timestamp 1649977179
transform 1 0 60444 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_657
timestamp 1649977179
transform 1 0 61548 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_669
timestamp 1649977179
transform 1 0 62652 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_673
timestamp 1649977179
transform 1 0 63020 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_685
timestamp 1649977179
transform 1 0 64124 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_696
timestamp 1649977179
transform 1 0 65136 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_101_701
timestamp 1649977179
transform 1 0 65596 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_713
timestamp 1649977179
transform 1 0 66700 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_717
timestamp 1649977179
transform 1 0 67068 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_724
timestamp 1649977179
transform 1 0 67712 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_729
timestamp 1649977179
transform 1 0 68172 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 68816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 68816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 68816 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 68816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 68816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 68816 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 68816 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 68816 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 68816 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 68816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 68816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 68816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 68816 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 68816 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 68816 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 68816 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 68816 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 68816 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 68816 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 68816 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 68816 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 68816 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 68816 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 68816 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 68816 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 68816 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 68816 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 68816 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 68816 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 68816 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 68816 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 68816 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 68816 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 68816 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 68816 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 68816 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 68816 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 68816 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 68816 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 68816 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1649977179
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1649977179
transform -1 0 68816 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1649977179
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1649977179
transform -1 0 68816 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1649977179
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1649977179
transform -1 0 68816 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1649977179
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1649977179
transform -1 0 68816 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1649977179
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1649977179
transform -1 0 68816 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1649977179
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1649977179
transform -1 0 68816 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1649977179
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1649977179
transform -1 0 68816 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1649977179
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1649977179
transform -1 0 68816 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1649977179
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1649977179
transform -1 0 68816 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1649977179
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1649977179
transform -1 0 68816 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1649977179
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1649977179
transform -1 0 68816 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1649977179
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1649977179
transform -1 0 68816 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1649977179
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1649977179
transform -1 0 68816 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1649977179
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1649977179
transform -1 0 68816 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1649977179
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1649977179
transform -1 0 68816 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1649977179
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1649977179
transform -1 0 68816 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1649977179
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1649977179
transform -1 0 68816 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1649977179
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1649977179
transform -1 0 68816 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1649977179
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1649977179
transform -1 0 68816 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1649977179
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1649977179
transform -1 0 68816 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1649977179
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1649977179
transform -1 0 68816 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1649977179
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1649977179
transform -1 0 68816 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1649977179
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1649977179
transform -1 0 68816 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1649977179
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1649977179
transform -1 0 68816 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1649977179
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1649977179
transform -1 0 68816 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1649977179
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1649977179
transform -1 0 68816 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1649977179
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1649977179
transform -1 0 68816 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1649977179
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1649977179
transform -1 0 68816 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1649977179
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1649977179
transform -1 0 68816 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1649977179
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1649977179
transform -1 0 68816 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1649977179
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1649977179
transform -1 0 68816 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1649977179
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1649977179
transform -1 0 68816 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1649977179
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1649977179
transform -1 0 68816 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1649977179
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1649977179
transform -1 0 68816 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1649977179
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1649977179
transform -1 0 68816 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1649977179
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1649977179
transform -1 0 68816 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1649977179
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1649977179
transform -1 0 68816 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1649977179
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1649977179
transform -1 0 68816 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1649977179
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1649977179
transform -1 0 68816 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1649977179
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1649977179
transform -1 0 68816 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1649977179
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1649977179
transform -1 0 68816 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1649977179
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1649977179
transform -1 0 68816 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1649977179
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1649977179
transform -1 0 68816 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1649977179
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1649977179
transform -1 0 68816 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1649977179
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1649977179
transform -1 0 68816 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1649977179
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1649977179
transform -1 0 68816 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1649977179
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1649977179
transform -1 0 68816 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1649977179
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1649977179
transform -1 0 68816 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1649977179
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1649977179
transform -1 0 68816 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1649977179
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1649977179
transform -1 0 68816 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1649977179
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1649977179
transform -1 0 68816 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1649977179
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1649977179
transform -1 0 68816 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1649977179
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1649977179
transform -1 0 68816 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1649977179
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1649977179
transform -1 0 68816 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1649977179
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1649977179
transform -1 0 68816 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1649977179
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1649977179
transform -1 0 68816 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1649977179
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1649977179
transform -1 0 68816 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1649977179
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1649977179
transform -1 0 68816 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1649977179
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1649977179
transform -1 0 68816 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1649977179
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1649977179
transform -1 0 68816 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1649977179
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1649977179
transform -1 0 68816 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1649977179
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1649977179
transform -1 0 68816 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1649977179
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1649977179
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1649977179
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1649977179
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1649977179
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1649977179
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1649977179
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1649977179
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1649977179
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1649977179
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1649977179
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1649977179
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1649977179
transform 1 0 60352 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1649977179
transform 1 0 65504 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1649977179
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1649977179
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1649977179
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1649977179
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1649977179
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1649977179
transform 1 0 62928 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1649977179
transform 1 0 68080 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1649977179
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1649977179
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1649977179
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1649977179
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1649977179
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1649977179
transform 1 0 60352 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1649977179
transform 1 0 65504 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1649977179
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1649977179
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1649977179
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1649977179
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1649977179
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1649977179
transform 1 0 62928 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1649977179
transform 1 0 68080 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1649977179
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1649977179
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1649977179
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1649977179
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1649977179
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1649977179
transform 1 0 60352 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1649977179
transform 1 0 65504 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1649977179
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1649977179
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1649977179
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1649977179
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1649977179
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1649977179
transform 1 0 62928 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1649977179
transform 1 0 68080 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1649977179
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1649977179
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1649977179
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1649977179
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1649977179
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1649977179
transform 1 0 60352 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1649977179
transform 1 0 65504 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1649977179
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1649977179
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1649977179
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1649977179
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1649977179
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1649977179
transform 1 0 62928 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1649977179
transform 1 0 68080 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1649977179
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1649977179
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1649977179
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1649977179
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1649977179
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1649977179
transform 1 0 60352 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1649977179
transform 1 0 65504 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1649977179
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1649977179
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1649977179
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1649977179
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1649977179
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1649977179
transform 1 0 62928 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1649977179
transform 1 0 68080 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1649977179
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1649977179
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1649977179
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1649977179
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1649977179
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1649977179
transform 1 0 60352 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1649977179
transform 1 0 65504 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1649977179
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1649977179
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1649977179
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1649977179
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1649977179
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1649977179
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1649977179
transform 1 0 62928 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1649977179
transform 1 0 68080 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1649977179
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1649977179
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1649977179
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1649977179
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1649977179
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1649977179
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1649977179
transform 1 0 60352 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1649977179
transform 1 0 65504 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1649977179
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1649977179
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1649977179
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1649977179
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1649977179
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1649977179
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1649977179
transform 1 0 62928 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1649977179
transform 1 0 68080 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1649977179
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1649977179
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1649977179
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1649977179
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1649977179
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1649977179
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1649977179
transform 1 0 60352 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1649977179
transform 1 0 65504 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1649977179
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1649977179
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1649977179
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1649977179
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1649977179
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1649977179
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1649977179
transform 1 0 62928 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1649977179
transform 1 0 68080 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1649977179
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1649977179
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1649977179
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1649977179
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1649977179
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1649977179
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1649977179
transform 1 0 60352 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1649977179
transform 1 0 65504 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1649977179
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1649977179
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1649977179
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1649977179
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1649977179
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1649977179
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1649977179
transform 1 0 62928 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1649977179
transform 1 0 68080 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1649977179
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1649977179
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1649977179
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1649977179
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1649977179
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1649977179
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1649977179
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1649977179
transform 1 0 60352 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1649977179
transform 1 0 65504 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1649977179
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1649977179
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1649977179
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1649977179
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1649977179
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1649977179
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1649977179
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1649977179
transform 1 0 62928 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1649977179
transform 1 0 68080 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1649977179
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1649977179
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1649977179
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1649977179
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1649977179
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1649977179
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1649977179
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1649977179
transform 1 0 60352 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1649977179
transform 1 0 65504 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1649977179
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1649977179
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1649977179
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1649977179
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1649977179
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1649977179
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1649977179
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1649977179
transform 1 0 62928 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1649977179
transform 1 0 68080 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1649977179
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1649977179
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1649977179
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1649977179
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1649977179
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1649977179
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1649977179
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1649977179
transform 1 0 60352 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1649977179
transform 1 0 65504 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1649977179
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1649977179
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1649977179
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1649977179
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1649977179
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1649977179
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1649977179
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1649977179
transform 1 0 62928 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1649977179
transform 1 0 68080 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1649977179
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1649977179
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1649977179
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1649977179
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1649977179
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1649977179
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1649977179
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1649977179
transform 1 0 60352 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1649977179
transform 1 0 65504 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1649977179
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1649977179
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1649977179
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1649977179
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1649977179
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1649977179
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1649977179
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1649977179
transform 1 0 62928 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1649977179
transform 1 0 68080 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1649977179
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1649977179
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1649977179
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1649977179
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1649977179
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1649977179
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1649977179
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1649977179
transform 1 0 60352 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1649977179
transform 1 0 65504 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1649977179
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1649977179
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1649977179
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1649977179
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1649977179
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1649977179
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1649977179
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1649977179
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1649977179
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1649977179
transform 1 0 62928 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1649977179
transform 1 0 68080 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1649977179
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1649977179
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1649977179
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1649977179
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1649977179
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1649977179
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1649977179
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1649977179
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1649977179
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1649977179
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1649977179
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1649977179
transform 1 0 60352 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1649977179
transform 1 0 65504 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1649977179
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1649977179
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1649977179
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1649977179
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1649977179
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1649977179
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1649977179
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1649977179
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1649977179
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1649977179
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1649977179
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1649977179
transform 1 0 62928 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1649977179
transform 1 0 68080 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1649977179
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1649977179
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1649977179
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1649977179
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1649977179
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1649977179
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1649977179
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1649977179
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1649977179
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1649977179
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1649977179
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1649977179
transform 1 0 60352 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1649977179
transform 1 0 65504 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1649977179
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1649977179
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1649977179
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1649977179
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1649977179
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1649977179
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1649977179
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1649977179
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1649977179
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1649977179
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1649977179
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1649977179
transform 1 0 62928 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1649977179
transform 1 0 68080 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1649977179
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1649977179
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1649977179
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1649977179
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1649977179
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1649977179
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1649977179
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1649977179
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1649977179
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1649977179
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1649977179
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1649977179
transform 1 0 60352 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1649977179
transform 1 0 65504 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1649977179
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1649977179
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1649977179
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1649977179
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1649977179
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1649977179
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1649977179
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1649977179
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1649977179
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1649977179
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1649977179
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1649977179
transform 1 0 62928 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1649977179
transform 1 0 68080 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1649977179
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1649977179
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1649977179
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1649977179
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1649977179
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1649977179
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1649977179
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1649977179
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1649977179
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1649977179
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1649977179
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1649977179
transform 1 0 60352 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1649977179
transform 1 0 65504 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1649977179
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1649977179
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1649977179
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1649977179
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1649977179
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1649977179
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1649977179
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1649977179
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1649977179
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1649977179
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1649977179
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1649977179
transform 1 0 62928 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1649977179
transform 1 0 68080 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1649977179
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1649977179
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1649977179
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1649977179
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1649977179
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1649977179
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1649977179
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1649977179
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1649977179
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1649977179
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1649977179
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1649977179
transform 1 0 60352 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1649977179
transform 1 0 65504 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1649977179
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1649977179
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1649977179
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1649977179
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1649977179
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1649977179
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1649977179
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1649977179
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1649977179
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1649977179
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1649977179
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1649977179
transform 1 0 62928 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1649977179
transform 1 0 68080 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1649977179
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1649977179
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1649977179
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1649977179
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1649977179
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1649977179
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1649977179
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1649977179
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1649977179
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1649977179
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1649977179
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1649977179
transform 1 0 60352 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1649977179
transform 1 0 65504 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1649977179
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1649977179
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1649977179
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1649977179
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1649977179
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1649977179
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1649977179
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1649977179
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1649977179
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1649977179
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1649977179
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1649977179
transform 1 0 62928 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1649977179
transform 1 0 68080 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1649977179
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1649977179
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1649977179
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1649977179
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1649977179
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1649977179
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1649977179
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1649977179
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1649977179
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1649977179
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1649977179
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1649977179
transform 1 0 60352 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1649977179
transform 1 0 65504 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1649977179
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1649977179
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1649977179
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1649977179
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1649977179
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1649977179
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1649977179
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1649977179
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1649977179
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1649977179
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1649977179
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1649977179
transform 1 0 62928 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1649977179
transform 1 0 68080 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1649977179
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1649977179
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1649977179
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1649977179
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1649977179
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1649977179
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1649977179
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1649977179
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1649977179
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1649977179
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1649977179
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1649977179
transform 1 0 60352 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1649977179
transform 1 0 65504 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1649977179
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1649977179
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1649977179
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1649977179
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1649977179
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1649977179
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1649977179
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1649977179
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1649977179
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1649977179
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1649977179
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1649977179
transform 1 0 62928 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1649977179
transform 1 0 68080 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1649977179
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1649977179
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1649977179
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1649977179
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1649977179
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1649977179
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1649977179
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1649977179
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1649977179
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1649977179
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1649977179
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1649977179
transform 1 0 60352 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1649977179
transform 1 0 65504 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1649977179
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1649977179
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1649977179
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1649977179
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1649977179
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1649977179
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1649977179
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1649977179
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1649977179
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1649977179
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1649977179
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1649977179
transform 1 0 62928 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1649977179
transform 1 0 68080 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1649977179
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1649977179
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1649977179
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1649977179
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1649977179
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1649977179
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1649977179
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1649977179
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1649977179
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1649977179
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1649977179
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1649977179
transform 1 0 60352 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1649977179
transform 1 0 65504 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1649977179
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1649977179
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1649977179
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1649977179
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1649977179
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1649977179
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1649977179
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1649977179
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1649977179
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1649977179
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1649977179
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1649977179
transform 1 0 62928 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1649977179
transform 1 0 68080 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1649977179
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1649977179
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1649977179
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1649977179
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1649977179
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1649977179
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1649977179
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1649977179
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1649977179
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1649977179
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1649977179
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1649977179
transform 1 0 60352 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1649977179
transform 1 0 65504 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1649977179
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1649977179
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1649977179
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1649977179
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1649977179
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1649977179
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1649977179
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1649977179
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1649977179
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1649977179
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1649977179
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1649977179
transform 1 0 62928 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1649977179
transform 1 0 68080 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1649977179
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1649977179
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1649977179
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1649977179
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1649977179
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1649977179
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1649977179
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1649977179
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1649977179
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1649977179
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1649977179
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1649977179
transform 1 0 60352 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1649977179
transform 1 0 65504 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1649977179
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1649977179
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1649977179
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1649977179
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1649977179
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1649977179
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1649977179
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1649977179
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1649977179
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1649977179
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1649977179
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1649977179
transform 1 0 62928 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1649977179
transform 1 0 68080 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1649977179
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1649977179
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1649977179
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1649977179
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1649977179
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1649977179
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1649977179
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1649977179
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1649977179
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1649977179
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1649977179
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1649977179
transform 1 0 60352 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1649977179
transform 1 0 65504 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1649977179
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1649977179
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1649977179
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1649977179
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1649977179
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1649977179
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1649977179
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1649977179
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1649977179
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1649977179
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1649977179
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1649977179
transform 1 0 62928 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1649977179
transform 1 0 68080 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1649977179
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1649977179
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1649977179
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1649977179
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1649977179
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1649977179
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1649977179
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1649977179
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1649977179
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1649977179
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1649977179
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1649977179
transform 1 0 60352 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1649977179
transform 1 0 65504 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1649977179
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1649977179
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1649977179
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1649977179
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1649977179
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1649977179
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1649977179
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1649977179
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1649977179
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1649977179
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1649977179
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1649977179
transform 1 0 62928 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1649977179
transform 1 0 68080 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1649977179
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1649977179
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1649977179
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1649977179
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1649977179
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1649977179
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1649977179
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1649977179
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1649977179
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1649977179
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1649977179
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1649977179
transform 1 0 60352 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1649977179
transform 1 0 65504 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1649977179
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1649977179
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1649977179
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1649977179
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1649977179
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1649977179
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1649977179
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1649977179
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1649977179
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1649977179
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1649977179
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1649977179
transform 1 0 62928 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1649977179
transform 1 0 68080 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1649977179
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1649977179
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1649977179
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1649977179
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1649977179
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1649977179
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1649977179
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1649977179
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1649977179
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1649977179
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1649977179
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1649977179
transform 1 0 60352 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1649977179
transform 1 0 65504 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1649977179
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1649977179
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1649977179
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1649977179
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1649977179
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1649977179
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1649977179
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1649977179
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1649977179
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1649977179
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1649977179
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1649977179
transform 1 0 62928 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1649977179
transform 1 0 68080 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1649977179
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1649977179
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1649977179
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1649977179
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1649977179
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1649977179
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1649977179
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1649977179
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1649977179
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1649977179
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1649977179
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1649977179
transform 1 0 60352 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1649977179
transform 1 0 65504 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1649977179
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1649977179
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1649977179
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1649977179
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1649977179
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1649977179
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1649977179
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1649977179
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1649977179
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1649977179
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1649977179
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1649977179
transform 1 0 62928 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1649977179
transform 1 0 68080 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1649977179
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1649977179
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1649977179
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1649977179
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1649977179
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1649977179
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1649977179
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1649977179
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1649977179
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1649977179
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1649977179
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1649977179
transform 1 0 60352 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1649977179
transform 1 0 65504 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1649977179
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1649977179
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1649977179
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1649977179
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1649977179
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1649977179
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1649977179
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1649977179
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1649977179
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1649977179
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1649977179
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1649977179
transform 1 0 62928 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1649977179
transform 1 0 68080 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1649977179
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1649977179
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1649977179
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1649977179
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1649977179
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1649977179
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1649977179
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1649977179
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1649977179
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1649977179
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1649977179
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1649977179
transform 1 0 60352 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1649977179
transform 1 0 65504 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1649977179
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1649977179
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1649977179
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1649977179
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1649977179
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1649977179
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1649977179
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1649977179
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1649977179
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1649977179
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1649977179
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1649977179
transform 1 0 62928 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1649977179
transform 1 0 68080 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1649977179
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1649977179
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1649977179
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1649977179
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1649977179
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1649977179
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1649977179
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1649977179
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1649977179
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1649977179
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1649977179
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1649977179
transform 1 0 60352 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1649977179
transform 1 0 65504 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1649977179
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1649977179
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1649977179
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1649977179
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1649977179
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1649977179
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1649977179
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1649977179
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1649977179
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1649977179
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1649977179
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1649977179
transform 1 0 62928 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1649977179
transform 1 0 68080 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1649977179
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1649977179
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1649977179
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1649977179
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1649977179
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1649977179
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1649977179
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1649977179
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1649977179
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1649977179
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1649977179
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1649977179
transform 1 0 60352 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1649977179
transform 1 0 65504 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1649977179
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1649977179
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1649977179
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1649977179
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1649977179
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1649977179
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1649977179
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1649977179
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1649977179
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1649977179
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1649977179
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1649977179
transform 1 0 62928 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1649977179
transform 1 0 68080 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1649977179
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1649977179
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1649977179
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1649977179
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1649977179
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1649977179
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1649977179
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1649977179
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1649977179
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1649977179
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1649977179
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1649977179
transform 1 0 60352 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1649977179
transform 1 0 65504 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1649977179
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1649977179
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1649977179
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1649977179
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1649977179
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1649977179
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1649977179
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1649977179
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1649977179
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1649977179
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1649977179
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1649977179
transform 1 0 62928 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1649977179
transform 1 0 68080 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1649977179
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1649977179
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1649977179
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1649977179
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1649977179
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1649977179
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1649977179
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1649977179
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1649977179
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1649977179
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1649977179
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1649977179
transform 1 0 60352 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1649977179
transform 1 0 65504 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1649977179
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1649977179
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1649977179
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1649977179
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1649977179
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1649977179
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1649977179
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1649977179
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1649977179
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1649977179
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1649977179
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1649977179
transform 1 0 62928 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1649977179
transform 1 0 68080 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1649977179
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1649977179
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1649977179
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1649977179
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1649977179
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1649977179
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1649977179
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1649977179
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1649977179
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1649977179
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1649977179
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1649977179
transform 1 0 60352 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1649977179
transform 1 0 65504 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1649977179
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1649977179
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1649977179
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1649977179
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1649977179
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1649977179
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1649977179
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1649977179
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1649977179
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1649977179
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1649977179
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1649977179
transform 1 0 62928 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1649977179
transform 1 0 68080 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1649977179
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1649977179
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1649977179
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1649977179
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1649977179
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1649977179
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1649977179
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1649977179
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1649977179
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1649977179
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1649977179
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1649977179
transform 1 0 60352 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1649977179
transform 1 0 65504 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1348
timestamp 1649977179
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1349
timestamp 1649977179
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1350
timestamp 1649977179
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1351
timestamp 1649977179
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1352
timestamp 1649977179
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1353
timestamp 1649977179
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1354
timestamp 1649977179
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1355
timestamp 1649977179
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1356
timestamp 1649977179
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1357
timestamp 1649977179
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1358
timestamp 1649977179
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1359
timestamp 1649977179
transform 1 0 62928 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1360
timestamp 1649977179
transform 1 0 68080 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1361
timestamp 1649977179
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1362
timestamp 1649977179
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1363
timestamp 1649977179
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1364
timestamp 1649977179
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1365
timestamp 1649977179
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1366
timestamp 1649977179
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1367
timestamp 1649977179
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1368
timestamp 1649977179
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1369
timestamp 1649977179
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1370
timestamp 1649977179
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1371
timestamp 1649977179
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1372
timestamp 1649977179
transform 1 0 60352 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1373
timestamp 1649977179
transform 1 0 65504 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1374
timestamp 1649977179
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1375
timestamp 1649977179
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1376
timestamp 1649977179
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1377
timestamp 1649977179
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1378
timestamp 1649977179
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1379
timestamp 1649977179
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1380
timestamp 1649977179
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1381
timestamp 1649977179
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1382
timestamp 1649977179
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1383
timestamp 1649977179
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1384
timestamp 1649977179
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1385
timestamp 1649977179
transform 1 0 62928 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1386
timestamp 1649977179
transform 1 0 68080 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1387
timestamp 1649977179
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1388
timestamp 1649977179
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1389
timestamp 1649977179
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1390
timestamp 1649977179
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1391
timestamp 1649977179
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1392
timestamp 1649977179
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1393
timestamp 1649977179
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1394
timestamp 1649977179
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1395
timestamp 1649977179
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1396
timestamp 1649977179
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1397
timestamp 1649977179
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1398
timestamp 1649977179
transform 1 0 60352 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1399
timestamp 1649977179
transform 1 0 65504 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1400
timestamp 1649977179
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1401
timestamp 1649977179
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1402
timestamp 1649977179
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1403
timestamp 1649977179
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1404
timestamp 1649977179
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1405
timestamp 1649977179
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1406
timestamp 1649977179
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1407
timestamp 1649977179
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1408
timestamp 1649977179
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1409
timestamp 1649977179
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1410
timestamp 1649977179
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1411
timestamp 1649977179
transform 1 0 62928 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1412
timestamp 1649977179
transform 1 0 68080 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1413
timestamp 1649977179
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1414
timestamp 1649977179
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1415
timestamp 1649977179
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1416
timestamp 1649977179
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1417
timestamp 1649977179
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1418
timestamp 1649977179
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1419
timestamp 1649977179
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1420
timestamp 1649977179
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1421
timestamp 1649977179
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1422
timestamp 1649977179
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1423
timestamp 1649977179
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1424
timestamp 1649977179
transform 1 0 60352 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1425
timestamp 1649977179
transform 1 0 65504 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1426
timestamp 1649977179
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1427
timestamp 1649977179
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1428
timestamp 1649977179
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1429
timestamp 1649977179
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1430
timestamp 1649977179
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1431
timestamp 1649977179
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1432
timestamp 1649977179
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1433
timestamp 1649977179
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1434
timestamp 1649977179
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1435
timestamp 1649977179
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1436
timestamp 1649977179
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1437
timestamp 1649977179
transform 1 0 62928 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1438
timestamp 1649977179
transform 1 0 68080 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1439
timestamp 1649977179
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1440
timestamp 1649977179
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1441
timestamp 1649977179
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1442
timestamp 1649977179
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1443
timestamp 1649977179
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1444
timestamp 1649977179
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1445
timestamp 1649977179
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1446
timestamp 1649977179
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1447
timestamp 1649977179
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1448
timestamp 1649977179
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1449
timestamp 1649977179
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1450
timestamp 1649977179
transform 1 0 60352 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1451
timestamp 1649977179
transform 1 0 65504 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1452
timestamp 1649977179
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1453
timestamp 1649977179
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1454
timestamp 1649977179
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1455
timestamp 1649977179
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1456
timestamp 1649977179
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1457
timestamp 1649977179
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1458
timestamp 1649977179
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1459
timestamp 1649977179
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1460
timestamp 1649977179
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1461
timestamp 1649977179
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1462
timestamp 1649977179
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1463
timestamp 1649977179
transform 1 0 62928 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1464
timestamp 1649977179
transform 1 0 68080 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1465
timestamp 1649977179
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1466
timestamp 1649977179
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1467
timestamp 1649977179
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1468
timestamp 1649977179
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1469
timestamp 1649977179
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1470
timestamp 1649977179
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1471
timestamp 1649977179
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1472
timestamp 1649977179
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1473
timestamp 1649977179
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1474
timestamp 1649977179
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1475
timestamp 1649977179
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1476
timestamp 1649977179
transform 1 0 60352 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1477
timestamp 1649977179
transform 1 0 65504 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1478
timestamp 1649977179
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1479
timestamp 1649977179
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1480
timestamp 1649977179
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1481
timestamp 1649977179
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1482
timestamp 1649977179
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1483
timestamp 1649977179
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1484
timestamp 1649977179
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1485
timestamp 1649977179
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1486
timestamp 1649977179
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1487
timestamp 1649977179
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1488
timestamp 1649977179
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1489
timestamp 1649977179
transform 1 0 62928 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1490
timestamp 1649977179
transform 1 0 68080 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1491
timestamp 1649977179
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1492
timestamp 1649977179
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1493
timestamp 1649977179
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1494
timestamp 1649977179
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1495
timestamp 1649977179
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1496
timestamp 1649977179
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1497
timestamp 1649977179
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1498
timestamp 1649977179
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1499
timestamp 1649977179
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1500
timestamp 1649977179
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1501
timestamp 1649977179
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1502
timestamp 1649977179
transform 1 0 60352 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1503
timestamp 1649977179
transform 1 0 65504 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1504
timestamp 1649977179
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1505
timestamp 1649977179
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1506
timestamp 1649977179
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1507
timestamp 1649977179
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1508
timestamp 1649977179
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1509
timestamp 1649977179
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1510
timestamp 1649977179
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1511
timestamp 1649977179
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1512
timestamp 1649977179
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1513
timestamp 1649977179
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1514
timestamp 1649977179
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1515
timestamp 1649977179
transform 1 0 62928 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1516
timestamp 1649977179
transform 1 0 68080 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1517
timestamp 1649977179
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1518
timestamp 1649977179
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1519
timestamp 1649977179
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1520
timestamp 1649977179
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1521
timestamp 1649977179
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1522
timestamp 1649977179
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1523
timestamp 1649977179
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1524
timestamp 1649977179
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1525
timestamp 1649977179
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1526
timestamp 1649977179
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1527
timestamp 1649977179
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1528
timestamp 1649977179
transform 1 0 60352 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1529
timestamp 1649977179
transform 1 0 65504 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1530
timestamp 1649977179
transform 1 0 3680 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1531
timestamp 1649977179
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1532
timestamp 1649977179
transform 1 0 8832 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1533
timestamp 1649977179
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1534
timestamp 1649977179
transform 1 0 13984 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1535
timestamp 1649977179
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1536
timestamp 1649977179
transform 1 0 19136 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1537
timestamp 1649977179
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1538
timestamp 1649977179
transform 1 0 24288 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1539
timestamp 1649977179
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1540
timestamp 1649977179
transform 1 0 29440 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1541
timestamp 1649977179
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1542
timestamp 1649977179
transform 1 0 34592 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1543
timestamp 1649977179
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1544
timestamp 1649977179
transform 1 0 39744 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1545
timestamp 1649977179
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1546
timestamp 1649977179
transform 1 0 44896 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1547
timestamp 1649977179
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1548
timestamp 1649977179
transform 1 0 50048 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1549
timestamp 1649977179
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1550
timestamp 1649977179
transform 1 0 55200 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1551
timestamp 1649977179
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1552
timestamp 1649977179
transform 1 0 60352 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1553
timestamp 1649977179
transform 1 0 62928 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1554
timestamp 1649977179
transform 1 0 65504 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1555
timestamp 1649977179
transform 1 0 68080 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _0790_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8832 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0791_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 7360 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__or4_4  _0792_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0793_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 13248 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0794_
timestamp 1649977179
transform -1 0 11776 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0795_
timestamp 1649977179
transform 1 0 12696 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0796_
timestamp 1649977179
transform 1 0 14168 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__or4_2  _0797_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _0798_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0799_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9752 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0800_
timestamp 1649977179
transform 1 0 10580 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0801_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 12236 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0802_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 6808 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0803_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0804_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 5704 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0805_
timestamp 1649977179
transform -1 0 5060 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0806_
timestamp 1649977179
transform 1 0 6900 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0807_
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0808_
timestamp 1649977179
transform 1 0 1840 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0809_
timestamp 1649977179
transform -1 0 2024 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0810_
timestamp 1649977179
transform -1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0811_
timestamp 1649977179
transform 1 0 1656 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0812_
timestamp 1649977179
transform 1 0 1656 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0813_
timestamp 1649977179
transform -1 0 2392 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0814_
timestamp 1649977179
transform 1 0 4784 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0815_
timestamp 1649977179
transform 1 0 1656 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0816_
timestamp 1649977179
transform -1 0 2208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0817_
timestamp 1649977179
transform 1 0 2024 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0818_
timestamp 1649977179
transform 1 0 1748 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0819_
timestamp 1649977179
transform -1 0 2484 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0820_
timestamp 1649977179
transform 1 0 7176 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0821_
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0822_
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0823_
timestamp 1649977179
transform -1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0824_
timestamp 1649977179
transform -1 0 8188 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0825_
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0826_
timestamp 1649977179
transform 1 0 18952 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0827_
timestamp 1649977179
transform -1 0 20056 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0828_
timestamp 1649977179
transform -1 0 18768 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0829_
timestamp 1649977179
transform 1 0 18492 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0830_
timestamp 1649977179
transform -1 0 19596 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0831_
timestamp 1649977179
transform 1 0 15456 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0832_
timestamp 1649977179
transform -1 0 15824 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0833_
timestamp 1649977179
transform -1 0 15272 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0834_
timestamp 1649977179
transform 1 0 6440 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0835_
timestamp 1649977179
transform -1 0 5888 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0836_
timestamp 1649977179
transform 1 0 4784 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0837_
timestamp 1649977179
transform 1 0 7176 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0838_
timestamp 1649977179
transform -1 0 6808 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0839_
timestamp 1649977179
transform -1 0 3312 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0840_
timestamp 1649977179
transform -1 0 5980 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0841_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 12788 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0842_
timestamp 1649977179
transform -1 0 6532 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__or4b_4  _0843_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11408 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_2  _0844_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0845_
timestamp 1649977179
transform 1 0 14168 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0846_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 6624 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0847_
timestamp 1649977179
transform -1 0 3680 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0848_
timestamp 1649977179
transform -1 0 5888 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0849_
timestamp 1649977179
transform 1 0 2116 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0850_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2852 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0851_
timestamp 1649977179
transform 1 0 6532 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0852_
timestamp 1649977179
transform -1 0 2944 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0853_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 3128 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0854_
timestamp 1649977179
transform 1 0 3588 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0855_
timestamp 1649977179
transform 1 0 3772 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0856_
timestamp 1649977179
transform -1 0 4508 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0857_
timestamp 1649977179
transform -1 0 1932 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0858_
timestamp 1649977179
transform 1 0 1564 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0859_
timestamp 1649977179
transform -1 0 2668 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0860_
timestamp 1649977179
transform 1 0 7268 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0861_
timestamp 1649977179
transform 1 0 2852 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0862_
timestamp 1649977179
transform -1 0 4508 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0863_
timestamp 1649977179
transform -1 0 3220 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0864_
timestamp 1649977179
transform 1 0 1656 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0865_
timestamp 1649977179
transform -1 0 2576 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0866_
timestamp 1649977179
transform 1 0 5704 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0867_
timestamp 1649977179
transform -1 0 3312 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0868_
timestamp 1649977179
transform 1 0 2024 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0869_
timestamp 1649977179
transform 1 0 1472 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0870_
timestamp 1649977179
transform -1 0 2668 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0871_
timestamp 1649977179
transform -1 0 3036 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0872_
timestamp 1649977179
transform -1 0 12696 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0873_
timestamp 1649977179
transform 1 0 1840 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0874_
timestamp 1649977179
transform -1 0 2944 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0875_
timestamp 1649977179
transform 1 0 13156 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0876_
timestamp 1649977179
transform 1 0 1380 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0877_
timestamp 1649977179
transform -1 0 3772 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0878_
timestamp 1649977179
transform -1 0 13708 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0879_
timestamp 1649977179
transform 1 0 1564 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0880_
timestamp 1649977179
transform -1 0 3036 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0881_
timestamp 1649977179
transform -1 0 7452 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0882_
timestamp 1649977179
transform 1 0 1656 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0883_
timestamp 1649977179
transform -1 0 2484 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0884_
timestamp 1649977179
transform -1 0 9568 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0885_
timestamp 1649977179
transform -1 0 5520 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0886_
timestamp 1649977179
transform -1 0 2668 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0887_
timestamp 1649977179
transform 1 0 4692 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_4  _0888_
timestamp 1649977179
transform 1 0 11776 0 -1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _0889_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12512 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0890_
timestamp 1649977179
transform -1 0 9016 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0891_
timestamp 1649977179
transform -1 0 6624 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0892_
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0893_
timestamp 1649977179
transform -1 0 16468 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0894_
timestamp 1649977179
transform -1 0 7636 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0895_
timestamp 1649977179
transform 1 0 4508 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0896_
timestamp 1649977179
transform -1 0 4600 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0897_
timestamp 1649977179
transform -1 0 2576 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0898_
timestamp 1649977179
transform 1 0 2116 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0899_
timestamp 1649977179
transform -1 0 2852 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0900_
timestamp 1649977179
transform -1 0 2208 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0901_
timestamp 1649977179
transform -1 0 2576 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0902_
timestamp 1649977179
transform 1 0 4600 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0903_
timestamp 1649977179
transform -1 0 5060 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0904_
timestamp 1649977179
transform -1 0 2208 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0905_
timestamp 1649977179
transform -1 0 2300 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0906_
timestamp 1649977179
transform -1 0 2484 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0907_
timestamp 1649977179
transform -1 0 2760 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0908_
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0909_
timestamp 1649977179
transform -1 0 2300 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0910_
timestamp 1649977179
transform -1 0 2484 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0911_
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0912_
timestamp 1649977179
transform -1 0 2760 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0913_
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0914_
timestamp 1649977179
transform -1 0 2576 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0915_
timestamp 1649977179
transform -1 0 2392 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0916_
timestamp 1649977179
transform -1 0 2668 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0917_
timestamp 1649977179
transform -1 0 2484 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0918_
timestamp 1649977179
transform -1 0 14168 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0919_
timestamp 1649977179
transform 1 0 6992 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0920_
timestamp 1649977179
transform -1 0 6716 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0921_
timestamp 1649977179
transform -1 0 2668 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0922_
timestamp 1649977179
transform 1 0 4232 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0923_
timestamp 1649977179
transform -1 0 5796 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_2  _0924_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11776 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0925_
timestamp 1649977179
transform 1 0 13064 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0926_
timestamp 1649977179
transform 1 0 9936 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0927_
timestamp 1649977179
transform -1 0 9200 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0928_
timestamp 1649977179
transform 1 0 7544 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0929_
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0930_
timestamp 1649977179
transform -1 0 7176 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0931_
timestamp 1649977179
transform 1 0 1840 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0932_
timestamp 1649977179
transform -1 0 2760 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0933_
timestamp 1649977179
transform 1 0 1840 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0934_
timestamp 1649977179
transform -1 0 2760 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0935_
timestamp 1649977179
transform -1 0 6808 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0936_
timestamp 1649977179
transform -1 0 5888 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0937_
timestamp 1649977179
transform 1 0 7452 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0938_
timestamp 1649977179
transform 1 0 6992 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0939_
timestamp 1649977179
transform -1 0 7912 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0940_
timestamp 1649977179
transform -1 0 7636 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0941_
timestamp 1649977179
transform -1 0 7360 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0942_
timestamp 1649977179
transform -1 0 8004 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0943_
timestamp 1649977179
transform 1 0 6440 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0944_
timestamp 1649977179
transform -1 0 8188 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0945_
timestamp 1649977179
transform -1 0 8372 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0946_
timestamp 1649977179
transform 1 0 7176 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0947_
timestamp 1649977179
transform -1 0 8188 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0948_
timestamp 1649977179
transform 1 0 6164 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0949_
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0950_
timestamp 1649977179
transform -1 0 5888 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0951_
timestamp 1649977179
transform 1 0 6164 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0952_
timestamp 1649977179
transform 1 0 6164 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0953_
timestamp 1649977179
transform 1 0 7912 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0954_
timestamp 1649977179
transform -1 0 8280 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0955_
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0956_
timestamp 1649977179
transform -1 0 8464 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_4  _0957_
timestamp 1649977179
transform 1 0 13432 0 -1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_2  _0958_
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0959_
timestamp 1649977179
transform 1 0 15732 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0960_
timestamp 1649977179
transform -1 0 6808 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0961_
timestamp 1649977179
transform -1 0 7360 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0962_
timestamp 1649977179
transform 1 0 6900 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0963_
timestamp 1649977179
transform -1 0 7176 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0964_
timestamp 1649977179
transform -1 0 8372 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0965_
timestamp 1649977179
transform -1 0 8188 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0966_
timestamp 1649977179
transform -1 0 7544 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0967_
timestamp 1649977179
transform -1 0 7176 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0968_
timestamp 1649977179
transform 1 0 9476 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0969_
timestamp 1649977179
transform 1 0 6808 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0970_
timestamp 1649977179
transform -1 0 10304 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0971_
timestamp 1649977179
transform 1 0 9660 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0972_
timestamp 1649977179
transform -1 0 10212 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0973_
timestamp 1649977179
transform -1 0 9844 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0974_
timestamp 1649977179
transform -1 0 8004 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0975_
timestamp 1649977179
transform 1 0 6900 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0976_
timestamp 1649977179
transform -1 0 8372 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0977_
timestamp 1649977179
transform 1 0 8924 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0978_
timestamp 1649977179
transform -1 0 8464 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0979_
timestamp 1649977179
transform -1 0 8188 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0980_
timestamp 1649977179
transform 1 0 6992 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0981_
timestamp 1649977179
transform 1 0 8004 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0982_
timestamp 1649977179
transform -1 0 7360 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0983_
timestamp 1649977179
transform -1 0 9200 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0984_
timestamp 1649977179
transform -1 0 7636 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0985_
timestamp 1649977179
transform -1 0 8924 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0986_
timestamp 1649977179
transform 1 0 8924 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0987_
timestamp 1649977179
transform -1 0 9568 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0988_
timestamp 1649977179
transform -1 0 8372 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0989_
timestamp 1649977179
transform 1 0 6808 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _0990_
timestamp 1649977179
transform -1 0 15732 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0991_
timestamp 1649977179
transform -1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0992_
timestamp 1649977179
transform 1 0 7360 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0993_
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0994_
timestamp 1649977179
transform 1 0 8004 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0995_
timestamp 1649977179
transform 1 0 8188 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0996_
timestamp 1649977179
transform -1 0 9384 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0997_
timestamp 1649977179
transform 1 0 7728 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0998_
timestamp 1649977179
transform 1 0 9844 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0999_
timestamp 1649977179
transform 1 0 14444 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1000_
timestamp 1649977179
transform -1 0 12696 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1001_
timestamp 1649977179
transform 1 0 9568 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1002_
timestamp 1649977179
transform 1 0 11592 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1003_
timestamp 1649977179
transform -1 0 12420 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1004_
timestamp 1649977179
transform -1 0 11960 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1005_
timestamp 1649977179
transform -1 0 11040 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1006_
timestamp 1649977179
transform 1 0 8004 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1007_
timestamp 1649977179
transform -1 0 9200 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1008_
timestamp 1649977179
transform 1 0 9660 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1009_
timestamp 1649977179
transform -1 0 10488 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1010_
timestamp 1649977179
transform 1 0 12788 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1011_
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1012_
timestamp 1649977179
transform 1 0 10488 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1013_
timestamp 1649977179
transform 1 0 12328 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1014_
timestamp 1649977179
transform -1 0 10948 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1015_
timestamp 1649977179
transform 1 0 12788 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1016_
timestamp 1649977179
transform -1 0 14076 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1017_
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1018_
timestamp 1649977179
transform 1 0 12604 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1019_
timestamp 1649977179
transform 1 0 11684 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1020_
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1021_
timestamp 1649977179
transform 1 0 8832 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1022_
timestamp 1649977179
transform -1 0 10120 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1023_
timestamp 1649977179
transform 1 0 22172 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1024_
timestamp 1649977179
transform 1 0 22080 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1025_
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1026_
timestamp 1649977179
transform -1 0 26496 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1027_
timestamp 1649977179
transform 1 0 24012 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1028_
timestamp 1649977179
transform 1 0 24840 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1029_
timestamp 1649977179
transform 1 0 22816 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1030_
timestamp 1649977179
transform -1 0 23920 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1031_
timestamp 1649977179
transform 1 0 24564 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1032_
timestamp 1649977179
transform -1 0 25668 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1033_
timestamp 1649977179
transform 1 0 24748 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1034_
timestamp 1649977179
transform 1 0 23000 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1035_
timestamp 1649977179
transform 1 0 24288 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1036_
timestamp 1649977179
transform 1 0 24656 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1037_
timestamp 1649977179
transform 1 0 25760 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1038_
timestamp 1649977179
transform 1 0 24932 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1039_
timestamp 1649977179
transform -1 0 26128 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1040_
timestamp 1649977179
transform 1 0 24380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1041_
timestamp 1649977179
transform 1 0 25300 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1042_
timestamp 1649977179
transform -1 0 26036 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1043_
timestamp 1649977179
transform 1 0 21068 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1044_
timestamp 1649977179
transform 1 0 25668 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1045_
timestamp 1649977179
transform -1 0 26864 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1046_
timestamp 1649977179
transform 1 0 23736 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1047_
timestamp 1649977179
transform -1 0 25208 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1048_
timestamp 1649977179
transform -1 0 24656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1049_
timestamp 1649977179
transform 1 0 29256 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1050_
timestamp 1649977179
transform -1 0 25944 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1051_
timestamp 1649977179
transform -1 0 30268 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1052_
timestamp 1649977179
transform 1 0 27876 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1053_
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1054_
timestamp 1649977179
transform -1 0 30544 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1055_
timestamp 1649977179
transform 1 0 26312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1056_
timestamp 1649977179
transform 1 0 28612 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1057_
timestamp 1649977179
transform -1 0 29808 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1058_
timestamp 1649977179
transform 1 0 24840 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1059_
timestamp 1649977179
transform 1 0 25576 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1060_
timestamp 1649977179
transform -1 0 27140 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1061_
timestamp 1649977179
transform 1 0 25484 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1062_
timestamp 1649977179
transform 1 0 24288 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1063_
timestamp 1649977179
transform 1 0 25116 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1064_
timestamp 1649977179
transform 1 0 20700 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1065_
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1066_
timestamp 1649977179
transform -1 0 25576 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1067_
timestamp 1649977179
transform 1 0 24104 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1068_
timestamp 1649977179
transform 1 0 15548 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1069_
timestamp 1649977179
transform -1 0 26404 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1070_
timestamp 1649977179
transform 1 0 29624 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1071_
timestamp 1649977179
transform 1 0 32752 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1072_
timestamp 1649977179
transform 1 0 17020 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1073_
timestamp 1649977179
transform 1 0 28796 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1074_
timestamp 1649977179
transform -1 0 32384 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1075_
timestamp 1649977179
transform 1 0 33948 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1076_
timestamp 1649977179
transform -1 0 35788 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1077_
timestamp 1649977179
transform 1 0 34500 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1078_
timestamp 1649977179
transform -1 0 35696 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1079_
timestamp 1649977179
transform 1 0 32936 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1080_
timestamp 1649977179
transform -1 0 33672 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1081_
timestamp 1649977179
transform 1 0 34684 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1082_
timestamp 1649977179
transform -1 0 35880 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1083_
timestamp 1649977179
transform -1 0 34500 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1084_
timestamp 1649977179
transform 1 0 31648 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1085_
timestamp 1649977179
transform -1 0 31648 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1086_
timestamp 1649977179
transform -1 0 33948 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1087_
timestamp 1649977179
transform 1 0 29624 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1088_
timestamp 1649977179
transform 1 0 28796 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1089_
timestamp 1649977179
transform 1 0 25116 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1090_
timestamp 1649977179
transform 1 0 25760 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1091_
timestamp 1649977179
transform -1 0 28888 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1092_
timestamp 1649977179
transform 1 0 27324 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1093_
timestamp 1649977179
transform -1 0 24932 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1094_
timestamp 1649977179
transform 1 0 25024 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1095_
timestamp 1649977179
transform 1 0 24840 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1096_
timestamp 1649977179
transform -1 0 26220 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1097_
timestamp 1649977179
transform 1 0 29532 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1098_
timestamp 1649977179
transform -1 0 31280 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1099_
timestamp 1649977179
transform 1 0 29532 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1100_
timestamp 1649977179
transform 1 0 30820 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1101_
timestamp 1649977179
transform -1 0 31556 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_4  _1102_
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_2  _1103_
timestamp 1649977179
transform 1 0 18308 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1104_
timestamp 1649977179
transform -1 0 36248 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1105_
timestamp 1649977179
transform -1 0 35788 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1106_
timestamp 1649977179
transform 1 0 35880 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1107_
timestamp 1649977179
transform 1 0 35052 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1108_
timestamp 1649977179
transform -1 0 37536 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1109_
timestamp 1649977179
transform 1 0 37352 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1110_
timestamp 1649977179
transform -1 0 38364 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1111_
timestamp 1649977179
transform 1 0 38456 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1112_
timestamp 1649977179
transform -1 0 38456 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1113_
timestamp 1649977179
transform 1 0 36524 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1114_
timestamp 1649977179
transform -1 0 38088 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1115_
timestamp 1649977179
transform 1 0 36340 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1116_
timestamp 1649977179
transform -1 0 37168 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1117_
timestamp 1649977179
transform -1 0 38180 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1118_
timestamp 1649977179
transform 1 0 37904 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1119_
timestamp 1649977179
transform -1 0 38732 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1120_
timestamp 1649977179
transform -1 0 35604 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1121_
timestamp 1649977179
transform -1 0 34960 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1122_
timestamp 1649977179
transform 1 0 37260 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1123_
timestamp 1649977179
transform -1 0 38824 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1124_
timestamp 1649977179
transform 1 0 37260 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1125_
timestamp 1649977179
transform -1 0 37812 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1126_
timestamp 1649977179
transform 1 0 35788 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1127_
timestamp 1649977179
transform 1 0 35788 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1128_
timestamp 1649977179
transform -1 0 33212 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1129_
timestamp 1649977179
transform -1 0 33948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1130_
timestamp 1649977179
transform 1 0 32844 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1131_
timestamp 1649977179
transform -1 0 35144 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1132_
timestamp 1649977179
transform 1 0 33948 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1133_
timestamp 1649977179
transform -1 0 33580 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1134_
timestamp 1649977179
transform 1 0 33120 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1135_
timestamp 1649977179
transform 1 0 18400 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1136_
timestamp 1649977179
transform 1 0 35420 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1137_
timestamp 1649977179
transform -1 0 34960 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1138_
timestamp 1649977179
transform 1 0 35328 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1139_
timestamp 1649977179
transform -1 0 35144 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1140_
timestamp 1649977179
transform 1 0 34776 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1141_
timestamp 1649977179
transform -1 0 34868 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1142_
timestamp 1649977179
transform -1 0 36064 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1143_
timestamp 1649977179
transform -1 0 35972 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1144_
timestamp 1649977179
transform 1 0 35052 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1145_
timestamp 1649977179
transform 1 0 38732 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1146_
timestamp 1649977179
transform 1 0 37260 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1147_
timestamp 1649977179
transform -1 0 38548 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1148_
timestamp 1649977179
transform -1 0 39008 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1149_
timestamp 1649977179
transform -1 0 38364 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1150_
timestamp 1649977179
transform 1 0 37628 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1151_
timestamp 1649977179
transform -1 0 38548 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1152_
timestamp 1649977179
transform 1 0 35696 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1153_
timestamp 1649977179
transform -1 0 35144 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1154_
timestamp 1649977179
transform -1 0 38640 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1155_
timestamp 1649977179
transform -1 0 38640 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1156_
timestamp 1649977179
transform 1 0 38456 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1157_
timestamp 1649977179
transform -1 0 38640 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1158_
timestamp 1649977179
transform -1 0 36708 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1159_
timestamp 1649977179
transform -1 0 31648 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1160_
timestamp 1649977179
transform 1 0 31188 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1161_
timestamp 1649977179
transform 1 0 35144 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1162_
timestamp 1649977179
transform -1 0 34040 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1163_
timestamp 1649977179
transform 1 0 33488 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1164_
timestamp 1649977179
transform -1 0 34868 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1165_
timestamp 1649977179
transform 1 0 33580 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1166_
timestamp 1649977179
transform -1 0 33672 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1167_
timestamp 1649977179
transform 1 0 33212 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1168_
timestamp 1649977179
transform 1 0 15916 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1169_
timestamp 1649977179
transform 1 0 29532 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1170_
timestamp 1649977179
transform -1 0 29072 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1171_
timestamp 1649977179
transform 1 0 35236 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1172_
timestamp 1649977179
transform -1 0 31372 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1173_
timestamp 1649977179
transform -1 0 35972 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1174_
timestamp 1649977179
transform -1 0 36892 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1175_
timestamp 1649977179
transform 1 0 35328 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1176_
timestamp 1649977179
transform 1 0 37444 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1177_
timestamp 1649977179
transform 1 0 33120 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1178_
timestamp 1649977179
transform -1 0 38272 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1179_
timestamp 1649977179
transform 1 0 37720 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1180_
timestamp 1649977179
transform -1 0 39284 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1181_
timestamp 1649977179
transform 1 0 38916 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1182_
timestamp 1649977179
transform -1 0 38548 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1183_
timestamp 1649977179
transform 1 0 37720 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1184_
timestamp 1649977179
transform -1 0 38548 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1185_
timestamp 1649977179
transform -1 0 33120 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1186_
timestamp 1649977179
transform -1 0 30912 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1187_
timestamp 1649977179
transform 1 0 33488 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1188_
timestamp 1649977179
transform -1 0 34592 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1189_
timestamp 1649977179
transform 1 0 32200 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1190_
timestamp 1649977179
transform -1 0 32844 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1191_
timestamp 1649977179
transform -1 0 33212 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1192_
timestamp 1649977179
transform 1 0 31832 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1193_
timestamp 1649977179
transform 1 0 32200 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1194_
timestamp 1649977179
transform 1 0 32108 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1195_
timestamp 1649977179
transform -1 0 33304 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1196_
timestamp 1649977179
transform 1 0 31188 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1197_
timestamp 1649977179
transform 1 0 32384 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1198_
timestamp 1649977179
transform 1 0 32108 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1199_
timestamp 1649977179
transform -1 0 33028 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1200_
timestamp 1649977179
transform 1 0 20976 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1201_
timestamp 1649977179
transform 1 0 17756 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1202_
timestamp 1649977179
transform -1 0 15548 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1203_
timestamp 1649977179
transform 1 0 20424 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1204_
timestamp 1649977179
transform -1 0 23460 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1205_
timestamp 1649977179
transform -1 0 23644 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1206_
timestamp 1649977179
transform 1 0 20884 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1207_
timestamp 1649977179
transform -1 0 22908 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1208_
timestamp 1649977179
transform 1 0 23368 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1209_
timestamp 1649977179
transform -1 0 24932 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1210_
timestamp 1649977179
transform 1 0 23460 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1211_
timestamp 1649977179
transform -1 0 21896 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1212_
timestamp 1649977179
transform 1 0 23460 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1213_
timestamp 1649977179
transform -1 0 24932 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1214_
timestamp 1649977179
transform -1 0 25208 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1215_
timestamp 1649977179
transform 1 0 26128 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1216_
timestamp 1649977179
transform -1 0 25760 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1217_
timestamp 1649977179
transform 1 0 25484 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1218_
timestamp 1649977179
transform 1 0 24656 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1219_
timestamp 1649977179
transform -1 0 25852 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1220_
timestamp 1649977179
transform -1 0 17020 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1221_
timestamp 1649977179
transform 1 0 23092 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1222_
timestamp 1649977179
transform -1 0 23920 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1223_
timestamp 1649977179
transform -1 0 15916 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1224_
timestamp 1649977179
transform -1 0 22724 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1225_
timestamp 1649977179
transform 1 0 20884 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1226_
timestamp 1649977179
transform 1 0 20332 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1227_
timestamp 1649977179
transform -1 0 25024 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1228_
timestamp 1649977179
transform -1 0 20976 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1229_
timestamp 1649977179
transform 1 0 13064 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1230_
timestamp 1649977179
transform 1 0 18308 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1231_
timestamp 1649977179
transform -1 0 19964 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1232_
timestamp 1649977179
transform -1 0 14444 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1233_
timestamp 1649977179
transform -1 0 18216 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1234_
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1235_
timestamp 1649977179
transform -1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1236_
timestamp 1649977179
transform 1 0 15180 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1237_
timestamp 1649977179
transform 1 0 15456 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1238_
timestamp 1649977179
transform -1 0 13800 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1239_
timestamp 1649977179
transform -1 0 14996 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1240_
timestamp 1649977179
transform 1 0 15364 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1241_
timestamp 1649977179
transform -1 0 16008 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1242_
timestamp 1649977179
transform 1 0 22356 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1243_
timestamp 1649977179
transform -1 0 21988 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1244_
timestamp 1649977179
transform -1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1245_
timestamp 1649977179
transform -1 0 23368 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _1246_
timestamp 1649977179
transform 1 0 13616 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _1247_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16284 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1248_
timestamp 1649977179
transform -1 0 28244 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1249_
timestamp 1649977179
transform -1 0 28796 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1250_
timestamp 1649977179
transform 1 0 29532 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1251_
timestamp 1649977179
transform 1 0 15824 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1252_
timestamp 1649977179
transform 1 0 28612 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1253_
timestamp 1649977179
transform -1 0 31096 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1254_
timestamp 1649977179
transform -1 0 30360 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1255_
timestamp 1649977179
transform 1 0 28796 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1256_
timestamp 1649977179
transform 1 0 30728 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1257_
timestamp 1649977179
transform -1 0 31648 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1258_
timestamp 1649977179
transform 1 0 31188 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1259_
timestamp 1649977179
transform -1 0 30820 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1260_
timestamp 1649977179
transform 1 0 30912 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1261_
timestamp 1649977179
transform -1 0 31832 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1262_
timestamp 1649977179
transform 1 0 29992 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1263_
timestamp 1649977179
transform 1 0 26220 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1264_
timestamp 1649977179
transform -1 0 30912 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1265_
timestamp 1649977179
transform 1 0 29164 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1266_
timestamp 1649977179
transform -1 0 29808 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1267_
timestamp 1649977179
transform 1 0 29992 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1268_
timestamp 1649977179
transform -1 0 31188 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1269_
timestamp 1649977179
transform 1 0 30268 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1270_
timestamp 1649977179
transform -1 0 31832 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1271_
timestamp 1649977179
transform -1 0 29992 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1272_
timestamp 1649977179
transform -1 0 29072 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1273_
timestamp 1649977179
transform -1 0 27784 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1274_
timestamp 1649977179
transform -1 0 27140 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1275_
timestamp 1649977179
transform -1 0 28152 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1276_
timestamp 1649977179
transform -1 0 25668 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1277_
timestamp 1649977179
transform 1 0 26956 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1278_
timestamp 1649977179
transform -1 0 29440 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1279_
timestamp 1649977179
transform -1 0 28152 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1280_
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1281_
timestamp 1649977179
transform 1 0 17848 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1282_
timestamp 1649977179
transform 1 0 19228 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1283_
timestamp 1649977179
transform 1 0 20148 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1284_
timestamp 1649977179
transform -1 0 18768 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1285_
timestamp 1649977179
transform -1 0 21252 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1286_
timestamp 1649977179
transform 1 0 21804 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1287_
timestamp 1649977179
transform -1 0 22632 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1288_
timestamp 1649977179
transform 1 0 20516 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1289_
timestamp 1649977179
transform 1 0 21344 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1290_
timestamp 1649977179
transform 1 0 23092 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1291_
timestamp 1649977179
transform -1 0 24196 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1292_
timestamp 1649977179
transform -1 0 19688 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1293_
timestamp 1649977179
transform -1 0 21068 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1294_
timestamp 1649977179
transform -1 0 20792 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1295_
timestamp 1649977179
transform 1 0 22080 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1296_
timestamp 1649977179
transform 1 0 21988 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1297_
timestamp 1649977179
transform 1 0 19964 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1298_
timestamp 1649977179
transform 1 0 19228 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1299_
timestamp 1649977179
transform 1 0 20148 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1300_
timestamp 1649977179
transform -1 0 22540 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1301_
timestamp 1649977179
transform 1 0 18676 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1302_
timestamp 1649977179
transform -1 0 20240 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1303_
timestamp 1649977179
transform 1 0 19228 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1304_
timestamp 1649977179
transform -1 0 20148 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1305_
timestamp 1649977179
transform 1 0 18032 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1306_
timestamp 1649977179
transform 1 0 21804 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1307_
timestamp 1649977179
transform 1 0 19228 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1308_
timestamp 1649977179
transform 1 0 18308 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1309_
timestamp 1649977179
transform 1 0 18584 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1310_
timestamp 1649977179
transform 1 0 18124 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1311_
timestamp 1649977179
transform 1 0 18952 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1312_
timestamp 1649977179
transform 1 0 13064 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1313_
timestamp 1649977179
transform 1 0 15272 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1314_
timestamp 1649977179
transform 1 0 17480 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1315_
timestamp 1649977179
transform -1 0 16192 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1316_
timestamp 1649977179
transform -1 0 15088 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1317_
timestamp 1649977179
transform -1 0 15456 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1318_
timestamp 1649977179
transform 1 0 19228 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1319_
timestamp 1649977179
transform -1 0 20056 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1320_
timestamp 1649977179
transform 1 0 17388 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1321_
timestamp 1649977179
transform 1 0 18216 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1322_
timestamp 1649977179
transform 1 0 15088 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1323_
timestamp 1649977179
transform 1 0 14536 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1324_
timestamp 1649977179
transform -1 0 15824 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1325_
timestamp 1649977179
transform 1 0 15088 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1326_
timestamp 1649977179
transform 1 0 12788 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1327_
timestamp 1649977179
transform 1 0 13156 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1328_
timestamp 1649977179
transform -1 0 12512 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1329_
timestamp 1649977179
transform 1 0 12880 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1330_
timestamp 1649977179
transform -1 0 16376 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1331_
timestamp 1649977179
transform -1 0 14904 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1332_
timestamp 1649977179
transform 1 0 16652 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1333_
timestamp 1649977179
transform 1 0 15180 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1334_
timestamp 1649977179
transform 1 0 12420 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1335_
timestamp 1649977179
transform 1 0 14076 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1336_
timestamp 1649977179
transform 1 0 12328 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1337_
timestamp 1649977179
transform 1 0 21896 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1338_
timestamp 1649977179
transform 1 0 12880 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1339_
timestamp 1649977179
transform 1 0 14260 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1340_
timestamp 1649977179
transform -1 0 15548 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1341_
timestamp 1649977179
transform 1 0 12420 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1342_
timestamp 1649977179
transform 1 0 13248 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1343_
timestamp 1649977179
transform -1 0 13616 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1344_
timestamp 1649977179
transform 1 0 15456 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1345_
timestamp 1649977179
transform 1 0 15272 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1346_
timestamp 1649977179
transform 1 0 22724 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1347_
timestamp 1649977179
transform -1 0 22816 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1348_
timestamp 1649977179
transform 1 0 25300 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1349_
timestamp 1649977179
transform 1 0 20608 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1350_
timestamp 1649977179
transform -1 0 24656 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1351_
timestamp 1649977179
transform 1 0 26956 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1352_
timestamp 1649977179
transform -1 0 28428 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1353_
timestamp 1649977179
transform 1 0 28060 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1354_
timestamp 1649977179
transform 1 0 21988 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1355_
timestamp 1649977179
transform -1 0 28336 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1356_
timestamp 1649977179
transform 1 0 26956 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1357_
timestamp 1649977179
transform -1 0 27784 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1358_
timestamp 1649977179
transform 1 0 26496 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1359_
timestamp 1649977179
transform -1 0 27692 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1360_
timestamp 1649977179
transform 1 0 25392 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1361_
timestamp 1649977179
transform -1 0 26312 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1362_
timestamp 1649977179
transform 1 0 22540 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1363_
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1364_
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1365_
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1366_
timestamp 1649977179
transform 1 0 19320 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1367_
timestamp 1649977179
transform 1 0 17388 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1368_
timestamp 1649977179
transform -1 0 22172 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1369_
timestamp 1649977179
transform -1 0 19688 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1370_
timestamp 1649977179
transform 1 0 18032 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1371_
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1372_
timestamp 1649977179
transform 1 0 16468 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1373_
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1374_
timestamp 1649977179
transform 1 0 16560 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1375_
timestamp 1649977179
transform 1 0 24380 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1376_
timestamp 1649977179
transform -1 0 23920 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1377_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13064 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1378_
timestamp 1649977179
transform -1 0 18768 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1379_
timestamp 1649977179
transform 1 0 22356 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1380_
timestamp 1649977179
transform -1 0 22080 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1381_
timestamp 1649977179
transform 1 0 20056 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1382_
timestamp 1649977179
transform -1 0 21160 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1383_
timestamp 1649977179
transform -1 0 19596 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1384_
timestamp 1649977179
transform 1 0 18124 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1385_
timestamp 1649977179
transform -1 0 18676 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1386_
timestamp 1649977179
transform 1 0 18032 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1387_
timestamp 1649977179
transform -1 0 18216 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1388_
timestamp 1649977179
transform 1 0 18032 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1389_
timestamp 1649977179
transform 1 0 20516 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1390_
timestamp 1649977179
transform -1 0 20148 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1391_
timestamp 1649977179
transform 1 0 19688 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1392_
timestamp 1649977179
transform -1 0 20424 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1393_
timestamp 1649977179
transform 1 0 19228 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1394_
timestamp 1649977179
transform -1 0 20516 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1395_
timestamp 1649977179
transform -1 0 21712 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1396_
timestamp 1649977179
transform -1 0 20976 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1397_
timestamp 1649977179
transform -1 0 25116 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1398_
timestamp 1649977179
transform 1 0 20424 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1399_
timestamp 1649977179
transform -1 0 25300 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1400_
timestamp 1649977179
transform 1 0 27324 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1401_
timestamp 1649977179
transform -1 0 28060 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1402_
timestamp 1649977179
transform 1 0 26036 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1403_
timestamp 1649977179
transform -1 0 27232 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1404_
timestamp 1649977179
transform 1 0 23092 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1405_
timestamp 1649977179
transform -1 0 23920 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1406_
timestamp 1649977179
transform 1 0 23092 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1407_
timestamp 1649977179
transform 1 0 23276 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1408_
timestamp 1649977179
transform -1 0 20424 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1409_
timestamp 1649977179
transform 1 0 10672 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1410_
timestamp 1649977179
transform -1 0 20608 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1411_
timestamp 1649977179
transform 1 0 19228 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1412_
timestamp 1649977179
transform -1 0 20148 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1413_
timestamp 1649977179
transform -1 0 11040 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1414_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 14536 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1415_
timestamp 1649977179
transform -1 0 10028 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor4b_2  _1416_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 10120 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1417_
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _1418_
timestamp 1649977179
transform -1 0 9384 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _1419_
timestamp 1649977179
transform -1 0 10764 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_2  _1420_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1421_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 9844 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1422_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 36524 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1423_
timestamp 1649977179
transform -1 0 29992 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1424_
timestamp 1649977179
transform 1 0 21712 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1425_
timestamp 1649977179
transform 1 0 5060 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1426_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21988 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1427_
timestamp 1649977179
transform -1 0 17664 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1428_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18952 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1429_
timestamp 1649977179
transform 1 0 23276 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1430_
timestamp 1649977179
transform -1 0 26036 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1431_
timestamp 1649977179
transform -1 0 22540 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1432_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12052 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1433_
timestamp 1649977179
transform -1 0 35512 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1434_
timestamp 1649977179
transform -1 0 31464 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1435_
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1436_
timestamp 1649977179
transform 1 0 4876 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1437_
timestamp 1649977179
transform -1 0 22356 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1438_
timestamp 1649977179
transform -1 0 17480 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1439_
timestamp 1649977179
transform 1 0 19228 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1440_
timestamp 1649977179
transform 1 0 23184 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1441_
timestamp 1649977179
transform -1 0 25668 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1442_
timestamp 1649977179
transform -1 0 21344 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1443_
timestamp 1649977179
transform 1 0 9016 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1444_
timestamp 1649977179
transform 1 0 10212 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1445_
timestamp 1649977179
transform -1 0 7544 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1446_
timestamp 1649977179
transform -1 0 12788 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1447_
timestamp 1649977179
transform -1 0 36064 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1448_
timestamp 1649977179
transform -1 0 31464 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1449_
timestamp 1649977179
transform 1 0 22356 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1450_
timestamp 1649977179
transform 1 0 27324 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1451_
timestamp 1649977179
transform -1 0 27600 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1452_
timestamp 1649977179
transform 1 0 6440 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1453_
timestamp 1649977179
transform -1 0 27416 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1454_
timestamp 1649977179
transform 1 0 15364 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1455_
timestamp 1649977179
transform 1 0 18032 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1456_
timestamp 1649977179
transform 1 0 23276 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1457_
timestamp 1649977179
transform 1 0 25116 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1458_
timestamp 1649977179
transform -1 0 26128 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1459_
timestamp 1649977179
transform -1 0 7820 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1460_
timestamp 1649977179
transform 1 0 13616 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1461_
timestamp 1649977179
transform 1 0 13708 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1462_
timestamp 1649977179
transform 1 0 37260 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1463_
timestamp 1649977179
transform 1 0 35788 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1464_
timestamp 1649977179
transform -1 0 37628 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1465_
timestamp 1649977179
transform 1 0 28796 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1466_
timestamp 1649977179
transform 1 0 28796 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1467_
timestamp 1649977179
transform -1 0 30176 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1468_
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1469_
timestamp 1649977179
transform 1 0 28336 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1470_
timestamp 1649977179
transform 1 0 10488 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1471_
timestamp 1649977179
transform 1 0 10120 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1472_
timestamp 1649977179
transform 1 0 9476 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1473_
timestamp 1649977179
transform 1 0 29348 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1474_
timestamp 1649977179
transform -1 0 13984 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1475_
timestamp 1649977179
transform 1 0 14076 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1476_
timestamp 1649977179
transform 1 0 12512 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1477_
timestamp 1649977179
transform 1 0 16744 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1478_
timestamp 1649977179
transform 1 0 18400 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1479_
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1480_
timestamp 1649977179
transform -1 0 19872 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1481_
timestamp 1649977179
transform -1 0 25760 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1482_
timestamp 1649977179
transform -1 0 18676 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1483_
timestamp 1649977179
transform -1 0 8648 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1484_
timestamp 1649977179
transform -1 0 12236 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1485_
timestamp 1649977179
transform 1 0 11868 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1486_
timestamp 1649977179
transform -1 0 37536 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1487_
timestamp 1649977179
transform -1 0 29072 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1488_
timestamp 1649977179
transform 1 0 27232 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1489_
timestamp 1649977179
transform 1 0 10212 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1490_
timestamp 1649977179
transform 1 0 27968 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1491_
timestamp 1649977179
transform -1 0 17664 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1492_
timestamp 1649977179
transform 1 0 16652 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1493_
timestamp 1649977179
transform 1 0 12972 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1494_
timestamp 1649977179
transform 1 0 16744 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1495_
timestamp 1649977179
transform 1 0 20424 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1496_
timestamp 1649977179
transform 1 0 20516 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1497_
timestamp 1649977179
transform 1 0 18952 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1498_
timestamp 1649977179
transform -1 0 20700 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1499_
timestamp 1649977179
transform -1 0 17664 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1500_
timestamp 1649977179
transform -1 0 8464 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1501_
timestamp 1649977179
transform -1 0 16192 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1502_
timestamp 1649977179
transform -1 0 37812 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1503_
timestamp 1649977179
transform -1 0 30176 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1504_
timestamp 1649977179
transform 1 0 28244 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1505_
timestamp 1649977179
transform 1 0 10120 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1506_
timestamp 1649977179
transform -1 0 29072 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1507_
timestamp 1649977179
transform 1 0 14076 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1508_
timestamp 1649977179
transform 1 0 16744 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1509_
timestamp 1649977179
transform 1 0 18124 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1510_
timestamp 1649977179
transform -1 0 20884 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1511_
timestamp 1649977179
transform -1 0 17664 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1512_
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1513_
timestamp 1649977179
transform -1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1514_
timestamp 1649977179
transform 1 0 12144 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1515_
timestamp 1649977179
transform -1 0 37260 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1516_
timestamp 1649977179
transform -1 0 29808 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1517_
timestamp 1649977179
transform 1 0 28336 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1518_
timestamp 1649977179
transform 1 0 9660 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1519_
timestamp 1649977179
transform 1 0 28888 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1520_
timestamp 1649977179
transform 1 0 13248 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1521_
timestamp 1649977179
transform 1 0 17020 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1522_
timestamp 1649977179
transform 1 0 18860 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1523_
timestamp 1649977179
transform -1 0 21160 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1524_
timestamp 1649977179
transform -1 0 17940 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1525_
timestamp 1649977179
transform -1 0 9936 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1526_
timestamp 1649977179
transform 1 0 17848 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1527_
timestamp 1649977179
transform 1 0 16836 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1528_
timestamp 1649977179
transform -1 0 36432 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1529_
timestamp 1649977179
transform -1 0 30176 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1530_
timestamp 1649977179
transform 1 0 27324 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1531_
timestamp 1649977179
transform 1 0 9936 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1532_
timestamp 1649977179
transform 1 0 27968 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1533_
timestamp 1649977179
transform 1 0 12052 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1534_
timestamp 1649977179
transform 1 0 16652 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1535_
timestamp 1649977179
transform 1 0 18124 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1536_
timestamp 1649977179
transform 1 0 19596 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1537_
timestamp 1649977179
transform -1 0 18032 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1538_
timestamp 1649977179
transform 1 0 17112 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1539_
timestamp 1649977179
transform -1 0 17480 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1540_
timestamp 1649977179
transform -1 0 32752 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1541_
timestamp 1649977179
transform -1 0 28520 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1542_
timestamp 1649977179
transform 1 0 26312 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1543_
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1544_
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1545_
timestamp 1649977179
transform 1 0 15088 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1546_
timestamp 1649977179
transform 1 0 17112 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1547_
timestamp 1649977179
transform 1 0 14996 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1548_
timestamp 1649977179
transform 1 0 19412 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1549_
timestamp 1649977179
transform -1 0 19688 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1550_
timestamp 1649977179
transform 1 0 15640 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1551_
timestamp 1649977179
transform -1 0 16008 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1552_
timestamp 1649977179
transform -1 0 34500 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1553_
timestamp 1649977179
transform -1 0 28428 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1554_
timestamp 1649977179
transform 1 0 23184 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1555_
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1556_
timestamp 1649977179
transform 1 0 23644 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1557_
timestamp 1649977179
transform 1 0 13616 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1558_
timestamp 1649977179
transform 1 0 14628 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1559_
timestamp 1649977179
transform 1 0 14812 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1560_
timestamp 1649977179
transform 1 0 15824 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1561_
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1562_
timestamp 1649977179
transform -1 0 8188 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1563_
timestamp 1649977179
transform 1 0 10304 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1564_
timestamp 1649977179
transform -1 0 31464 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1565_
timestamp 1649977179
transform -1 0 28704 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1566_
timestamp 1649977179
transform 1 0 22908 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1567_
timestamp 1649977179
transform 1 0 11500 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1568_
timestamp 1649977179
transform 1 0 23552 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1569_
timestamp 1649977179
transform 1 0 14904 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1570_
timestamp 1649977179
transform 1 0 16284 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1571_
timestamp 1649977179
transform 1 0 16376 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1572_
timestamp 1649977179
transform -1 0 17756 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1573_
timestamp 1649977179
transform 1 0 17112 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1574_
timestamp 1649977179
transform -1 0 8464 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1575_
timestamp 1649977179
transform 1 0 9108 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1576_
timestamp 1649977179
transform 1 0 18308 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1577_
timestamp 1649977179
transform -1 0 14996 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1578_
timestamp 1649977179
transform -1 0 8188 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1579_
timestamp 1649977179
transform -1 0 6164 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1580_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4784 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1581_
timestamp 1649977179
transform 1 0 2576 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1582_
timestamp 1649977179
transform 1 0 2944 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1583_
timestamp 1649977179
transform 1 0 2760 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1584_
timestamp 1649977179
transform 1 0 2852 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1585_
timestamp 1649977179
transform 1 0 4416 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1586_
timestamp 1649977179
transform -1 0 22540 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1587_
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1588_
timestamp 1649977179
transform -1 0 18124 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1589_
timestamp 1649977179
transform 1 0 4416 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1590_
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1591_
timestamp 1649977179
transform 1 0 4416 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1592_
timestamp 1649977179
transform 1 0 4048 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1593_
timestamp 1649977179
transform -1 0 4324 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1594_
timestamp 1649977179
transform 1 0 4048 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1595_
timestamp 1649977179
transform 1 0 5428 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1596_
timestamp 1649977179
transform -1 0 4324 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1597_
timestamp 1649977179
transform 1 0 4416 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1598_
timestamp 1649977179
transform 1 0 3772 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1599_
timestamp 1649977179
transform 1 0 3772 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1600_
timestamp 1649977179
transform 1 0 2852 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1601_
timestamp 1649977179
transform 1 0 4416 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1602_
timestamp 1649977179
transform 1 0 2944 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1603_
timestamp 1649977179
transform 1 0 3404 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1604_
timestamp 1649977179
transform 1 0 2760 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1605_
timestamp 1649977179
transform 1 0 5428 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1606_
timestamp 1649977179
transform 1 0 2668 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1607_
timestamp 1649977179
transform 1 0 3128 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1608_
timestamp 1649977179
transform 1 0 2576 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1609_
timestamp 1649977179
transform 1 0 3772 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1610_
timestamp 1649977179
transform 1 0 3128 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1611_
timestamp 1649977179
transform 1 0 3128 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1612_
timestamp 1649977179
transform 1 0 5060 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1613_
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1614_
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1615_
timestamp 1649977179
transform -1 0 7820 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1616_
timestamp 1649977179
transform 1 0 8280 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1617_
timestamp 1649977179
transform 1 0 8924 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1618_
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1619_
timestamp 1649977179
transform 1 0 8004 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1620_
timestamp 1649977179
transform 1 0 5612 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1621_
timestamp 1649977179
transform -1 0 6624 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1622_
timestamp 1649977179
transform 1 0 8372 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1623_
timestamp 1649977179
transform 1 0 9384 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1624_
timestamp 1649977179
transform 1 0 7728 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1625_
timestamp 1649977179
transform 1 0 6716 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1626_
timestamp 1649977179
transform 1 0 9568 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1627_
timestamp 1649977179
transform 1 0 9936 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1628_
timestamp 1649977179
transform 1 0 7544 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1629_
timestamp 1649977179
transform 1 0 8924 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1630_
timestamp 1649977179
transform 1 0 5336 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1631_
timestamp 1649977179
transform 1 0 9568 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1632_
timestamp 1649977179
transform 1 0 9384 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1633_
timestamp 1649977179
transform 1 0 9752 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1634_
timestamp 1649977179
transform 1 0 6624 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1635_
timestamp 1649977179
transform 1 0 7636 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1636_
timestamp 1649977179
transform 1 0 9568 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1637_
timestamp 1649977179
transform 1 0 12420 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1638_
timestamp 1649977179
transform 1 0 12420 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1639_
timestamp 1649977179
transform 1 0 9200 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1640_
timestamp 1649977179
transform 1 0 10948 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1641_
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1642_
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1643_
timestamp 1649977179
transform 1 0 12512 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1644_
timestamp 1649977179
transform 1 0 10580 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1645_
timestamp 1649977179
transform 1 0 12696 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1646_
timestamp 1649977179
transform -1 0 23552 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1647_
timestamp 1649977179
transform -1 0 23920 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1648_
timestamp 1649977179
transform 1 0 26220 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1649_
timestamp 1649977179
transform 1 0 26496 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1650_
timestamp 1649977179
transform 1 0 26036 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1651_
timestamp 1649977179
transform -1 0 31188 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1652_
timestamp 1649977179
transform -1 0 31648 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1653_
timestamp 1649977179
transform -1 0 31280 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1654_
timestamp 1649977179
transform -1 0 28520 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1655_
timestamp 1649977179
transform 1 0 22264 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1656_
timestamp 1649977179
transform 1 0 22080 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1657_
timestamp 1649977179
transform -1 0 38088 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1658_
timestamp 1649977179
transform -1 0 36800 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1659_
timestamp 1649977179
transform -1 0 34224 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1660_
timestamp 1649977179
transform -1 0 37076 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1661_
timestamp 1649977179
transform -1 0 34776 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1662_
timestamp 1649977179
transform -1 0 25852 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1663_
timestamp 1649977179
transform -1 0 27968 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1664_
timestamp 1649977179
transform -1 0 24380 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1665_
timestamp 1649977179
transform -1 0 28428 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1666_
timestamp 1649977179
transform 1 0 30176 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1667_
timestamp 1649977179
transform -1 0 32384 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1668_
timestamp 1649977179
transform -1 0 40388 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1669_
timestamp 1649977179
transform -1 0 40664 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1670_
timestamp 1649977179
transform -1 0 41308 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1671_
timestamp 1649977179
transform -1 0 40572 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1672_
timestamp 1649977179
transform -1 0 40572 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1673_
timestamp 1649977179
transform 1 0 38916 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1674_
timestamp 1649977179
transform -1 0 38824 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1675_
timestamp 1649977179
transform 1 0 35328 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1676_
timestamp 1649977179
transform -1 0 33212 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1677_
timestamp 1649977179
transform 1 0 33488 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1678_
timestamp 1649977179
transform 1 0 29808 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1679_
timestamp 1649977179
transform -1 0 36708 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1680_
timestamp 1649977179
transform -1 0 35512 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1681_
timestamp 1649977179
transform -1 0 41308 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1682_
timestamp 1649977179
transform -1 0 41308 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1683_
timestamp 1649977179
transform 1 0 39008 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1684_
timestamp 1649977179
transform 1 0 39836 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1685_
timestamp 1649977179
transform 1 0 39836 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1686_
timestamp 1649977179
transform 1 0 35328 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1687_
timestamp 1649977179
transform 1 0 31188 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1688_
timestamp 1649977179
transform 1 0 32016 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1689_
timestamp 1649977179
transform -1 0 33028 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1690_
timestamp 1649977179
transform 1 0 35328 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1691_
timestamp 1649977179
transform 1 0 38180 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1692_
timestamp 1649977179
transform 1 0 39100 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1693_
timestamp 1649977179
transform 1 0 39008 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1694_
timestamp 1649977179
transform 1 0 39192 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1695_
timestamp 1649977179
transform -1 0 36708 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1696_
timestamp 1649977179
transform -1 0 34224 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1697_
timestamp 1649977179
transform -1 0 31648 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1698_
timestamp 1649977179
transform -1 0 34500 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1699_
timestamp 1649977179
transform -1 0 32016 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1700_
timestamp 1649977179
transform -1 0 34500 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1701_
timestamp 1649977179
transform -1 0 23920 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1702_
timestamp 1649977179
transform -1 0 26128 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1703_
timestamp 1649977179
transform 1 0 25760 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1704_
timestamp 1649977179
transform -1 0 27048 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1705_
timestamp 1649977179
transform -1 0 25208 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1706_
timestamp 1649977179
transform -1 0 22816 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1707_
timestamp 1649977179
transform -1 0 20148 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1708_
timestamp 1649977179
transform 1 0 16836 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1709_
timestamp 1649977179
transform -1 0 15548 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1710_
timestamp 1649977179
transform -1 0 15548 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1711_
timestamp 1649977179
transform -1 0 24656 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1712_
timestamp 1649977179
transform 1 0 28520 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1713_
timestamp 1649977179
transform -1 0 33488 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1714_
timestamp 1649977179
transform 1 0 30360 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1715_
timestamp 1649977179
transform -1 0 34040 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1716_
timestamp 1649977179
transform 1 0 31556 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1717_
timestamp 1649977179
transform 1 0 30912 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1718_
timestamp 1649977179
transform -1 0 33580 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1719_
timestamp 1649977179
transform 1 0 29072 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1720_
timestamp 1649977179
transform 1 0 26956 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1721_
timestamp 1649977179
transform 1 0 26772 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1722_
timestamp 1649977179
transform 1 0 27600 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1723_
timestamp 1649977179
transform -1 0 24104 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1724_
timestamp 1649977179
transform -1 0 22816 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1725_
timestamp 1649977179
transform -1 0 25944 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1726_
timestamp 1649977179
transform -1 0 21528 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1727_
timestamp 1649977179
transform -1 0 23460 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1728_
timestamp 1649977179
transform -1 0 22816 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1729_
timestamp 1649977179
transform -1 0 22080 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1730_
timestamp 1649977179
transform 1 0 20516 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1731_
timestamp 1649977179
transform -1 0 20056 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1732_
timestamp 1649977179
transform -1 0 18124 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1733_
timestamp 1649977179
transform -1 0 18676 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1734_
timestamp 1649977179
transform -1 0 20976 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1735_
timestamp 1649977179
transform 1 0 16376 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1736_
timestamp 1649977179
transform 1 0 14076 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1737_
timestamp 1649977179
transform 1 0 11408 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1738_
timestamp 1649977179
transform -1 0 12972 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1739_
timestamp 1649977179
transform 1 0 11776 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1740_
timestamp 1649977179
transform 1 0 11040 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1741_
timestamp 1649977179
transform -1 0 11868 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1742_
timestamp 1649977179
transform -1 0 16192 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1743_
timestamp 1649977179
transform 1 0 11592 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1744_
timestamp 1649977179
transform -1 0 15548 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1745_
timestamp 1649977179
transform -1 0 27048 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1746_
timestamp 1649977179
transform -1 0 30728 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1747_
timestamp 1649977179
transform -1 0 29624 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1748_
timestamp 1649977179
transform -1 0 29072 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1749_
timestamp 1649977179
transform -1 0 28428 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1750_
timestamp 1649977179
transform -1 0 24472 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1751_
timestamp 1649977179
transform -1 0 23644 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1752_
timestamp 1649977179
transform 1 0 17296 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1753_
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1754_
timestamp 1649977179
transform 1 0 14536 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1755_
timestamp 1649977179
transform -1 0 26036 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1756_
timestamp 1649977179
transform 1 0 16376 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1757_
timestamp 1649977179
transform 1 0 18032 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1758_
timestamp 1649977179
transform 1 0 19872 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1759_
timestamp 1649977179
transform 1 0 19872 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1760_
timestamp 1649977179
transform 1 0 20976 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1761_
timestamp 1649977179
transform 1 0 25760 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1762_
timestamp 1649977179
transform -1 0 31004 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1763_
timestamp 1649977179
transform -1 0 29072 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1764_
timestamp 1649977179
transform 1 0 24288 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1765_
timestamp 1649977179
transform 1 0 22080 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1766_
timestamp 1649977179
transform 1 0 20516 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1767_
timestamp 1649977179
transform 1 0 20516 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1768_
timestamp 1649977179
transform -1 0 13616 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1769_
timestamp 1649977179
transform -1 0 11592 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1770_
timestamp 1649977179
transform -1 0 15824 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1771_
timestamp 1649977179
transform -1 0 12972 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1772_
timestamp 1649977179
transform -1 0 17020 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1773_
timestamp 1649977179
transform -1 0 14812 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1774_
timestamp 1649977179
transform -1 0 18952 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1775_
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1776_
timestamp 1649977179
transform 1 0 13340 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1777_
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1778_
timestamp 1649977179
transform 1 0 12144 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1779_
timestamp 1649977179
transform -1 0 16008 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1780_
timestamp 1649977179
transform -1 0 9936 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21896 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_wb_clk_i
timestamp 1649977179
transform -1 0 12236 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_wb_clk_i
timestamp 1649977179
transform 1 0 28612 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_0_wb_clk_i
timestamp 1649977179
transform 1 0 6716 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_1_wb_clk_i
timestamp 1649977179
transform 1 0 14352 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_2_wb_clk_i
timestamp 1649977179
transform 1 0 11776 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_3_wb_clk_i
timestamp 1649977179
transform 1 0 4416 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_4_wb_clk_i
timestamp 1649977179
transform 1 0 6716 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_5_wb_clk_i
timestamp 1649977179
transform -1 0 9384 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_6_wb_clk_i
timestamp 1649977179
transform 1 0 14444 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_7_wb_clk_i
timestamp 1649977179
transform 1 0 19504 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_8_wb_clk_i
timestamp 1649977179
transform 1 0 25484 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_9_wb_clk_i
timestamp 1649977179
transform -1 0 29164 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_10_wb_clk_i
timestamp 1649977179
transform 1 0 36340 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_11_wb_clk_i
timestamp 1649977179
transform 1 0 36340 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_12_wb_clk_i
timestamp 1649977179
transform 1 0 29256 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_13_wb_clk_i
timestamp 1649977179
transform 1 0 26772 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_14_wb_clk_i
timestamp 1649977179
transform -1 0 36892 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_15_wb_clk_i
timestamp 1649977179
transform 1 0 40204 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_16_wb_clk_i
timestamp 1649977179
transform 1 0 38732 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_17_wb_clk_i
timestamp 1649977179
transform -1 0 34224 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_18_wb_clk_i
timestamp 1649977179
transform -1 0 25944 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_19_wb_clk_i
timestamp 1649977179
transform 1 0 25760 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_20_wb_clk_i
timestamp 1649977179
transform 1 0 18492 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_21_wb_clk_i
timestamp 1649977179
transform 1 0 17020 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_22_wb_clk_i
timestamp 1649977179
transform -1 0 11776 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_23_wb_clk_i
timestamp 1649977179
transform 1 0 4140 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_24_wb_clk_i
timestamp 1649977179
transform 1 0 6716 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform -1 0 2024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform -1 0 5888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform -1 0 18584 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform -1 0 4508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform -1 0 18124 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform -1 0 18768 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1649977179
transform -1 0 6716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform -1 0 8464 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform -1 0 5152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform -1 0 10396 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform -1 0 7360 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform -1 0 2668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input15 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 10120 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input16
timestamp 1649977179
transform -1 0 15272 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform -1 0 13892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input18
timestamp 1649977179
transform -1 0 11040 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input19
timestamp 1649977179
transform -1 0 11040 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input20
timestamp 1649977179
transform 1 0 14444 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input21
timestamp 1649977179
transform 1 0 12788 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input22
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1649977179
transform -1 0 17756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1649977179
transform -1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1649977179
transform -1 0 16008 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input26
timestamp 1649977179
transform -1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1649977179
transform 1 0 10764 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform -1 0 5244 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1649977179
transform -1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1649977179
transform -1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1649977179
transform -1 0 11040 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1649977179
transform 1 0 15732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1649977179
transform -1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1649977179
transform -1 0 6992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1649977179
transform -1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1649977179
transform -1 0 7728 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1649977179
transform -1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1649977179
transform 1 0 18124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1649977179
transform -1 0 16744 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1649977179
transform -1 0 17020 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1649977179
transform -1 0 15272 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1649977179
transform 1 0 15456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_43 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 45264 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_44
timestamp 1649977179
transform -1 0 55568 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_45
timestamp 1649977179
transform -1 0 65136 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_46
timestamp 1649977179
transform -1 0 25392 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_47
timestamp 1649977179
transform -1 0 35328 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_48
timestamp 1649977179
transform -1 0 5520 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_49
timestamp 1649977179
transform -1 0 15456 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_50
timestamp 1649977179
transform 1 0 67896 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_51
timestamp 1649977179
transform 1 0 67436 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_52
timestamp 1649977179
transform 1 0 66792 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_53
timestamp 1649977179
transform 1 0 67436 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_54
timestamp 1649977179
transform -1 0 58788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_55
timestamp 1649977179
transform -1 0 58144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_56
timestamp 1649977179
transform -1 0 56488 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_57
timestamp 1649977179
transform -1 0 57500 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_58
timestamp 1649977179
transform -1 0 57132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_59
timestamp 1649977179
transform -1 0 59432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_60
timestamp 1649977179
transform -1 0 58144 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_61
timestamp 1649977179
transform -1 0 58788 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_62
timestamp 1649977179
transform -1 0 58788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_63
timestamp 1649977179
transform -1 0 59432 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_64
timestamp 1649977179
transform -1 0 60720 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_65
timestamp 1649977179
transform -1 0 58144 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_66
timestamp 1649977179
transform -1 0 60076 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_67
timestamp 1649977179
transform -1 0 57500 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_68
timestamp 1649977179
transform -1 0 58144 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_69
timestamp 1649977179
transform -1 0 59432 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_70
timestamp 1649977179
transform -1 0 61364 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_71
timestamp 1649977179
transform -1 0 58788 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_72
timestamp 1649977179
transform -1 0 58788 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_73
timestamp 1649977179
transform -1 0 60720 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_74
timestamp 1649977179
transform -1 0 59432 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_75
timestamp 1649977179
transform -1 0 60720 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_76
timestamp 1649977179
transform -1 0 60076 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_77
timestamp 1649977179
transform -1 0 62008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_78
timestamp 1649977179
transform -1 0 61364 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_79
timestamp 1649977179
transform -1 0 59432 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_80
timestamp 1649977179
transform -1 0 61364 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_81
timestamp 1649977179
transform -1 0 62008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_82
timestamp 1649977179
transform -1 0 63296 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_83
timestamp 1649977179
transform -1 0 60720 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_84
timestamp 1649977179
transform -1 0 59064 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_85
timestamp 1649977179
transform -1 0 59708 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_86
timestamp 1649977179
transform -1 0 60720 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_87
timestamp 1649977179
transform -1 0 62008 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_88
timestamp 1649977179
transform -1 0 63940 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_89
timestamp 1649977179
transform -1 0 61364 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_90
timestamp 1649977179
transform -1 0 60352 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_91
timestamp 1649977179
transform -1 0 63296 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_92
timestamp 1649977179
transform 1 0 67436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_93
timestamp 1649977179
transform 1 0 66792 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_94
timestamp 1649977179
transform 1 0 67896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_95
timestamp 1649977179
transform 1 0 67436 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_96
timestamp 1649977179
transform 1 0 67436 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_97
timestamp 1649977179
transform 1 0 67896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_98
timestamp 1649977179
transform 1 0 67896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_99
timestamp 1649977179
transform 1 0 67436 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_100
timestamp 1649977179
transform 1 0 67436 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_101
timestamp 1649977179
transform 1 0 67896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_102
timestamp 1649977179
transform 1 0 67896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_103
timestamp 1649977179
transform 1 0 67436 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_104
timestamp 1649977179
transform 1 0 67436 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_105
timestamp 1649977179
transform 1 0 67896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_106
timestamp 1649977179
transform 1 0 67896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_107
timestamp 1649977179
transform 1 0 67436 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_108
timestamp 1649977179
transform 1 0 67436 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_109
timestamp 1649977179
transform 1 0 67896 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_110
timestamp 1649977179
transform 1 0 67896 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_111
timestamp 1649977179
transform 1 0 67436 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_112
timestamp 1649977179
transform 1 0 67436 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_113
timestamp 1649977179
transform 1 0 67896 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_114
timestamp 1649977179
transform 1 0 67896 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_115
timestamp 1649977179
transform 1 0 67436 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_116
timestamp 1649977179
transform 1 0 67436 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_117
timestamp 1649977179
transform 1 0 67896 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_118
timestamp 1649977179
transform 1 0 67896 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_119
timestamp 1649977179
transform 1 0 67436 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_120
timestamp 1649977179
transform 1 0 67436 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_121
timestamp 1649977179
transform 1 0 67896 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_122
timestamp 1649977179
transform 1 0 67896 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_123
timestamp 1649977179
transform 1 0 67436 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_124
timestamp 1649977179
transform 1 0 67436 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_125
timestamp 1649977179
transform 1 0 67896 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_126
timestamp 1649977179
transform 1 0 67896 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_127
timestamp 1649977179
transform 1 0 67436 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_128
timestamp 1649977179
transform 1 0 67436 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_129
timestamp 1649977179
transform 1 0 67896 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_130
timestamp 1649977179
transform -1 0 56856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_131
timestamp 1649977179
transform -1 0 56856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_132
timestamp 1649977179
transform -1 0 58144 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_133
timestamp 1649977179
transform -1 0 20792 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_134
timestamp 1649977179
transform 1 0 19780 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_135
timestamp 1649977179
transform -1 0 21344 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_136
timestamp 1649977179
transform 1 0 20424 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_137
timestamp 1649977179
transform 1 0 19780 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_138
timestamp 1649977179
transform 1 0 21068 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_139
timestamp 1649977179
transform 1 0 20424 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_140
timestamp 1649977179
transform -1 0 22724 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_141
timestamp 1649977179
transform 1 0 21804 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_142
timestamp 1649977179
transform 1 0 21068 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_143
timestamp 1649977179
transform 1 0 22448 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_144
timestamp 1649977179
transform 1 0 22356 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_145
timestamp 1649977179
transform 1 0 23000 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_146
timestamp 1649977179
transform 1 0 22356 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_147
timestamp 1649977179
transform 1 0 23644 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_148
timestamp 1649977179
transform 1 0 23000 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_149
timestamp 1649977179
transform 1 0 24564 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_150
timestamp 1649977179
transform 1 0 24288 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_151
timestamp 1649977179
transform 1 0 23644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_152
timestamp 1649977179
transform 1 0 25208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_153
timestamp 1649977179
transform 1 0 24932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_154
timestamp 1649977179
transform 1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_155
timestamp 1649977179
transform 1 0 24932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_156
timestamp 1649977179
transform 1 0 25576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_157
timestamp 1649977179
transform 1 0 26220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_158
timestamp 1649977179
transform 1 0 25576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_159
timestamp 1649977179
transform 1 0 26220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_160
timestamp 1649977179
transform -1 0 28244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_161
timestamp 1649977179
transform 1 0 27508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_162
timestamp 1649977179
transform 1 0 27508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_163
timestamp 1649977179
transform -1 0 29072 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_164
timestamp 1649977179
transform 1 0 28152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_165
timestamp 1649977179
transform 1 0 28796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_166
timestamp 1649977179
transform -1 0 29900 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_167
timestamp 1649977179
transform 1 0 28152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_168
timestamp 1649977179
transform 1 0 29440 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_169
timestamp 1649977179
transform 1 0 28796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_170
timestamp 1649977179
transform 1 0 30452 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_171
timestamp 1649977179
transform 1 0 30084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_172
timestamp 1649977179
transform -1 0 31372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_173
timestamp 1649977179
transform 1 0 30728 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_174
timestamp 1649977179
transform 1 0 30084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_175
timestamp 1649977179
transform 1 0 31372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_176
timestamp 1649977179
transform 1 0 30728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_177
timestamp 1649977179
transform -1 0 32936 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_178
timestamp 1649977179
transform 1 0 31372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_179
timestamp 1649977179
transform 1 0 32660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_180
timestamp 1649977179
transform 1 0 32660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_181
timestamp 1649977179
transform 1 0 33304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_182
timestamp 1649977179
transform 1 0 33304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_183
timestamp 1649977179
transform 1 0 33948 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_184
timestamp 1649977179
transform -1 0 34868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_185
timestamp 1649977179
transform 1 0 33948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_186
timestamp 1649977179
transform 1 0 34684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_187
timestamp 1649977179
transform -1 0 35696 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_188
timestamp 1649977179
transform 1 0 35328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_189
timestamp 1649977179
transform -1 0 36248 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_190
timestamp 1649977179
transform -1 0 36524 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_191
timestamp 1649977179
transform -1 0 37536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_192
timestamp 1649977179
transform -1 0 37536 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_193
timestamp 1649977179
transform -1 0 38180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_194
timestamp 1649977179
transform -1 0 38180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_195
timestamp 1649977179
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_196
timestamp 1649977179
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_197
timestamp 1649977179
transform -1 0 40112 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_198
timestamp 1649977179
transform -1 0 39468 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_199
timestamp 1649977179
transform -1 0 40756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_200
timestamp 1649977179
transform -1 0 40112 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_201
timestamp 1649977179
transform -1 0 40112 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_202
timestamp 1649977179
transform -1 0 41400 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_203
timestamp 1649977179
transform -1 0 40756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_204
timestamp 1649977179
transform -1 0 40756 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_205
timestamp 1649977179
transform -1 0 41400 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_206
timestamp 1649977179
transform -1 0 42688 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_207
timestamp 1649977179
transform -1 0 41400 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_208
timestamp 1649977179
transform -1 0 42044 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_209
timestamp 1649977179
transform -1 0 43332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_210
timestamp 1649977179
transform -1 0 42688 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_211
timestamp 1649977179
transform -1 0 43976 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_212
timestamp 1649977179
transform -1 0 43332 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_213
timestamp 1649977179
transform -1 0 42872 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_214
timestamp 1649977179
transform -1 0 43976 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_215
timestamp 1649977179
transform -1 0 43516 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_216
timestamp 1649977179
transform -1 0 45264 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_217
timestamp 1649977179
transform -1 0 44620 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_218
timestamp 1649977179
transform -1 0 45908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_219
timestamp 1649977179
transform -1 0 45264 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_220
timestamp 1649977179
transform -1 0 46552 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_221
timestamp 1649977179
transform -1 0 45908 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_222
timestamp 1649977179
transform -1 0 45356 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_223
timestamp 1649977179
transform -1 0 46000 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_224
timestamp 1649977179
transform -1 0 46552 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_225
timestamp 1649977179
transform -1 0 47840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_226
timestamp 1649977179
transform -1 0 46644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_227
timestamp 1649977179
transform -1 0 48484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_228
timestamp 1649977179
transform -1 0 47840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_229
timestamp 1649977179
transform -1 0 47288 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_230
timestamp 1649977179
transform -1 0 49128 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_231
timestamp 1649977179
transform -1 0 48484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_232
timestamp 1649977179
transform -1 0 48116 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_233
timestamp 1649977179
transform -1 0 49128 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_234
timestamp 1649977179
transform -1 0 50416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_235
timestamp 1649977179
transform -1 0 49772 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_236
timestamp 1649977179
transform -1 0 49220 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_237
timestamp 1649977179
transform -1 0 51060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_238
timestamp 1649977179
transform -1 0 50416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_239
timestamp 1649977179
transform -1 0 51704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_240
timestamp 1649977179
transform -1 0 51060 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_241
timestamp 1649977179
transform -1 0 50600 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_242
timestamp 1649977179
transform -1 0 51704 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_243
timestamp 1649977179
transform -1 0 51244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_244
timestamp 1649977179
transform -1 0 52992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_245
timestamp 1649977179
transform -1 0 51888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_246
timestamp 1649977179
transform -1 0 53636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_247
timestamp 1649977179
transform -1 0 52992 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_248
timestamp 1649977179
transform -1 0 54280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_249
timestamp 1649977179
transform -1 0 53636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_250
timestamp 1649977179
transform -1 0 53084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_251
timestamp 1649977179
transform -1 0 53728 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_252
timestamp 1649977179
transform -1 0 54280 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_253
timestamp 1649977179
transform -1 0 55568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_254
timestamp 1649977179
transform -1 0 54924 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_255
timestamp 1649977179
transform -1 0 56212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_256
timestamp 1649977179
transform -1 0 55568 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_257
timestamp 1649977179
transform -1 0 55568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_258
timestamp 1649977179
transform -1 0 56856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_259
timestamp 1649977179
transform -1 0 56212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_260
timestamp 1649977179
transform -1 0 56212 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_261
timestamp 1649977179
transform 1 0 67436 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_262
timestamp 1649977179
transform 1 0 67896 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_263
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_264
timestamp 1649977179
transform -1 0 15640 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_265
timestamp 1649977179
transform 1 0 14352 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_266
timestamp 1649977179
transform 1 0 14996 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_267
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_268
timestamp 1649977179
transform 1 0 15640 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_269
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_270
timestamp 1649977179
transform 1 0 14352 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_271
timestamp 1649977179
transform 1 0 13340 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_272
timestamp 1649977179
transform -1 0 17848 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_273
timestamp 1649977179
transform 1 0 12696 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_274
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_275
timestamp 1649977179
transform 1 0 18032 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_276
timestamp 1649977179
transform -1 0 20332 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_277
timestamp 1649977179
transform 1 0 17112 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_278
timestamp 1649977179
transform 1 0 16652 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_279
timestamp 1649977179
transform 1 0 17296 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_280
timestamp 1649977179
transform -1 0 22080 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_281
timestamp 1649977179
transform 1 0 18492 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_282
timestamp 1649977179
transform 1 0 19136 0 -1 3264
box -38 -48 314 592
<< labels >>
flabel metal2 s 44914 59200 44970 60000 0 FreeSans 224 90 0 0 Sh
port 0 nsew signal tristate
flabel metal2 s 54850 59200 54906 60000 0 FreeSans 224 90 0 0 Sh_cmp
port 1 nsew signal tristate
flabel metal2 s 64786 59200 64842 60000 0 FreeSans 224 90 0 0 Sh_rst
port 2 nsew signal tristate
flabel metal2 s 25042 59200 25098 60000 0 FreeSans 224 90 0 0 Sw1
port 3 nsew signal tristate
flabel metal2 s 34978 59200 35034 60000 0 FreeSans 224 90 0 0 Sw2
port 4 nsew signal tristate
flabel metal2 s 5170 59200 5226 60000 0 FreeSans 224 90 0 0 Vd1
port 5 nsew signal tristate
flabel metal2 s 15106 59200 15162 60000 0 FreeSans 224 90 0 0 Vd2
port 6 nsew signal tristate
flabel metal3 s 69200 52368 70000 52488 0 FreeSans 480 0 0 0 clk_o
port 7 nsew signal tristate
flabel metal3 s 69200 59168 70000 59288 0 FreeSans 480 0 0 0 counter_rst
port 8 nsew signal tristate
flabel metal3 s 69200 57808 70000 57928 0 FreeSans 480 0 0 0 data_o
port 9 nsew signal tristate
flabel metal3 s 69200 55088 70000 55208 0 FreeSans 480 0 0 0 done_o
port 10 nsew signal tristate
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 io_in[0]
port 11 nsew signal input
flabel metal3 s 0 17144 800 17264 0 FreeSans 480 0 0 0 io_in[10]
port 12 nsew signal input
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 io_in[11]
port 13 nsew signal input
flabel metal3 s 0 20136 800 20256 0 FreeSans 480 0 0 0 io_in[12]
port 14 nsew signal input
flabel metal3 s 0 21632 800 21752 0 FreeSans 480 0 0 0 io_in[13]
port 15 nsew signal input
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 io_in[14]
port 16 nsew signal input
flabel metal3 s 0 24624 800 24744 0 FreeSans 480 0 0 0 io_in[15]
port 17 nsew signal input
flabel metal3 s 0 26120 800 26240 0 FreeSans 480 0 0 0 io_in[16]
port 18 nsew signal input
flabel metal3 s 0 27616 800 27736 0 FreeSans 480 0 0 0 io_in[17]
port 19 nsew signal input
flabel metal3 s 0 29112 800 29232 0 FreeSans 480 0 0 0 io_in[18]
port 20 nsew signal input
flabel metal3 s 0 30608 800 30728 0 FreeSans 480 0 0 0 io_in[19]
port 21 nsew signal input
flabel metal3 s 0 3680 800 3800 0 FreeSans 480 0 0 0 io_in[1]
port 22 nsew signal input
flabel metal3 s 0 32104 800 32224 0 FreeSans 480 0 0 0 io_in[20]
port 23 nsew signal input
flabel metal3 s 0 33600 800 33720 0 FreeSans 480 0 0 0 io_in[21]
port 24 nsew signal input
flabel metal3 s 0 35096 800 35216 0 FreeSans 480 0 0 0 io_in[22]
port 25 nsew signal input
flabel metal3 s 0 36592 800 36712 0 FreeSans 480 0 0 0 io_in[23]
port 26 nsew signal input
flabel metal3 s 0 38088 800 38208 0 FreeSans 480 0 0 0 io_in[24]
port 27 nsew signal input
flabel metal3 s 0 39584 800 39704 0 FreeSans 480 0 0 0 io_in[25]
port 28 nsew signal input
flabel metal3 s 0 41080 800 41200 0 FreeSans 480 0 0 0 io_in[26]
port 29 nsew signal input
flabel metal3 s 0 42576 800 42696 0 FreeSans 480 0 0 0 io_in[27]
port 30 nsew signal input
flabel metal3 s 0 44072 800 44192 0 FreeSans 480 0 0 0 io_in[28]
port 31 nsew signal input
flabel metal3 s 0 45568 800 45688 0 FreeSans 480 0 0 0 io_in[29]
port 32 nsew signal input
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 io_in[2]
port 33 nsew signal input
flabel metal3 s 0 47064 800 47184 0 FreeSans 480 0 0 0 io_in[30]
port 34 nsew signal input
flabel metal3 s 0 48560 800 48680 0 FreeSans 480 0 0 0 io_in[31]
port 35 nsew signal input
flabel metal3 s 0 50056 800 50176 0 FreeSans 480 0 0 0 io_in[32]
port 36 nsew signal input
flabel metal3 s 0 51552 800 51672 0 FreeSans 480 0 0 0 io_in[33]
port 37 nsew signal input
flabel metal3 s 0 53048 800 53168 0 FreeSans 480 0 0 0 io_in[34]
port 38 nsew signal input
flabel metal3 s 0 54544 800 54664 0 FreeSans 480 0 0 0 io_in[35]
port 39 nsew signal input
flabel metal3 s 0 56040 800 56160 0 FreeSans 480 0 0 0 io_in[36]
port 40 nsew signal input
flabel metal3 s 0 57536 800 57656 0 FreeSans 480 0 0 0 io_in[37]
port 41 nsew signal input
flabel metal3 s 0 6672 800 6792 0 FreeSans 480 0 0 0 io_in[3]
port 42 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 io_in[4]
port 43 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 io_in[5]
port 44 nsew signal input
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 io_in[6]
port 45 nsew signal input
flabel metal3 s 0 12656 800 12776 0 FreeSans 480 0 0 0 io_in[7]
port 46 nsew signal input
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 io_in[8]
port 47 nsew signal input
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 io_in[9]
port 48 nsew signal input
flabel metal2 s 55954 0 56010 800 0 FreeSans 224 90 0 0 io_oeb[0]
port 49 nsew signal tristate
flabel metal2 s 56874 0 56930 800 0 FreeSans 224 90 0 0 io_oeb[10]
port 50 nsew signal tristate
flabel metal2 s 56966 0 57022 800 0 FreeSans 224 90 0 0 io_oeb[11]
port 51 nsew signal tristate
flabel metal2 s 57058 0 57114 800 0 FreeSans 224 90 0 0 io_oeb[12]
port 52 nsew signal tristate
flabel metal2 s 57150 0 57206 800 0 FreeSans 224 90 0 0 io_oeb[13]
port 53 nsew signal tristate
flabel metal2 s 57242 0 57298 800 0 FreeSans 224 90 0 0 io_oeb[14]
port 54 nsew signal tristate
flabel metal2 s 57334 0 57390 800 0 FreeSans 224 90 0 0 io_oeb[15]
port 55 nsew signal tristate
flabel metal2 s 57426 0 57482 800 0 FreeSans 224 90 0 0 io_oeb[16]
port 56 nsew signal tristate
flabel metal2 s 57518 0 57574 800 0 FreeSans 224 90 0 0 io_oeb[17]
port 57 nsew signal tristate
flabel metal2 s 57610 0 57666 800 0 FreeSans 224 90 0 0 io_oeb[18]
port 58 nsew signal tristate
flabel metal2 s 57702 0 57758 800 0 FreeSans 224 90 0 0 io_oeb[19]
port 59 nsew signal tristate
flabel metal2 s 56046 0 56102 800 0 FreeSans 224 90 0 0 io_oeb[1]
port 60 nsew signal tristate
flabel metal2 s 57794 0 57850 800 0 FreeSans 224 90 0 0 io_oeb[20]
port 61 nsew signal tristate
flabel metal2 s 57886 0 57942 800 0 FreeSans 224 90 0 0 io_oeb[21]
port 62 nsew signal tristate
flabel metal2 s 57978 0 58034 800 0 FreeSans 224 90 0 0 io_oeb[22]
port 63 nsew signal tristate
flabel metal2 s 58070 0 58126 800 0 FreeSans 224 90 0 0 io_oeb[23]
port 64 nsew signal tristate
flabel metal2 s 58162 0 58218 800 0 FreeSans 224 90 0 0 io_oeb[24]
port 65 nsew signal tristate
flabel metal2 s 58254 0 58310 800 0 FreeSans 224 90 0 0 io_oeb[25]
port 66 nsew signal tristate
flabel metal2 s 58346 0 58402 800 0 FreeSans 224 90 0 0 io_oeb[26]
port 67 nsew signal tristate
flabel metal2 s 58438 0 58494 800 0 FreeSans 224 90 0 0 io_oeb[27]
port 68 nsew signal tristate
flabel metal2 s 58530 0 58586 800 0 FreeSans 224 90 0 0 io_oeb[28]
port 69 nsew signal tristate
flabel metal2 s 58622 0 58678 800 0 FreeSans 224 90 0 0 io_oeb[29]
port 70 nsew signal tristate
flabel metal2 s 56138 0 56194 800 0 FreeSans 224 90 0 0 io_oeb[2]
port 71 nsew signal tristate
flabel metal2 s 58714 0 58770 800 0 FreeSans 224 90 0 0 io_oeb[30]
port 72 nsew signal tristate
flabel metal2 s 58806 0 58862 800 0 FreeSans 224 90 0 0 io_oeb[31]
port 73 nsew signal tristate
flabel metal2 s 58898 0 58954 800 0 FreeSans 224 90 0 0 io_oeb[32]
port 74 nsew signal tristate
flabel metal2 s 58990 0 59046 800 0 FreeSans 224 90 0 0 io_oeb[33]
port 75 nsew signal tristate
flabel metal2 s 59082 0 59138 800 0 FreeSans 224 90 0 0 io_oeb[34]
port 76 nsew signal tristate
flabel metal2 s 59174 0 59230 800 0 FreeSans 224 90 0 0 io_oeb[35]
port 77 nsew signal tristate
flabel metal2 s 59266 0 59322 800 0 FreeSans 224 90 0 0 io_oeb[36]
port 78 nsew signal tristate
flabel metal2 s 59358 0 59414 800 0 FreeSans 224 90 0 0 io_oeb[37]
port 79 nsew signal tristate
flabel metal2 s 56230 0 56286 800 0 FreeSans 224 90 0 0 io_oeb[3]
port 80 nsew signal tristate
flabel metal2 s 56322 0 56378 800 0 FreeSans 224 90 0 0 io_oeb[4]
port 81 nsew signal tristate
flabel metal2 s 56414 0 56470 800 0 FreeSans 224 90 0 0 io_oeb[5]
port 82 nsew signal tristate
flabel metal2 s 56506 0 56562 800 0 FreeSans 224 90 0 0 io_oeb[6]
port 83 nsew signal tristate
flabel metal2 s 56598 0 56654 800 0 FreeSans 224 90 0 0 io_oeb[7]
port 84 nsew signal tristate
flabel metal2 s 56690 0 56746 800 0 FreeSans 224 90 0 0 io_oeb[8]
port 85 nsew signal tristate
flabel metal2 s 56782 0 56838 800 0 FreeSans 224 90 0 0 io_oeb[9]
port 86 nsew signal tristate
flabel metal3 s 69200 688 70000 808 0 FreeSans 480 0 0 0 io_out[0]
port 87 nsew signal tristate
flabel metal3 s 69200 14288 70000 14408 0 FreeSans 480 0 0 0 io_out[10]
port 88 nsew signal tristate
flabel metal3 s 69200 15648 70000 15768 0 FreeSans 480 0 0 0 io_out[11]
port 89 nsew signal tristate
flabel metal3 s 69200 17008 70000 17128 0 FreeSans 480 0 0 0 io_out[12]
port 90 nsew signal tristate
flabel metal3 s 69200 18368 70000 18488 0 FreeSans 480 0 0 0 io_out[13]
port 91 nsew signal tristate
flabel metal3 s 69200 19728 70000 19848 0 FreeSans 480 0 0 0 io_out[14]
port 92 nsew signal tristate
flabel metal3 s 69200 21088 70000 21208 0 FreeSans 480 0 0 0 io_out[15]
port 93 nsew signal tristate
flabel metal3 s 69200 22448 70000 22568 0 FreeSans 480 0 0 0 io_out[16]
port 94 nsew signal tristate
flabel metal3 s 69200 23808 70000 23928 0 FreeSans 480 0 0 0 io_out[17]
port 95 nsew signal tristate
flabel metal3 s 69200 25168 70000 25288 0 FreeSans 480 0 0 0 io_out[18]
port 96 nsew signal tristate
flabel metal3 s 69200 26528 70000 26648 0 FreeSans 480 0 0 0 io_out[19]
port 97 nsew signal tristate
flabel metal3 s 69200 2048 70000 2168 0 FreeSans 480 0 0 0 io_out[1]
port 98 nsew signal tristate
flabel metal3 s 69200 27888 70000 28008 0 FreeSans 480 0 0 0 io_out[20]
port 99 nsew signal tristate
flabel metal3 s 69200 29248 70000 29368 0 FreeSans 480 0 0 0 io_out[21]
port 100 nsew signal tristate
flabel metal3 s 69200 30608 70000 30728 0 FreeSans 480 0 0 0 io_out[22]
port 101 nsew signal tristate
flabel metal3 s 69200 31968 70000 32088 0 FreeSans 480 0 0 0 io_out[23]
port 102 nsew signal tristate
flabel metal3 s 69200 33328 70000 33448 0 FreeSans 480 0 0 0 io_out[24]
port 103 nsew signal tristate
flabel metal3 s 69200 34688 70000 34808 0 FreeSans 480 0 0 0 io_out[25]
port 104 nsew signal tristate
flabel metal3 s 69200 36048 70000 36168 0 FreeSans 480 0 0 0 io_out[26]
port 105 nsew signal tristate
flabel metal3 s 69200 37408 70000 37528 0 FreeSans 480 0 0 0 io_out[27]
port 106 nsew signal tristate
flabel metal3 s 69200 38768 70000 38888 0 FreeSans 480 0 0 0 io_out[28]
port 107 nsew signal tristate
flabel metal3 s 69200 40128 70000 40248 0 FreeSans 480 0 0 0 io_out[29]
port 108 nsew signal tristate
flabel metal3 s 69200 3408 70000 3528 0 FreeSans 480 0 0 0 io_out[2]
port 109 nsew signal tristate
flabel metal3 s 69200 41488 70000 41608 0 FreeSans 480 0 0 0 io_out[30]
port 110 nsew signal tristate
flabel metal3 s 69200 42848 70000 42968 0 FreeSans 480 0 0 0 io_out[31]
port 111 nsew signal tristate
flabel metal3 s 69200 44208 70000 44328 0 FreeSans 480 0 0 0 io_out[32]
port 112 nsew signal tristate
flabel metal3 s 69200 45568 70000 45688 0 FreeSans 480 0 0 0 io_out[33]
port 113 nsew signal tristate
flabel metal3 s 69200 46928 70000 47048 0 FreeSans 480 0 0 0 io_out[34]
port 114 nsew signal tristate
flabel metal3 s 69200 48288 70000 48408 0 FreeSans 480 0 0 0 io_out[35]
port 115 nsew signal tristate
flabel metal3 s 69200 49648 70000 49768 0 FreeSans 480 0 0 0 io_out[36]
port 116 nsew signal tristate
flabel metal3 s 69200 51008 70000 51128 0 FreeSans 480 0 0 0 io_out[37]
port 117 nsew signal tristate
flabel metal3 s 69200 4768 70000 4888 0 FreeSans 480 0 0 0 io_out[3]
port 118 nsew signal tristate
flabel metal3 s 69200 6128 70000 6248 0 FreeSans 480 0 0 0 io_out[4]
port 119 nsew signal tristate
flabel metal3 s 69200 7488 70000 7608 0 FreeSans 480 0 0 0 io_out[5]
port 120 nsew signal tristate
flabel metal3 s 69200 8848 70000 8968 0 FreeSans 480 0 0 0 io_out[6]
port 121 nsew signal tristate
flabel metal3 s 69200 10208 70000 10328 0 FreeSans 480 0 0 0 io_out[7]
port 122 nsew signal tristate
flabel metal3 s 69200 11568 70000 11688 0 FreeSans 480 0 0 0 io_out[8]
port 123 nsew signal tristate
flabel metal3 s 69200 12928 70000 13048 0 FreeSans 480 0 0 0 io_out[9]
port 124 nsew signal tristate
flabel metal2 s 55678 0 55734 800 0 FreeSans 224 90 0 0 irq[0]
port 125 nsew signal tristate
flabel metal2 s 55770 0 55826 800 0 FreeSans 224 90 0 0 irq[1]
port 126 nsew signal tristate
flabel metal2 s 55862 0 55918 800 0 FreeSans 224 90 0 0 irq[2]
port 127 nsew signal tristate
flabel metal2 s 20350 0 20406 800 0 FreeSans 224 90 0 0 la_data_in[0]
port 128 nsew signal input
flabel metal2 s 47950 0 48006 800 0 FreeSans 224 90 0 0 la_data_in[100]
port 129 nsew signal input
flabel metal2 s 48226 0 48282 800 0 FreeSans 224 90 0 0 la_data_in[101]
port 130 nsew signal input
flabel metal2 s 48502 0 48558 800 0 FreeSans 224 90 0 0 la_data_in[102]
port 131 nsew signal input
flabel metal2 s 48778 0 48834 800 0 FreeSans 224 90 0 0 la_data_in[103]
port 132 nsew signal input
flabel metal2 s 49054 0 49110 800 0 FreeSans 224 90 0 0 la_data_in[104]
port 133 nsew signal input
flabel metal2 s 49330 0 49386 800 0 FreeSans 224 90 0 0 la_data_in[105]
port 134 nsew signal input
flabel metal2 s 49606 0 49662 800 0 FreeSans 224 90 0 0 la_data_in[106]
port 135 nsew signal input
flabel metal2 s 49882 0 49938 800 0 FreeSans 224 90 0 0 la_data_in[107]
port 136 nsew signal input
flabel metal2 s 50158 0 50214 800 0 FreeSans 224 90 0 0 la_data_in[108]
port 137 nsew signal input
flabel metal2 s 50434 0 50490 800 0 FreeSans 224 90 0 0 la_data_in[109]
port 138 nsew signal input
flabel metal2 s 23110 0 23166 800 0 FreeSans 224 90 0 0 la_data_in[10]
port 139 nsew signal input
flabel metal2 s 50710 0 50766 800 0 FreeSans 224 90 0 0 la_data_in[110]
port 140 nsew signal input
flabel metal2 s 50986 0 51042 800 0 FreeSans 224 90 0 0 la_data_in[111]
port 141 nsew signal input
flabel metal2 s 51262 0 51318 800 0 FreeSans 224 90 0 0 la_data_in[112]
port 142 nsew signal input
flabel metal2 s 51538 0 51594 800 0 FreeSans 224 90 0 0 la_data_in[113]
port 143 nsew signal input
flabel metal2 s 51814 0 51870 800 0 FreeSans 224 90 0 0 la_data_in[114]
port 144 nsew signal input
flabel metal2 s 52090 0 52146 800 0 FreeSans 224 90 0 0 la_data_in[115]
port 145 nsew signal input
flabel metal2 s 52366 0 52422 800 0 FreeSans 224 90 0 0 la_data_in[116]
port 146 nsew signal input
flabel metal2 s 52642 0 52698 800 0 FreeSans 224 90 0 0 la_data_in[117]
port 147 nsew signal input
flabel metal2 s 52918 0 52974 800 0 FreeSans 224 90 0 0 la_data_in[118]
port 148 nsew signal input
flabel metal2 s 53194 0 53250 800 0 FreeSans 224 90 0 0 la_data_in[119]
port 149 nsew signal input
flabel metal2 s 23386 0 23442 800 0 FreeSans 224 90 0 0 la_data_in[11]
port 150 nsew signal input
flabel metal2 s 53470 0 53526 800 0 FreeSans 224 90 0 0 la_data_in[120]
port 151 nsew signal input
flabel metal2 s 53746 0 53802 800 0 FreeSans 224 90 0 0 la_data_in[121]
port 152 nsew signal input
flabel metal2 s 54022 0 54078 800 0 FreeSans 224 90 0 0 la_data_in[122]
port 153 nsew signal input
flabel metal2 s 54298 0 54354 800 0 FreeSans 224 90 0 0 la_data_in[123]
port 154 nsew signal input
flabel metal2 s 54574 0 54630 800 0 FreeSans 224 90 0 0 la_data_in[124]
port 155 nsew signal input
flabel metal2 s 54850 0 54906 800 0 FreeSans 224 90 0 0 la_data_in[125]
port 156 nsew signal input
flabel metal2 s 55126 0 55182 800 0 FreeSans 224 90 0 0 la_data_in[126]
port 157 nsew signal input
flabel metal2 s 55402 0 55458 800 0 FreeSans 224 90 0 0 la_data_in[127]
port 158 nsew signal input
flabel metal2 s 23662 0 23718 800 0 FreeSans 224 90 0 0 la_data_in[12]
port 159 nsew signal input
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 la_data_in[13]
port 160 nsew signal input
flabel metal2 s 24214 0 24270 800 0 FreeSans 224 90 0 0 la_data_in[14]
port 161 nsew signal input
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 la_data_in[15]
port 162 nsew signal input
flabel metal2 s 24766 0 24822 800 0 FreeSans 224 90 0 0 la_data_in[16]
port 163 nsew signal input
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 la_data_in[17]
port 164 nsew signal input
flabel metal2 s 25318 0 25374 800 0 FreeSans 224 90 0 0 la_data_in[18]
port 165 nsew signal input
flabel metal2 s 25594 0 25650 800 0 FreeSans 224 90 0 0 la_data_in[19]
port 166 nsew signal input
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 la_data_in[1]
port 167 nsew signal input
flabel metal2 s 25870 0 25926 800 0 FreeSans 224 90 0 0 la_data_in[20]
port 168 nsew signal input
flabel metal2 s 26146 0 26202 800 0 FreeSans 224 90 0 0 la_data_in[21]
port 169 nsew signal input
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 la_data_in[22]
port 170 nsew signal input
flabel metal2 s 26698 0 26754 800 0 FreeSans 224 90 0 0 la_data_in[23]
port 171 nsew signal input
flabel metal2 s 26974 0 27030 800 0 FreeSans 224 90 0 0 la_data_in[24]
port 172 nsew signal input
flabel metal2 s 27250 0 27306 800 0 FreeSans 224 90 0 0 la_data_in[25]
port 173 nsew signal input
flabel metal2 s 27526 0 27582 800 0 FreeSans 224 90 0 0 la_data_in[26]
port 174 nsew signal input
flabel metal2 s 27802 0 27858 800 0 FreeSans 224 90 0 0 la_data_in[27]
port 175 nsew signal input
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 la_data_in[28]
port 176 nsew signal input
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 la_data_in[29]
port 177 nsew signal input
flabel metal2 s 20902 0 20958 800 0 FreeSans 224 90 0 0 la_data_in[2]
port 178 nsew signal input
flabel metal2 s 28630 0 28686 800 0 FreeSans 224 90 0 0 la_data_in[30]
port 179 nsew signal input
flabel metal2 s 28906 0 28962 800 0 FreeSans 224 90 0 0 la_data_in[31]
port 180 nsew signal input
flabel metal2 s 29182 0 29238 800 0 FreeSans 224 90 0 0 la_data_in[32]
port 181 nsew signal input
flabel metal2 s 29458 0 29514 800 0 FreeSans 224 90 0 0 la_data_in[33]
port 182 nsew signal input
flabel metal2 s 29734 0 29790 800 0 FreeSans 224 90 0 0 la_data_in[34]
port 183 nsew signal input
flabel metal2 s 30010 0 30066 800 0 FreeSans 224 90 0 0 la_data_in[35]
port 184 nsew signal input
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 la_data_in[36]
port 185 nsew signal input
flabel metal2 s 30562 0 30618 800 0 FreeSans 224 90 0 0 la_data_in[37]
port 186 nsew signal input
flabel metal2 s 30838 0 30894 800 0 FreeSans 224 90 0 0 la_data_in[38]
port 187 nsew signal input
flabel metal2 s 31114 0 31170 800 0 FreeSans 224 90 0 0 la_data_in[39]
port 188 nsew signal input
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 la_data_in[3]
port 189 nsew signal input
flabel metal2 s 31390 0 31446 800 0 FreeSans 224 90 0 0 la_data_in[40]
port 190 nsew signal input
flabel metal2 s 31666 0 31722 800 0 FreeSans 224 90 0 0 la_data_in[41]
port 191 nsew signal input
flabel metal2 s 31942 0 31998 800 0 FreeSans 224 90 0 0 la_data_in[42]
port 192 nsew signal input
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 la_data_in[43]
port 193 nsew signal input
flabel metal2 s 32494 0 32550 800 0 FreeSans 224 90 0 0 la_data_in[44]
port 194 nsew signal input
flabel metal2 s 32770 0 32826 800 0 FreeSans 224 90 0 0 la_data_in[45]
port 195 nsew signal input
flabel metal2 s 33046 0 33102 800 0 FreeSans 224 90 0 0 la_data_in[46]
port 196 nsew signal input
flabel metal2 s 33322 0 33378 800 0 FreeSans 224 90 0 0 la_data_in[47]
port 197 nsew signal input
flabel metal2 s 33598 0 33654 800 0 FreeSans 224 90 0 0 la_data_in[48]
port 198 nsew signal input
flabel metal2 s 33874 0 33930 800 0 FreeSans 224 90 0 0 la_data_in[49]
port 199 nsew signal input
flabel metal2 s 21454 0 21510 800 0 FreeSans 224 90 0 0 la_data_in[4]
port 200 nsew signal input
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 la_data_in[50]
port 201 nsew signal input
flabel metal2 s 34426 0 34482 800 0 FreeSans 224 90 0 0 la_data_in[51]
port 202 nsew signal input
flabel metal2 s 34702 0 34758 800 0 FreeSans 224 90 0 0 la_data_in[52]
port 203 nsew signal input
flabel metal2 s 34978 0 35034 800 0 FreeSans 224 90 0 0 la_data_in[53]
port 204 nsew signal input
flabel metal2 s 35254 0 35310 800 0 FreeSans 224 90 0 0 la_data_in[54]
port 205 nsew signal input
flabel metal2 s 35530 0 35586 800 0 FreeSans 224 90 0 0 la_data_in[55]
port 206 nsew signal input
flabel metal2 s 35806 0 35862 800 0 FreeSans 224 90 0 0 la_data_in[56]
port 207 nsew signal input
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 la_data_in[57]
port 208 nsew signal input
flabel metal2 s 36358 0 36414 800 0 FreeSans 224 90 0 0 la_data_in[58]
port 209 nsew signal input
flabel metal2 s 36634 0 36690 800 0 FreeSans 224 90 0 0 la_data_in[59]
port 210 nsew signal input
flabel metal2 s 21730 0 21786 800 0 FreeSans 224 90 0 0 la_data_in[5]
port 211 nsew signal input
flabel metal2 s 36910 0 36966 800 0 FreeSans 224 90 0 0 la_data_in[60]
port 212 nsew signal input
flabel metal2 s 37186 0 37242 800 0 FreeSans 224 90 0 0 la_data_in[61]
port 213 nsew signal input
flabel metal2 s 37462 0 37518 800 0 FreeSans 224 90 0 0 la_data_in[62]
port 214 nsew signal input
flabel metal2 s 37738 0 37794 800 0 FreeSans 224 90 0 0 la_data_in[63]
port 215 nsew signal input
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 la_data_in[64]
port 216 nsew signal input
flabel metal2 s 38290 0 38346 800 0 FreeSans 224 90 0 0 la_data_in[65]
port 217 nsew signal input
flabel metal2 s 38566 0 38622 800 0 FreeSans 224 90 0 0 la_data_in[66]
port 218 nsew signal input
flabel metal2 s 38842 0 38898 800 0 FreeSans 224 90 0 0 la_data_in[67]
port 219 nsew signal input
flabel metal2 s 39118 0 39174 800 0 FreeSans 224 90 0 0 la_data_in[68]
port 220 nsew signal input
flabel metal2 s 39394 0 39450 800 0 FreeSans 224 90 0 0 la_data_in[69]
port 221 nsew signal input
flabel metal2 s 22006 0 22062 800 0 FreeSans 224 90 0 0 la_data_in[6]
port 222 nsew signal input
flabel metal2 s 39670 0 39726 800 0 FreeSans 224 90 0 0 la_data_in[70]
port 223 nsew signal input
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 la_data_in[71]
port 224 nsew signal input
flabel metal2 s 40222 0 40278 800 0 FreeSans 224 90 0 0 la_data_in[72]
port 225 nsew signal input
flabel metal2 s 40498 0 40554 800 0 FreeSans 224 90 0 0 la_data_in[73]
port 226 nsew signal input
flabel metal2 s 40774 0 40830 800 0 FreeSans 224 90 0 0 la_data_in[74]
port 227 nsew signal input
flabel metal2 s 41050 0 41106 800 0 FreeSans 224 90 0 0 la_data_in[75]
port 228 nsew signal input
flabel metal2 s 41326 0 41382 800 0 FreeSans 224 90 0 0 la_data_in[76]
port 229 nsew signal input
flabel metal2 s 41602 0 41658 800 0 FreeSans 224 90 0 0 la_data_in[77]
port 230 nsew signal input
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 la_data_in[78]
port 231 nsew signal input
flabel metal2 s 42154 0 42210 800 0 FreeSans 224 90 0 0 la_data_in[79]
port 232 nsew signal input
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 la_data_in[7]
port 233 nsew signal input
flabel metal2 s 42430 0 42486 800 0 FreeSans 224 90 0 0 la_data_in[80]
port 234 nsew signal input
flabel metal2 s 42706 0 42762 800 0 FreeSans 224 90 0 0 la_data_in[81]
port 235 nsew signal input
flabel metal2 s 42982 0 43038 800 0 FreeSans 224 90 0 0 la_data_in[82]
port 236 nsew signal input
flabel metal2 s 43258 0 43314 800 0 FreeSans 224 90 0 0 la_data_in[83]
port 237 nsew signal input
flabel metal2 s 43534 0 43590 800 0 FreeSans 224 90 0 0 la_data_in[84]
port 238 nsew signal input
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 la_data_in[85]
port 239 nsew signal input
flabel metal2 s 44086 0 44142 800 0 FreeSans 224 90 0 0 la_data_in[86]
port 240 nsew signal input
flabel metal2 s 44362 0 44418 800 0 FreeSans 224 90 0 0 la_data_in[87]
port 241 nsew signal input
flabel metal2 s 44638 0 44694 800 0 FreeSans 224 90 0 0 la_data_in[88]
port 242 nsew signal input
flabel metal2 s 44914 0 44970 800 0 FreeSans 224 90 0 0 la_data_in[89]
port 243 nsew signal input
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 la_data_in[8]
port 244 nsew signal input
flabel metal2 s 45190 0 45246 800 0 FreeSans 224 90 0 0 la_data_in[90]
port 245 nsew signal input
flabel metal2 s 45466 0 45522 800 0 FreeSans 224 90 0 0 la_data_in[91]
port 246 nsew signal input
flabel metal2 s 45742 0 45798 800 0 FreeSans 224 90 0 0 la_data_in[92]
port 247 nsew signal input
flabel metal2 s 46018 0 46074 800 0 FreeSans 224 90 0 0 la_data_in[93]
port 248 nsew signal input
flabel metal2 s 46294 0 46350 800 0 FreeSans 224 90 0 0 la_data_in[94]
port 249 nsew signal input
flabel metal2 s 46570 0 46626 800 0 FreeSans 224 90 0 0 la_data_in[95]
port 250 nsew signal input
flabel metal2 s 46846 0 46902 800 0 FreeSans 224 90 0 0 la_data_in[96]
port 251 nsew signal input
flabel metal2 s 47122 0 47178 800 0 FreeSans 224 90 0 0 la_data_in[97]
port 252 nsew signal input
flabel metal2 s 47398 0 47454 800 0 FreeSans 224 90 0 0 la_data_in[98]
port 253 nsew signal input
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 la_data_in[99]
port 254 nsew signal input
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 la_data_in[9]
port 255 nsew signal input
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 la_data_out[0]
port 256 nsew signal tristate
flabel metal2 s 48042 0 48098 800 0 FreeSans 224 90 0 0 la_data_out[100]
port 257 nsew signal tristate
flabel metal2 s 48318 0 48374 800 0 FreeSans 224 90 0 0 la_data_out[101]
port 258 nsew signal tristate
flabel metal2 s 48594 0 48650 800 0 FreeSans 224 90 0 0 la_data_out[102]
port 259 nsew signal tristate
flabel metal2 s 48870 0 48926 800 0 FreeSans 224 90 0 0 la_data_out[103]
port 260 nsew signal tristate
flabel metal2 s 49146 0 49202 800 0 FreeSans 224 90 0 0 la_data_out[104]
port 261 nsew signal tristate
flabel metal2 s 49422 0 49478 800 0 FreeSans 224 90 0 0 la_data_out[105]
port 262 nsew signal tristate
flabel metal2 s 49698 0 49754 800 0 FreeSans 224 90 0 0 la_data_out[106]
port 263 nsew signal tristate
flabel metal2 s 49974 0 50030 800 0 FreeSans 224 90 0 0 la_data_out[107]
port 264 nsew signal tristate
flabel metal2 s 50250 0 50306 800 0 FreeSans 224 90 0 0 la_data_out[108]
port 265 nsew signal tristate
flabel metal2 s 50526 0 50582 800 0 FreeSans 224 90 0 0 la_data_out[109]
port 266 nsew signal tristate
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 la_data_out[10]
port 267 nsew signal tristate
flabel metal2 s 50802 0 50858 800 0 FreeSans 224 90 0 0 la_data_out[110]
port 268 nsew signal tristate
flabel metal2 s 51078 0 51134 800 0 FreeSans 224 90 0 0 la_data_out[111]
port 269 nsew signal tristate
flabel metal2 s 51354 0 51410 800 0 FreeSans 224 90 0 0 la_data_out[112]
port 270 nsew signal tristate
flabel metal2 s 51630 0 51686 800 0 FreeSans 224 90 0 0 la_data_out[113]
port 271 nsew signal tristate
flabel metal2 s 51906 0 51962 800 0 FreeSans 224 90 0 0 la_data_out[114]
port 272 nsew signal tristate
flabel metal2 s 52182 0 52238 800 0 FreeSans 224 90 0 0 la_data_out[115]
port 273 nsew signal tristate
flabel metal2 s 52458 0 52514 800 0 FreeSans 224 90 0 0 la_data_out[116]
port 274 nsew signal tristate
flabel metal2 s 52734 0 52790 800 0 FreeSans 224 90 0 0 la_data_out[117]
port 275 nsew signal tristate
flabel metal2 s 53010 0 53066 800 0 FreeSans 224 90 0 0 la_data_out[118]
port 276 nsew signal tristate
flabel metal2 s 53286 0 53342 800 0 FreeSans 224 90 0 0 la_data_out[119]
port 277 nsew signal tristate
flabel metal2 s 23478 0 23534 800 0 FreeSans 224 90 0 0 la_data_out[11]
port 278 nsew signal tristate
flabel metal2 s 53562 0 53618 800 0 FreeSans 224 90 0 0 la_data_out[120]
port 279 nsew signal tristate
flabel metal2 s 53838 0 53894 800 0 FreeSans 224 90 0 0 la_data_out[121]
port 280 nsew signal tristate
flabel metal2 s 54114 0 54170 800 0 FreeSans 224 90 0 0 la_data_out[122]
port 281 nsew signal tristate
flabel metal2 s 54390 0 54446 800 0 FreeSans 224 90 0 0 la_data_out[123]
port 282 nsew signal tristate
flabel metal2 s 54666 0 54722 800 0 FreeSans 224 90 0 0 la_data_out[124]
port 283 nsew signal tristate
flabel metal2 s 54942 0 54998 800 0 FreeSans 224 90 0 0 la_data_out[125]
port 284 nsew signal tristate
flabel metal2 s 55218 0 55274 800 0 FreeSans 224 90 0 0 la_data_out[126]
port 285 nsew signal tristate
flabel metal2 s 55494 0 55550 800 0 FreeSans 224 90 0 0 la_data_out[127]
port 286 nsew signal tristate
flabel metal2 s 23754 0 23810 800 0 FreeSans 224 90 0 0 la_data_out[12]
port 287 nsew signal tristate
flabel metal2 s 24030 0 24086 800 0 FreeSans 224 90 0 0 la_data_out[13]
port 288 nsew signal tristate
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 la_data_out[14]
port 289 nsew signal tristate
flabel metal2 s 24582 0 24638 800 0 FreeSans 224 90 0 0 la_data_out[15]
port 290 nsew signal tristate
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 la_data_out[16]
port 291 nsew signal tristate
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 la_data_out[17]
port 292 nsew signal tristate
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 la_data_out[18]
port 293 nsew signal tristate
flabel metal2 s 25686 0 25742 800 0 FreeSans 224 90 0 0 la_data_out[19]
port 294 nsew signal tristate
flabel metal2 s 20718 0 20774 800 0 FreeSans 224 90 0 0 la_data_out[1]
port 295 nsew signal tristate
flabel metal2 s 25962 0 26018 800 0 FreeSans 224 90 0 0 la_data_out[20]
port 296 nsew signal tristate
flabel metal2 s 26238 0 26294 800 0 FreeSans 224 90 0 0 la_data_out[21]
port 297 nsew signal tristate
flabel metal2 s 26514 0 26570 800 0 FreeSans 224 90 0 0 la_data_out[22]
port 298 nsew signal tristate
flabel metal2 s 26790 0 26846 800 0 FreeSans 224 90 0 0 la_data_out[23]
port 299 nsew signal tristate
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 la_data_out[24]
port 300 nsew signal tristate
flabel metal2 s 27342 0 27398 800 0 FreeSans 224 90 0 0 la_data_out[25]
port 301 nsew signal tristate
flabel metal2 s 27618 0 27674 800 0 FreeSans 224 90 0 0 la_data_out[26]
port 302 nsew signal tristate
flabel metal2 s 27894 0 27950 800 0 FreeSans 224 90 0 0 la_data_out[27]
port 303 nsew signal tristate
flabel metal2 s 28170 0 28226 800 0 FreeSans 224 90 0 0 la_data_out[28]
port 304 nsew signal tristate
flabel metal2 s 28446 0 28502 800 0 FreeSans 224 90 0 0 la_data_out[29]
port 305 nsew signal tristate
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 la_data_out[2]
port 306 nsew signal tristate
flabel metal2 s 28722 0 28778 800 0 FreeSans 224 90 0 0 la_data_out[30]
port 307 nsew signal tristate
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 la_data_out[31]
port 308 nsew signal tristate
flabel metal2 s 29274 0 29330 800 0 FreeSans 224 90 0 0 la_data_out[32]
port 309 nsew signal tristate
flabel metal2 s 29550 0 29606 800 0 FreeSans 224 90 0 0 la_data_out[33]
port 310 nsew signal tristate
flabel metal2 s 29826 0 29882 800 0 FreeSans 224 90 0 0 la_data_out[34]
port 311 nsew signal tristate
flabel metal2 s 30102 0 30158 800 0 FreeSans 224 90 0 0 la_data_out[35]
port 312 nsew signal tristate
flabel metal2 s 30378 0 30434 800 0 FreeSans 224 90 0 0 la_data_out[36]
port 313 nsew signal tristate
flabel metal2 s 30654 0 30710 800 0 FreeSans 224 90 0 0 la_data_out[37]
port 314 nsew signal tristate
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 la_data_out[38]
port 315 nsew signal tristate
flabel metal2 s 31206 0 31262 800 0 FreeSans 224 90 0 0 la_data_out[39]
port 316 nsew signal tristate
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 la_data_out[3]
port 317 nsew signal tristate
flabel metal2 s 31482 0 31538 800 0 FreeSans 224 90 0 0 la_data_out[40]
port 318 nsew signal tristate
flabel metal2 s 31758 0 31814 800 0 FreeSans 224 90 0 0 la_data_out[41]
port 319 nsew signal tristate
flabel metal2 s 32034 0 32090 800 0 FreeSans 224 90 0 0 la_data_out[42]
port 320 nsew signal tristate
flabel metal2 s 32310 0 32366 800 0 FreeSans 224 90 0 0 la_data_out[43]
port 321 nsew signal tristate
flabel metal2 s 32586 0 32642 800 0 FreeSans 224 90 0 0 la_data_out[44]
port 322 nsew signal tristate
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 la_data_out[45]
port 323 nsew signal tristate
flabel metal2 s 33138 0 33194 800 0 FreeSans 224 90 0 0 la_data_out[46]
port 324 nsew signal tristate
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 la_data_out[47]
port 325 nsew signal tristate
flabel metal2 s 33690 0 33746 800 0 FreeSans 224 90 0 0 la_data_out[48]
port 326 nsew signal tristate
flabel metal2 s 33966 0 34022 800 0 FreeSans 224 90 0 0 la_data_out[49]
port 327 nsew signal tristate
flabel metal2 s 21546 0 21602 800 0 FreeSans 224 90 0 0 la_data_out[4]
port 328 nsew signal tristate
flabel metal2 s 34242 0 34298 800 0 FreeSans 224 90 0 0 la_data_out[50]
port 329 nsew signal tristate
flabel metal2 s 34518 0 34574 800 0 FreeSans 224 90 0 0 la_data_out[51]
port 330 nsew signal tristate
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 la_data_out[52]
port 331 nsew signal tristate
flabel metal2 s 35070 0 35126 800 0 FreeSans 224 90 0 0 la_data_out[53]
port 332 nsew signal tristate
flabel metal2 s 35346 0 35402 800 0 FreeSans 224 90 0 0 la_data_out[54]
port 333 nsew signal tristate
flabel metal2 s 35622 0 35678 800 0 FreeSans 224 90 0 0 la_data_out[55]
port 334 nsew signal tristate
flabel metal2 s 35898 0 35954 800 0 FreeSans 224 90 0 0 la_data_out[56]
port 335 nsew signal tristate
flabel metal2 s 36174 0 36230 800 0 FreeSans 224 90 0 0 la_data_out[57]
port 336 nsew signal tristate
flabel metal2 s 36450 0 36506 800 0 FreeSans 224 90 0 0 la_data_out[58]
port 337 nsew signal tristate
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 la_data_out[59]
port 338 nsew signal tristate
flabel metal2 s 21822 0 21878 800 0 FreeSans 224 90 0 0 la_data_out[5]
port 339 nsew signal tristate
flabel metal2 s 37002 0 37058 800 0 FreeSans 224 90 0 0 la_data_out[60]
port 340 nsew signal tristate
flabel metal2 s 37278 0 37334 800 0 FreeSans 224 90 0 0 la_data_out[61]
port 341 nsew signal tristate
flabel metal2 s 37554 0 37610 800 0 FreeSans 224 90 0 0 la_data_out[62]
port 342 nsew signal tristate
flabel metal2 s 37830 0 37886 800 0 FreeSans 224 90 0 0 la_data_out[63]
port 343 nsew signal tristate
flabel metal2 s 38106 0 38162 800 0 FreeSans 224 90 0 0 la_data_out[64]
port 344 nsew signal tristate
flabel metal2 s 38382 0 38438 800 0 FreeSans 224 90 0 0 la_data_out[65]
port 345 nsew signal tristate
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 la_data_out[66]
port 346 nsew signal tristate
flabel metal2 s 38934 0 38990 800 0 FreeSans 224 90 0 0 la_data_out[67]
port 347 nsew signal tristate
flabel metal2 s 39210 0 39266 800 0 FreeSans 224 90 0 0 la_data_out[68]
port 348 nsew signal tristate
flabel metal2 s 39486 0 39542 800 0 FreeSans 224 90 0 0 la_data_out[69]
port 349 nsew signal tristate
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 la_data_out[6]
port 350 nsew signal tristate
flabel metal2 s 39762 0 39818 800 0 FreeSans 224 90 0 0 la_data_out[70]
port 351 nsew signal tristate
flabel metal2 s 40038 0 40094 800 0 FreeSans 224 90 0 0 la_data_out[71]
port 352 nsew signal tristate
flabel metal2 s 40314 0 40370 800 0 FreeSans 224 90 0 0 la_data_out[72]
port 353 nsew signal tristate
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 la_data_out[73]
port 354 nsew signal tristate
flabel metal2 s 40866 0 40922 800 0 FreeSans 224 90 0 0 la_data_out[74]
port 355 nsew signal tristate
flabel metal2 s 41142 0 41198 800 0 FreeSans 224 90 0 0 la_data_out[75]
port 356 nsew signal tristate
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 la_data_out[76]
port 357 nsew signal tristate
flabel metal2 s 41694 0 41750 800 0 FreeSans 224 90 0 0 la_data_out[77]
port 358 nsew signal tristate
flabel metal2 s 41970 0 42026 800 0 FreeSans 224 90 0 0 la_data_out[78]
port 359 nsew signal tristate
flabel metal2 s 42246 0 42302 800 0 FreeSans 224 90 0 0 la_data_out[79]
port 360 nsew signal tristate
flabel metal2 s 22374 0 22430 800 0 FreeSans 224 90 0 0 la_data_out[7]
port 361 nsew signal tristate
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 la_data_out[80]
port 362 nsew signal tristate
flabel metal2 s 42798 0 42854 800 0 FreeSans 224 90 0 0 la_data_out[81]
port 363 nsew signal tristate
flabel metal2 s 43074 0 43130 800 0 FreeSans 224 90 0 0 la_data_out[82]
port 364 nsew signal tristate
flabel metal2 s 43350 0 43406 800 0 FreeSans 224 90 0 0 la_data_out[83]
port 365 nsew signal tristate
flabel metal2 s 43626 0 43682 800 0 FreeSans 224 90 0 0 la_data_out[84]
port 366 nsew signal tristate
flabel metal2 s 43902 0 43958 800 0 FreeSans 224 90 0 0 la_data_out[85]
port 367 nsew signal tristate
flabel metal2 s 44178 0 44234 800 0 FreeSans 224 90 0 0 la_data_out[86]
port 368 nsew signal tristate
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 la_data_out[87]
port 369 nsew signal tristate
flabel metal2 s 44730 0 44786 800 0 FreeSans 224 90 0 0 la_data_out[88]
port 370 nsew signal tristate
flabel metal2 s 45006 0 45062 800 0 FreeSans 224 90 0 0 la_data_out[89]
port 371 nsew signal tristate
flabel metal2 s 22650 0 22706 800 0 FreeSans 224 90 0 0 la_data_out[8]
port 372 nsew signal tristate
flabel metal2 s 45282 0 45338 800 0 FreeSans 224 90 0 0 la_data_out[90]
port 373 nsew signal tristate
flabel metal2 s 45558 0 45614 800 0 FreeSans 224 90 0 0 la_data_out[91]
port 374 nsew signal tristate
flabel metal2 s 45834 0 45890 800 0 FreeSans 224 90 0 0 la_data_out[92]
port 375 nsew signal tristate
flabel metal2 s 46110 0 46166 800 0 FreeSans 224 90 0 0 la_data_out[93]
port 376 nsew signal tristate
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 la_data_out[94]
port 377 nsew signal tristate
flabel metal2 s 46662 0 46718 800 0 FreeSans 224 90 0 0 la_data_out[95]
port 378 nsew signal tristate
flabel metal2 s 46938 0 46994 800 0 FreeSans 224 90 0 0 la_data_out[96]
port 379 nsew signal tristate
flabel metal2 s 47214 0 47270 800 0 FreeSans 224 90 0 0 la_data_out[97]
port 380 nsew signal tristate
flabel metal2 s 47490 0 47546 800 0 FreeSans 224 90 0 0 la_data_out[98]
port 381 nsew signal tristate
flabel metal2 s 47766 0 47822 800 0 FreeSans 224 90 0 0 la_data_out[99]
port 382 nsew signal tristate
flabel metal2 s 22926 0 22982 800 0 FreeSans 224 90 0 0 la_data_out[9]
port 383 nsew signal tristate
flabel metal2 s 20534 0 20590 800 0 FreeSans 224 90 0 0 la_oenb[0]
port 384 nsew signal input
flabel metal2 s 48134 0 48190 800 0 FreeSans 224 90 0 0 la_oenb[100]
port 385 nsew signal input
flabel metal2 s 48410 0 48466 800 0 FreeSans 224 90 0 0 la_oenb[101]
port 386 nsew signal input
flabel metal2 s 48686 0 48742 800 0 FreeSans 224 90 0 0 la_oenb[102]
port 387 nsew signal input
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 la_oenb[103]
port 388 nsew signal input
flabel metal2 s 49238 0 49294 800 0 FreeSans 224 90 0 0 la_oenb[104]
port 389 nsew signal input
flabel metal2 s 49514 0 49570 800 0 FreeSans 224 90 0 0 la_oenb[105]
port 390 nsew signal input
flabel metal2 s 49790 0 49846 800 0 FreeSans 224 90 0 0 la_oenb[106]
port 391 nsew signal input
flabel metal2 s 50066 0 50122 800 0 FreeSans 224 90 0 0 la_oenb[107]
port 392 nsew signal input
flabel metal2 s 50342 0 50398 800 0 FreeSans 224 90 0 0 la_oenb[108]
port 393 nsew signal input
flabel metal2 s 50618 0 50674 800 0 FreeSans 224 90 0 0 la_oenb[109]
port 394 nsew signal input
flabel metal2 s 23294 0 23350 800 0 FreeSans 224 90 0 0 la_oenb[10]
port 395 nsew signal input
flabel metal2 s 50894 0 50950 800 0 FreeSans 224 90 0 0 la_oenb[110]
port 396 nsew signal input
flabel metal2 s 51170 0 51226 800 0 FreeSans 224 90 0 0 la_oenb[111]
port 397 nsew signal input
flabel metal2 s 51446 0 51502 800 0 FreeSans 224 90 0 0 la_oenb[112]
port 398 nsew signal input
flabel metal2 s 51722 0 51778 800 0 FreeSans 224 90 0 0 la_oenb[113]
port 399 nsew signal input
flabel metal2 s 51998 0 52054 800 0 FreeSans 224 90 0 0 la_oenb[114]
port 400 nsew signal input
flabel metal2 s 52274 0 52330 800 0 FreeSans 224 90 0 0 la_oenb[115]
port 401 nsew signal input
flabel metal2 s 52550 0 52606 800 0 FreeSans 224 90 0 0 la_oenb[116]
port 402 nsew signal input
flabel metal2 s 52826 0 52882 800 0 FreeSans 224 90 0 0 la_oenb[117]
port 403 nsew signal input
flabel metal2 s 53102 0 53158 800 0 FreeSans 224 90 0 0 la_oenb[118]
port 404 nsew signal input
flabel metal2 s 53378 0 53434 800 0 FreeSans 224 90 0 0 la_oenb[119]
port 405 nsew signal input
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 la_oenb[11]
port 406 nsew signal input
flabel metal2 s 53654 0 53710 800 0 FreeSans 224 90 0 0 la_oenb[120]
port 407 nsew signal input
flabel metal2 s 53930 0 53986 800 0 FreeSans 224 90 0 0 la_oenb[121]
port 408 nsew signal input
flabel metal2 s 54206 0 54262 800 0 FreeSans 224 90 0 0 la_oenb[122]
port 409 nsew signal input
flabel metal2 s 54482 0 54538 800 0 FreeSans 224 90 0 0 la_oenb[123]
port 410 nsew signal input
flabel metal2 s 54758 0 54814 800 0 FreeSans 224 90 0 0 la_oenb[124]
port 411 nsew signal input
flabel metal2 s 55034 0 55090 800 0 FreeSans 224 90 0 0 la_oenb[125]
port 412 nsew signal input
flabel metal2 s 55310 0 55366 800 0 FreeSans 224 90 0 0 la_oenb[126]
port 413 nsew signal input
flabel metal2 s 55586 0 55642 800 0 FreeSans 224 90 0 0 la_oenb[127]
port 414 nsew signal input
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 la_oenb[12]
port 415 nsew signal input
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 la_oenb[13]
port 416 nsew signal input
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 la_oenb[14]
port 417 nsew signal input
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 la_oenb[15]
port 418 nsew signal input
flabel metal2 s 24950 0 25006 800 0 FreeSans 224 90 0 0 la_oenb[16]
port 419 nsew signal input
flabel metal2 s 25226 0 25282 800 0 FreeSans 224 90 0 0 la_oenb[17]
port 420 nsew signal input
flabel metal2 s 25502 0 25558 800 0 FreeSans 224 90 0 0 la_oenb[18]
port 421 nsew signal input
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 la_oenb[19]
port 422 nsew signal input
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 la_oenb[1]
port 423 nsew signal input
flabel metal2 s 26054 0 26110 800 0 FreeSans 224 90 0 0 la_oenb[20]
port 424 nsew signal input
flabel metal2 s 26330 0 26386 800 0 FreeSans 224 90 0 0 la_oenb[21]
port 425 nsew signal input
flabel metal2 s 26606 0 26662 800 0 FreeSans 224 90 0 0 la_oenb[22]
port 426 nsew signal input
flabel metal2 s 26882 0 26938 800 0 FreeSans 224 90 0 0 la_oenb[23]
port 427 nsew signal input
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 la_oenb[24]
port 428 nsew signal input
flabel metal2 s 27434 0 27490 800 0 FreeSans 224 90 0 0 la_oenb[25]
port 429 nsew signal input
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 la_oenb[26]
port 430 nsew signal input
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 la_oenb[27]
port 431 nsew signal input
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 la_oenb[28]
port 432 nsew signal input
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 la_oenb[29]
port 433 nsew signal input
flabel metal2 s 21086 0 21142 800 0 FreeSans 224 90 0 0 la_oenb[2]
port 434 nsew signal input
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 la_oenb[30]
port 435 nsew signal input
flabel metal2 s 29090 0 29146 800 0 FreeSans 224 90 0 0 la_oenb[31]
port 436 nsew signal input
flabel metal2 s 29366 0 29422 800 0 FreeSans 224 90 0 0 la_oenb[32]
port 437 nsew signal input
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 la_oenb[33]
port 438 nsew signal input
flabel metal2 s 29918 0 29974 800 0 FreeSans 224 90 0 0 la_oenb[34]
port 439 nsew signal input
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 la_oenb[35]
port 440 nsew signal input
flabel metal2 s 30470 0 30526 800 0 FreeSans 224 90 0 0 la_oenb[36]
port 441 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 la_oenb[37]
port 442 nsew signal input
flabel metal2 s 31022 0 31078 800 0 FreeSans 224 90 0 0 la_oenb[38]
port 443 nsew signal input
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 la_oenb[39]
port 444 nsew signal input
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 la_oenb[3]
port 445 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 la_oenb[40]
port 446 nsew signal input
flabel metal2 s 31850 0 31906 800 0 FreeSans 224 90 0 0 la_oenb[41]
port 447 nsew signal input
flabel metal2 s 32126 0 32182 800 0 FreeSans 224 90 0 0 la_oenb[42]
port 448 nsew signal input
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 la_oenb[43]
port 449 nsew signal input
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 la_oenb[44]
port 450 nsew signal input
flabel metal2 s 32954 0 33010 800 0 FreeSans 224 90 0 0 la_oenb[45]
port 451 nsew signal input
flabel metal2 s 33230 0 33286 800 0 FreeSans 224 90 0 0 la_oenb[46]
port 452 nsew signal input
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 la_oenb[47]
port 453 nsew signal input
flabel metal2 s 33782 0 33838 800 0 FreeSans 224 90 0 0 la_oenb[48]
port 454 nsew signal input
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 la_oenb[49]
port 455 nsew signal input
flabel metal2 s 21638 0 21694 800 0 FreeSans 224 90 0 0 la_oenb[4]
port 456 nsew signal input
flabel metal2 s 34334 0 34390 800 0 FreeSans 224 90 0 0 la_oenb[50]
port 457 nsew signal input
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 la_oenb[51]
port 458 nsew signal input
flabel metal2 s 34886 0 34942 800 0 FreeSans 224 90 0 0 la_oenb[52]
port 459 nsew signal input
flabel metal2 s 35162 0 35218 800 0 FreeSans 224 90 0 0 la_oenb[53]
port 460 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 la_oenb[54]
port 461 nsew signal input
flabel metal2 s 35714 0 35770 800 0 FreeSans 224 90 0 0 la_oenb[55]
port 462 nsew signal input
flabel metal2 s 35990 0 36046 800 0 FreeSans 224 90 0 0 la_oenb[56]
port 463 nsew signal input
flabel metal2 s 36266 0 36322 800 0 FreeSans 224 90 0 0 la_oenb[57]
port 464 nsew signal input
flabel metal2 s 36542 0 36598 800 0 FreeSans 224 90 0 0 la_oenb[58]
port 465 nsew signal input
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 la_oenb[59]
port 466 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 la_oenb[5]
port 467 nsew signal input
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 la_oenb[60]
port 468 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 la_oenb[61]
port 469 nsew signal input
flabel metal2 s 37646 0 37702 800 0 FreeSans 224 90 0 0 la_oenb[62]
port 470 nsew signal input
flabel metal2 s 37922 0 37978 800 0 FreeSans 224 90 0 0 la_oenb[63]
port 471 nsew signal input
flabel metal2 s 38198 0 38254 800 0 FreeSans 224 90 0 0 la_oenb[64]
port 472 nsew signal input
flabel metal2 s 38474 0 38530 800 0 FreeSans 224 90 0 0 la_oenb[65]
port 473 nsew signal input
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 la_oenb[66]
port 474 nsew signal input
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 la_oenb[67]
port 475 nsew signal input
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 la_oenb[68]
port 476 nsew signal input
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 la_oenb[69]
port 477 nsew signal input
flabel metal2 s 22190 0 22246 800 0 FreeSans 224 90 0 0 la_oenb[6]
port 478 nsew signal input
flabel metal2 s 39854 0 39910 800 0 FreeSans 224 90 0 0 la_oenb[70]
port 479 nsew signal input
flabel metal2 s 40130 0 40186 800 0 FreeSans 224 90 0 0 la_oenb[71]
port 480 nsew signal input
flabel metal2 s 40406 0 40462 800 0 FreeSans 224 90 0 0 la_oenb[72]
port 481 nsew signal input
flabel metal2 s 40682 0 40738 800 0 FreeSans 224 90 0 0 la_oenb[73]
port 482 nsew signal input
flabel metal2 s 40958 0 41014 800 0 FreeSans 224 90 0 0 la_oenb[74]
port 483 nsew signal input
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 la_oenb[75]
port 484 nsew signal input
flabel metal2 s 41510 0 41566 800 0 FreeSans 224 90 0 0 la_oenb[76]
port 485 nsew signal input
flabel metal2 s 41786 0 41842 800 0 FreeSans 224 90 0 0 la_oenb[77]
port 486 nsew signal input
flabel metal2 s 42062 0 42118 800 0 FreeSans 224 90 0 0 la_oenb[78]
port 487 nsew signal input
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 la_oenb[79]
port 488 nsew signal input
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 la_oenb[7]
port 489 nsew signal input
flabel metal2 s 42614 0 42670 800 0 FreeSans 224 90 0 0 la_oenb[80]
port 490 nsew signal input
flabel metal2 s 42890 0 42946 800 0 FreeSans 224 90 0 0 la_oenb[81]
port 491 nsew signal input
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 la_oenb[82]
port 492 nsew signal input
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 la_oenb[83]
port 493 nsew signal input
flabel metal2 s 43718 0 43774 800 0 FreeSans 224 90 0 0 la_oenb[84]
port 494 nsew signal input
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 la_oenb[85]
port 495 nsew signal input
flabel metal2 s 44270 0 44326 800 0 FreeSans 224 90 0 0 la_oenb[86]
port 496 nsew signal input
flabel metal2 s 44546 0 44602 800 0 FreeSans 224 90 0 0 la_oenb[87]
port 497 nsew signal input
flabel metal2 s 44822 0 44878 800 0 FreeSans 224 90 0 0 la_oenb[88]
port 498 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 la_oenb[89]
port 499 nsew signal input
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 la_oenb[8]
port 500 nsew signal input
flabel metal2 s 45374 0 45430 800 0 FreeSans 224 90 0 0 la_oenb[90]
port 501 nsew signal input
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 la_oenb[91]
port 502 nsew signal input
flabel metal2 s 45926 0 45982 800 0 FreeSans 224 90 0 0 la_oenb[92]
port 503 nsew signal input
flabel metal2 s 46202 0 46258 800 0 FreeSans 224 90 0 0 la_oenb[93]
port 504 nsew signal input
flabel metal2 s 46478 0 46534 800 0 FreeSans 224 90 0 0 la_oenb[94]
port 505 nsew signal input
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 la_oenb[95]
port 506 nsew signal input
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 la_oenb[96]
port 507 nsew signal input
flabel metal2 s 47306 0 47362 800 0 FreeSans 224 90 0 0 la_oenb[97]
port 508 nsew signal input
flabel metal2 s 47582 0 47638 800 0 FreeSans 224 90 0 0 la_oenb[98]
port 509 nsew signal input
flabel metal2 s 47858 0 47914 800 0 FreeSans 224 90 0 0 la_oenb[99]
port 510 nsew signal input
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 la_oenb[9]
port 511 nsew signal input
flabel metal3 s 69200 53728 70000 53848 0 FreeSans 480 0 0 0 rst_o
port 512 nsew signal tristate
flabel metal3 s 69200 56448 70000 56568 0 FreeSans 480 0 0 0 start_o
port 513 nsew signal tristate
flabel metal4 s 4208 2128 4528 57712 0 FreeSans 1920 90 0 0 vccd1
port 514 nsew power bidirectional
flabel metal4 s 34928 2128 35248 57712 0 FreeSans 1920 90 0 0 vccd1
port 514 nsew power bidirectional
flabel metal4 s 65648 2128 65968 57712 0 FreeSans 1920 90 0 0 vccd1
port 514 nsew power bidirectional
flabel metal4 s 19568 2128 19888 57712 0 FreeSans 1920 90 0 0 vssd1
port 515 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 57712 0 FreeSans 1920 90 0 0 vssd1
port 515 nsew ground bidirectional
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 wb_clk_i
port 516 nsew signal input
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 wb_rst_i
port 517 nsew signal input
flabel metal2 s 10782 0 10838 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 518 nsew signal tristate
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 519 nsew signal input
flabel metal2 s 14278 0 14334 800 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 520 nsew signal input
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 521 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 522 nsew signal input
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 523 nsew signal input
flabel metal2 s 15382 0 15438 800 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 524 nsew signal input
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 525 nsew signal input
flabel metal2 s 15934 0 15990 800 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 526 nsew signal input
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 527 nsew signal input
flabel metal2 s 16486 0 16542 800 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 528 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 529 nsew signal input
flabel metal2 s 11518 0 11574 800 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 530 nsew signal input
flabel metal2 s 17038 0 17094 800 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 531 nsew signal input
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 532 nsew signal input
flabel metal2 s 17590 0 17646 800 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 533 nsew signal input
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 534 nsew signal input
flabel metal2 s 18142 0 18198 800 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 535 nsew signal input
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 536 nsew signal input
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 537 nsew signal input
flabel metal2 s 18970 0 19026 800 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 538 nsew signal input
flabel metal2 s 19246 0 19302 800 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 539 nsew signal input
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 540 nsew signal input
flabel metal2 s 11886 0 11942 800 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 541 nsew signal input
flabel metal2 s 19798 0 19854 800 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 542 nsew signal input
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 543 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 544 nsew signal input
flabel metal2 s 12622 0 12678 800 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 545 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 546 nsew signal input
flabel metal2 s 13174 0 13230 800 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 547 nsew signal input
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 548 nsew signal input
flabel metal2 s 13726 0 13782 800 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 549 nsew signal input
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 550 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 551 nsew signal input
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 552 nsew signal input
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 553 nsew signal input
flabel metal2 s 14646 0 14702 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 554 nsew signal input
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 555 nsew signal input
flabel metal2 s 15198 0 15254 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 556 nsew signal input
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 557 nsew signal input
flabel metal2 s 15750 0 15806 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 558 nsew signal input
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 559 nsew signal input
flabel metal2 s 16302 0 16358 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 560 nsew signal input
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 561 nsew signal input
flabel metal2 s 16854 0 16910 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 562 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 563 nsew signal input
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 564 nsew signal input
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 565 nsew signal input
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 566 nsew signal input
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 567 nsew signal input
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 568 nsew signal input
flabel metal2 s 18510 0 18566 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 569 nsew signal input
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 570 nsew signal input
flabel metal2 s 19062 0 19118 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 571 nsew signal input
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 572 nsew signal input
flabel metal2 s 19614 0 19670 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 573 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 574 nsew signal input
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 575 nsew signal input
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 576 nsew signal input
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 577 nsew signal input
flabel metal2 s 12714 0 12770 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 578 nsew signal input
flabel metal2 s 12990 0 13046 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 579 nsew signal input
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 580 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 581 nsew signal input
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 582 nsew signal input
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 583 nsew signal input
flabel metal2 s 11334 0 11390 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 584 nsew signal tristate
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 585 nsew signal tristate
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 586 nsew signal tristate
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 587 nsew signal tristate
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 588 nsew signal tristate
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 589 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 590 nsew signal tristate
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 591 nsew signal tristate
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 592 nsew signal tristate
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 593 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 594 nsew signal tristate
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 595 nsew signal tristate
flabel metal2 s 17222 0 17278 800 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 596 nsew signal tristate
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 597 nsew signal tristate
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 598 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 599 nsew signal tristate
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 600 nsew signal tristate
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 601 nsew signal tristate
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 602 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 603 nsew signal tristate
flabel metal2 s 19430 0 19486 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 604 nsew signal tristate
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 605 nsew signal tristate
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 606 nsew signal tristate
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 607 nsew signal tristate
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 608 nsew signal tristate
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 609 nsew signal tristate
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 610 nsew signal tristate
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 611 nsew signal tristate
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 612 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 613 nsew signal tristate
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 614 nsew signal tristate
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 615 nsew signal tristate
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 wbs_sel_i[0]
port 616 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 wbs_sel_i[1]
port 617 nsew signal input
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 wbs_sel_i[2]
port 618 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 wbs_sel_i[3]
port 619 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 wbs_stb_i
port 620 nsew signal input
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 wbs_we_i
port 621 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 70000 60000
<< end >>
