magic
tech sky130B
magscale 1 2
timestamp 1668103391
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 196618 700612 196624 700664
rect 196676 700652 196682 700664
rect 218974 700652 218980 700664
rect 196676 700624 218980 700652
rect 196676 700612 196682 700624
rect 218974 700612 218980 700624
rect 219032 700612 219038 700664
rect 193858 700544 193864 700596
rect 193916 700584 193922 700596
rect 283834 700584 283840 700596
rect 193916 700556 283840 700584
rect 193916 700544 193922 700556
rect 283834 700544 283840 700556
rect 283892 700544 283898 700596
rect 192478 700476 192484 700528
rect 192536 700516 192542 700528
rect 348786 700516 348792 700528
rect 192536 700488 348792 700516
rect 192536 700476 192542 700488
rect 348786 700476 348792 700488
rect 348844 700476 348850 700528
rect 189718 700408 189724 700460
rect 189776 700448 189782 700460
rect 413646 700448 413652 700460
rect 189776 700420 413652 700448
rect 189776 700408 189782 700420
rect 413646 700408 413652 700420
rect 413704 700408 413710 700460
rect 188338 700340 188344 700392
rect 188396 700380 188402 700392
rect 478506 700380 478512 700392
rect 188396 700352 478512 700380
rect 188396 700340 188402 700352
rect 478506 700340 478512 700352
rect 478564 700340 478570 700392
rect 89162 700272 89168 700324
rect 89220 700312 89226 700324
rect 180794 700312 180800 700324
rect 89220 700284 180800 700312
rect 89220 700272 89226 700284
rect 180794 700272 180800 700284
rect 180852 700272 180858 700324
rect 185578 700272 185584 700324
rect 185636 700312 185642 700324
rect 543458 700312 543464 700324
rect 185636 700284 543464 700312
rect 185636 700272 185642 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106918 699700 106924 699712
rect 105504 699672 106924 699700
rect 105504 699660 105510 699672
rect 106918 699660 106924 699672
rect 106976 699660 106982 699712
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 2774 683680 2780 683732
rect 2832 683720 2838 683732
rect 4798 683720 4804 683732
rect 2832 683692 4804 683720
rect 2832 683680 2838 683692
rect 4798 683680 4804 683692
rect 4856 683680 4862 683732
rect 184198 683136 184204 683188
rect 184256 683176 184262 683188
rect 579614 683176 579620 683188
rect 184256 683148 579620 683176
rect 184256 683136 184262 683148
rect 579614 683136 579620 683148
rect 579672 683136 579678 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 180886 670732 180892 670744
rect 3568 670704 180892 670732
rect 3568 670692 3574 670704
rect 180886 670692 180892 670704
rect 180944 670692 180950 670744
rect 182818 643084 182824 643136
rect 182876 643124 182882 643136
rect 580166 643124 580172 643136
rect 182876 643096 580172 643124
rect 182876 643084 182882 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3510 632068 3516 632120
rect 3568 632108 3574 632120
rect 7558 632108 7564 632120
rect 3568 632080 7564 632108
rect 3568 632068 3574 632080
rect 7558 632068 7564 632080
rect 7616 632068 7622 632120
rect 184290 630640 184296 630692
rect 184348 630680 184354 630692
rect 579706 630680 579712 630692
rect 184348 630652 579712 630680
rect 184348 630640 184354 630652
rect 579706 630640 579712 630652
rect 579764 630640 579770 630692
rect 3510 618264 3516 618316
rect 3568 618304 3574 618316
rect 180978 618304 180984 618316
rect 3568 618276 180984 618304
rect 3568 618264 3574 618276
rect 180978 618264 180984 618276
rect 181036 618264 181042 618316
rect 120718 616836 120724 616888
rect 120776 616876 120782 616888
rect 580166 616876 580172 616888
rect 120776 616848 580172 616876
rect 120776 616836 120782 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3510 579640 3516 579692
rect 3568 579680 3574 579692
rect 17218 579680 17224 579692
rect 3568 579652 17224 579680
rect 3568 579640 3574 579652
rect 17218 579640 17224 579652
rect 17276 579640 17282 579692
rect 184382 576852 184388 576904
rect 184440 576892 184446 576904
rect 580166 576892 580172 576904
rect 184440 576864 580172 576892
rect 184440 576852 184446 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3050 565836 3056 565888
rect 3108 565876 3114 565888
rect 179414 565876 179420 565888
rect 3108 565848 179420 565876
rect 3108 565836 3114 565848
rect 179414 565836 179420 565848
rect 179472 565836 179478 565888
rect 120810 563048 120816 563100
rect 120868 563088 120874 563100
rect 580166 563088 580172 563100
rect 120868 563060 580172 563088
rect 120868 563048 120874 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 180058 536800 180064 536852
rect 180116 536840 180122 536852
rect 580166 536840 580172 536852
rect 180116 536812 580172 536840
rect 180116 536800 180122 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 3510 527824 3516 527876
rect 3568 527864 3574 527876
rect 8938 527864 8944 527876
rect 3568 527836 8944 527864
rect 3568 527824 3574 527836
rect 8938 527824 8944 527836
rect 8996 527824 9002 527876
rect 214558 524424 214564 524476
rect 214616 524464 214622 524476
rect 579798 524464 579804 524476
rect 214616 524436 579804 524464
rect 214616 524424 214622 524436
rect 579798 524424 579804 524436
rect 579856 524424 579862 524476
rect 3510 514768 3516 514820
rect 3568 514808 3574 514820
rect 181070 514808 181076 514820
rect 3568 514780 181076 514808
rect 3568 514768 3574 514780
rect 181070 514768 181076 514780
rect 181128 514768 181134 514820
rect 120902 510620 120908 510672
rect 120960 510660 120966 510672
rect 579982 510660 579988 510672
rect 120960 510632 579988 510660
rect 120960 510620 120966 510632
rect 579982 510620 579988 510632
rect 580040 510620 580046 510672
rect 182910 484372 182916 484424
rect 182968 484412 182974 484424
rect 580166 484412 580172 484424
rect 182968 484384 580172 484412
rect 182968 484372 182974 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 3510 474716 3516 474768
rect 3568 474756 3574 474768
rect 10318 474756 10324 474768
rect 3568 474728 10324 474756
rect 3568 474716 3574 474728
rect 10318 474716 10324 474728
rect 10376 474716 10382 474768
rect 211798 470568 211804 470620
rect 211856 470608 211862 470620
rect 579614 470608 579620 470620
rect 211856 470580 579620 470608
rect 211856 470568 211862 470580
rect 579614 470568 579620 470580
rect 579672 470568 579678 470620
rect 120994 456764 121000 456816
rect 121052 456804 121058 456816
rect 579614 456804 579620 456816
rect 121052 456776 579620 456804
rect 121052 456764 121058 456776
rect 579614 456764 579620 456776
rect 579672 456764 579678 456816
rect 118694 431196 118700 431248
rect 118752 431236 118758 431248
rect 580534 431236 580540 431248
rect 118752 431208 580540 431236
rect 118752 431196 118758 431208
rect 580534 431196 580540 431208
rect 580592 431196 580598 431248
rect 2958 422288 2964 422340
rect 3016 422328 3022 422340
rect 13078 422328 13084 422340
rect 3016 422300 13084 422328
rect 3016 422288 3022 422300
rect 13078 422288 13084 422300
rect 13136 422288 13142 422340
rect 183002 418140 183008 418192
rect 183060 418180 183066 418192
rect 580166 418180 580172 418192
rect 183060 418152 580172 418180
rect 183060 418140 183066 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 3050 409844 3056 409896
rect 3108 409884 3114 409896
rect 179506 409884 179512 409896
rect 3108 409856 179512 409884
rect 3108 409844 3114 409856
rect 179506 409844 179512 409856
rect 179564 409844 179570 409896
rect 118602 404336 118608 404388
rect 118660 404376 118666 404388
rect 580166 404376 580172 404388
rect 118660 404348 580172 404376
rect 118660 404336 118666 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3326 371220 3332 371272
rect 3384 371260 3390 371272
rect 84838 371260 84844 371272
rect 3384 371232 84844 371260
rect 3384 371220 3390 371232
rect 84838 371220 84844 371232
rect 84896 371220 84902 371272
rect 224218 364352 224224 364404
rect 224276 364392 224282 364404
rect 580166 364392 580172 364404
rect 224276 364364 580172 364392
rect 224276 364352 224282 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 3326 357416 3332 357468
rect 3384 357456 3390 357468
rect 181162 357456 181168 357468
rect 3384 357428 181168 357456
rect 3384 357416 3390 357428
rect 181162 357416 181168 357428
rect 181220 357416 181226 357468
rect 118510 351908 118516 351960
rect 118568 351948 118574 351960
rect 580166 351948 580172 351960
rect 118568 351920 580172 351948
rect 118568 351908 118574 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 3326 318792 3332 318844
rect 3384 318832 3390 318844
rect 14458 318832 14464 318844
rect 3384 318804 14464 318832
rect 3384 318792 3390 318804
rect 14458 318792 14464 318804
rect 14516 318792 14522 318844
rect 221458 311856 221464 311908
rect 221516 311896 221522 311908
rect 580166 311896 580172 311908
rect 221516 311868 580172 311896
rect 221516 311856 221522 311868
rect 580166 311856 580172 311868
rect 580224 311856 580230 311908
rect 3326 304988 3332 305040
rect 3384 305028 3390 305040
rect 182174 305028 182180 305040
rect 3384 305000 182180 305028
rect 3384 304988 3390 305000
rect 182174 304988 182180 305000
rect 182232 304988 182238 305040
rect 146938 298120 146944 298172
rect 146996 298160 147002 298172
rect 580166 298160 580172 298172
rect 146996 298132 580172 298160
rect 146996 298120 147002 298132
rect 580166 298120 580172 298132
rect 580224 298120 580230 298172
rect 183094 271872 183100 271924
rect 183152 271912 183158 271924
rect 580166 271912 580172 271924
rect 183152 271884 580172 271912
rect 183152 271872 183158 271884
rect 580166 271872 580172 271884
rect 580224 271872 580230 271924
rect 3326 266364 3332 266416
rect 3384 266404 3390 266416
rect 18598 266404 18604 266416
rect 3384 266376 18604 266404
rect 3384 266364 3390 266376
rect 18598 266364 18604 266376
rect 18656 266364 18662 266416
rect 220078 258068 220084 258120
rect 220136 258108 220142 258120
rect 579614 258108 579620 258120
rect 220136 258080 579620 258108
rect 220136 258068 220142 258080
rect 579614 258068 579620 258080
rect 579672 258068 579678 258120
rect 3326 253920 3332 253972
rect 3384 253960 3390 253972
rect 178678 253960 178684 253972
rect 3384 253932 178684 253960
rect 3384 253920 3390 253932
rect 178678 253920 178684 253932
rect 178736 253920 178742 253972
rect 126238 244264 126244 244316
rect 126296 244304 126302 244316
rect 580166 244304 580172 244316
rect 126296 244276 580172 244304
rect 126296 244264 126302 244276
rect 580166 244264 580172 244276
rect 580224 244264 580230 244316
rect 3326 240116 3332 240168
rect 3384 240156 3390 240168
rect 82078 240156 82084 240168
rect 3384 240128 82084 240156
rect 3384 240116 3390 240128
rect 82078 240116 82084 240128
rect 82136 240116 82142 240168
rect 217318 218016 217324 218068
rect 217376 218056 217382 218068
rect 580166 218056 580172 218068
rect 217376 218028 580172 218056
rect 217376 218016 217382 218028
rect 580166 218016 580172 218028
rect 580224 218016 580230 218068
rect 3326 213936 3332 213988
rect 3384 213976 3390 213988
rect 31018 213976 31024 213988
rect 3384 213948 31024 213976
rect 3384 213936 3390 213948
rect 31018 213936 31024 213948
rect 31076 213936 31082 213988
rect 122098 205640 122104 205692
rect 122156 205680 122162 205692
rect 580166 205680 580172 205692
rect 122156 205652 580172 205680
rect 122156 205640 122162 205652
rect 580166 205640 580172 205652
rect 580224 205640 580230 205692
rect 3326 201492 3332 201544
rect 3384 201532 3390 201544
rect 178770 201532 178776 201544
rect 3384 201504 178776 201532
rect 3384 201492 3390 201504
rect 178770 201492 178776 201504
rect 178828 201492 178834 201544
rect 3326 187688 3332 187740
rect 3384 187728 3390 187740
rect 119338 187728 119344 187740
rect 3384 187700 119344 187728
rect 3384 187688 3390 187700
rect 119338 187688 119344 187700
rect 119396 187688 119402 187740
rect 215938 178032 215944 178084
rect 215996 178072 216002 178084
rect 580166 178072 580172 178084
rect 215996 178044 580172 178072
rect 215996 178032 216002 178044
rect 580166 178032 580172 178044
rect 580224 178032 580230 178084
rect 3510 166268 3516 166320
rect 3568 166308 3574 166320
rect 179690 166308 179696 166320
rect 3568 166280 179696 166308
rect 3568 166268 3574 166280
rect 179690 166268 179696 166280
rect 179748 166268 179754 166320
rect 122190 165588 122196 165640
rect 122248 165628 122254 165640
rect 580166 165628 580172 165640
rect 122248 165600 580172 165628
rect 122248 165588 122254 165600
rect 580166 165588 580172 165600
rect 580224 165588 580230 165640
rect 3510 162868 3516 162920
rect 3568 162908 3574 162920
rect 21358 162908 21364 162920
rect 3568 162880 21364 162908
rect 3568 162868 3574 162880
rect 21358 162868 21364 162880
rect 21416 162868 21422 162920
rect 183186 151784 183192 151836
rect 183244 151824 183250 151836
rect 579982 151824 579988 151836
rect 183244 151796 579988 151824
rect 183244 151784 183250 151796
rect 579982 151784 579988 151796
rect 580040 151784 580046 151836
rect 3510 149064 3516 149116
rect 3568 149104 3574 149116
rect 179598 149104 179604 149116
rect 3568 149076 179604 149104
rect 3568 149064 3574 149076
rect 179598 149064 179604 149076
rect 179656 149064 179662 149116
rect 119062 145596 119068 145648
rect 119120 145636 119126 145648
rect 234614 145636 234620 145648
rect 119120 145608 234620 145636
rect 119120 145596 119126 145608
rect 234614 145596 234620 145608
rect 234672 145596 234678 145648
rect 23474 145528 23480 145580
rect 23532 145568 23538 145580
rect 179782 145568 179788 145580
rect 23532 145540 179788 145568
rect 23532 145528 23538 145540
rect 179782 145528 179788 145540
rect 179840 145528 179846 145580
rect 119154 144168 119160 144220
rect 119212 144208 119218 144220
rect 299474 144208 299480 144220
rect 119212 144180 299480 144208
rect 119212 144168 119218 144180
rect 299474 144168 299480 144180
rect 299532 144168 299538 144220
rect 118234 142876 118240 142928
rect 118292 142916 118298 142928
rect 146938 142916 146944 142928
rect 118292 142888 146944 142916
rect 118292 142876 118298 142888
rect 146938 142876 146944 142888
rect 146996 142876 147002 142928
rect 153194 142876 153200 142928
rect 153252 142916 153258 142928
rect 181438 142916 181444 142928
rect 153252 142888 181444 142916
rect 153252 142876 153258 142888
rect 181438 142876 181444 142888
rect 181496 142876 181502 142928
rect 118970 142808 118976 142860
rect 119028 142848 119034 142860
rect 429194 142848 429200 142860
rect 119028 142820 429200 142848
rect 119028 142808 119034 142820
rect 429194 142808 429200 142820
rect 429252 142808 429258 142860
rect 118142 141516 118148 141568
rect 118200 141556 118206 141568
rect 126238 141556 126244 141568
rect 118200 141528 126244 141556
rect 118200 141516 118206 141528
rect 126238 141516 126244 141528
rect 126296 141516 126302 141568
rect 136634 141516 136640 141568
rect 136692 141556 136698 141568
rect 181346 141556 181352 141568
rect 136692 141528 181352 141556
rect 136692 141516 136698 141528
rect 181346 141516 181352 141528
rect 181404 141516 181410 141568
rect 118050 141448 118056 141500
rect 118108 141488 118114 141500
rect 169754 141488 169760 141500
rect 118108 141460 169760 141488
rect 118108 141448 118114 141460
rect 169754 141448 169760 141460
rect 169812 141448 169818 141500
rect 118878 141380 118884 141432
rect 118936 141420 118942 141432
rect 494054 141420 494060 141432
rect 118936 141392 494060 141420
rect 118936 141380 118942 141392
rect 494054 141380 494060 141392
rect 494112 141380 494118 141432
rect 119246 140088 119252 140140
rect 119304 140128 119310 140140
rect 364334 140128 364340 140140
rect 119304 140100 364340 140128
rect 119304 140088 119310 140100
rect 364334 140088 364340 140100
rect 364392 140088 364398 140140
rect 118786 140020 118792 140072
rect 118844 140060 118850 140072
rect 558914 140060 558920 140072
rect 118844 140032 558920 140060
rect 118844 140020 118850 140032
rect 558914 140020 558920 140032
rect 558972 140020 558978 140072
rect 118326 139544 118332 139596
rect 118384 139584 118390 139596
rect 122098 139584 122104 139596
rect 118384 139556 122104 139584
rect 118384 139544 118390 139556
rect 122098 139544 122104 139556
rect 122156 139544 122162 139596
rect 118418 139476 118424 139528
rect 118476 139516 118482 139528
rect 122190 139516 122196 139528
rect 118476 139488 122196 139516
rect 118476 139476 118482 139488
rect 122190 139476 122196 139488
rect 122248 139476 122254 139528
rect 3326 139408 3332 139460
rect 3384 139448 3390 139460
rect 181530 139448 181536 139460
rect 3384 139420 181536 139448
rect 3384 139408 3390 139420
rect 181530 139408 181536 139420
rect 181588 139408 181594 139460
rect 178678 139340 178684 139392
rect 178736 139380 178742 139392
rect 182266 139380 182272 139392
rect 178736 139352 182272 139380
rect 178736 139340 178742 139352
rect 182266 139340 182272 139352
rect 182324 139340 182330 139392
rect 178770 139272 178776 139324
rect 178828 139312 178834 139324
rect 182358 139312 182364 139324
rect 178828 139284 182364 139312
rect 178828 139272 178834 139284
rect 182358 139272 182364 139284
rect 182416 139272 182422 139324
rect 196710 137980 196716 138032
rect 196768 138020 196774 138032
rect 580166 138020 580172 138032
rect 196768 137992 580172 138020
rect 196768 137980 196774 137992
rect 580166 137980 580172 137992
rect 580224 137980 580230 138032
rect 3510 137776 3516 137828
rect 3568 137816 3574 137828
rect 121086 137816 121092 137828
rect 3568 137788 121092 137816
rect 3568 137776 3574 137788
rect 121086 137776 121092 137788
rect 121144 137776 121150 137828
rect 7650 136688 7656 136740
rect 7708 136728 7714 136740
rect 117314 136728 117320 136740
rect 7708 136700 117320 136728
rect 7708 136688 7714 136700
rect 117314 136688 117320 136700
rect 117372 136688 117378 136740
rect 9030 135260 9036 135312
rect 9088 135300 9094 135312
rect 117314 135300 117320 135312
rect 9088 135272 117320 135300
rect 9088 135260 9094 135272
rect 117314 135260 117320 135272
rect 117372 135260 117378 135312
rect 3418 135056 3424 135108
rect 3476 135056 3482 135108
rect 3436 134904 3464 135056
rect 3418 134852 3424 134904
rect 3476 134852 3482 134904
rect 22738 133900 22744 133952
rect 22796 133940 22802 133952
rect 117314 133940 117320 133952
rect 22796 133912 117320 133940
rect 22796 133900 22802 133912
rect 117314 133900 117320 133912
rect 117372 133900 117378 133952
rect 21358 133832 21364 133884
rect 21416 133872 21422 133884
rect 117406 133872 117412 133884
rect 21416 133844 117412 133872
rect 21416 133832 21422 133844
rect 117406 133832 117412 133844
rect 117464 133832 117470 133884
rect 31018 132404 31024 132456
rect 31076 132444 31082 132456
rect 117314 132444 117320 132456
rect 31076 132416 117320 132444
rect 31076 132404 31082 132416
rect 117314 132404 117320 132416
rect 117372 132404 117378 132456
rect 18598 131044 18604 131096
rect 18656 131084 18662 131096
rect 117314 131084 117320 131096
rect 18656 131056 117320 131084
rect 18656 131044 18662 131056
rect 117314 131044 117320 131056
rect 117372 131044 117378 131096
rect 14458 129684 14464 129736
rect 14516 129724 14522 129736
rect 117314 129724 117320 129736
rect 14516 129696 117320 129724
rect 14516 129684 14522 129696
rect 117314 129684 117320 129696
rect 117372 129684 117378 129736
rect 84838 128256 84844 128308
rect 84896 128296 84902 128308
rect 117314 128296 117320 128308
rect 84896 128268 117320 128296
rect 84896 128256 84902 128268
rect 117314 128256 117320 128268
rect 117372 128256 117378 128308
rect 13078 126896 13084 126948
rect 13136 126936 13142 126948
rect 117314 126936 117320 126948
rect 13136 126908 117320 126936
rect 13136 126896 13142 126908
rect 117314 126896 117320 126908
rect 117372 126896 117378 126948
rect 10318 124108 10324 124160
rect 10376 124148 10382 124160
rect 117314 124148 117320 124160
rect 10376 124120 117320 124148
rect 10376 124108 10382 124120
rect 117314 124108 117320 124120
rect 117372 124108 117378 124160
rect 8938 122748 8944 122800
rect 8996 122788 9002 122800
rect 117314 122788 117320 122800
rect 8996 122760 117320 122788
rect 8996 122748 9002 122760
rect 117314 122748 117320 122760
rect 117372 122748 117378 122800
rect 17218 121388 17224 121440
rect 17276 121428 17282 121440
rect 117314 121428 117320 121440
rect 17276 121400 117320 121428
rect 17276 121388 17282 121400
rect 117314 121388 117320 121400
rect 117372 121388 117378 121440
rect 7558 120028 7564 120080
rect 7616 120068 7622 120080
rect 117314 120068 117320 120080
rect 7616 120040 117320 120068
rect 7616 120028 7622 120040
rect 117314 120028 117320 120040
rect 117372 120028 117378 120080
rect 4798 118600 4804 118652
rect 4856 118640 4862 118652
rect 117314 118640 117320 118652
rect 4856 118612 117320 118640
rect 4856 118600 4862 118612
rect 117314 118600 117320 118612
rect 117372 118600 117378 118652
rect 40034 117240 40040 117292
rect 40092 117280 40098 117292
rect 117314 117280 117320 117292
rect 40092 117252 117320 117280
rect 40092 117240 40098 117252
rect 117314 117240 117320 117252
rect 117372 117240 117378 117292
rect 106918 115880 106924 115932
rect 106976 115920 106982 115932
rect 117314 115920 117320 115932
rect 106976 115892 117320 115920
rect 106976 115880 106982 115892
rect 117314 115880 117320 115892
rect 117372 115880 117378 115932
rect 180150 111800 180156 111852
rect 180208 111840 180214 111852
rect 579982 111840 579988 111852
rect 180208 111812 579988 111840
rect 180208 111800 180214 111812
rect 579982 111800 579988 111812
rect 580040 111800 580046 111852
rect 3326 111732 3332 111784
rect 3384 111772 3390 111784
rect 22738 111772 22744 111784
rect 3384 111744 22744 111772
rect 3384 111732 3390 111744
rect 22738 111732 22744 111744
rect 22796 111732 22802 111784
rect 183462 108944 183468 108996
rect 183520 108984 183526 108996
rect 196618 108984 196624 108996
rect 183520 108956 196624 108984
rect 183520 108944 183526 108956
rect 196618 108944 196624 108956
rect 196676 108944 196682 108996
rect 183462 107584 183468 107636
rect 183520 107624 183526 107636
rect 193858 107624 193864 107636
rect 183520 107596 193864 107624
rect 183520 107584 183526 107596
rect 193858 107584 193864 107596
rect 193916 107584 193922 107636
rect 183462 106224 183468 106276
rect 183520 106264 183526 106276
rect 192478 106264 192484 106276
rect 183520 106236 192484 106264
rect 183520 106224 183526 106236
rect 192478 106224 192484 106236
rect 192536 106224 192542 106276
rect 182726 104796 182732 104848
rect 182784 104836 182790 104848
rect 189718 104836 189724 104848
rect 182784 104808 189724 104836
rect 182784 104796 182790 104808
rect 189718 104796 189724 104808
rect 189776 104796 189782 104848
rect 183462 102620 183468 102672
rect 183520 102660 183526 102672
rect 188338 102660 188344 102672
rect 183520 102632 188344 102660
rect 183520 102620 183526 102632
rect 188338 102620 188344 102632
rect 188396 102620 188402 102672
rect 182266 101464 182272 101516
rect 182324 101504 182330 101516
rect 185578 101504 185584 101516
rect 182324 101476 185584 101504
rect 182324 101464 182330 101476
rect 185578 101464 185584 101476
rect 185636 101464 185642 101516
rect 182450 99968 182456 100020
rect 182508 100008 182514 100020
rect 184198 100008 184204 100020
rect 182508 99980 184204 100008
rect 182508 99968 182514 99980
rect 184198 99968 184204 99980
rect 184256 99968 184262 100020
rect 193858 99356 193864 99408
rect 193916 99396 193922 99408
rect 580166 99396 580172 99408
rect 193916 99368 580172 99396
rect 193916 99356 193922 99368
rect 580166 99356 580172 99368
rect 580224 99356 580230 99408
rect 182174 98472 182180 98524
rect 182232 98512 182238 98524
rect 184290 98512 184296 98524
rect 182232 98484 184296 98512
rect 182232 98472 182238 98484
rect 184290 98472 184296 98484
rect 184348 98472 184354 98524
rect 182542 97384 182548 97436
rect 182600 97424 182606 97436
rect 184382 97424 184388 97436
rect 182600 97396 184388 97424
rect 182600 97384 182606 97396
rect 184382 97384 184388 97396
rect 184440 97384 184446 97436
rect 183462 96568 183468 96620
rect 183520 96608 183526 96620
rect 214558 96608 214564 96620
rect 183520 96580 214564 96608
rect 183520 96568 183526 96580
rect 214558 96568 214564 96580
rect 214616 96568 214622 96620
rect 183462 95140 183468 95192
rect 183520 95180 183526 95192
rect 211798 95180 211804 95192
rect 183520 95152 211804 95180
rect 183520 95140 183526 95152
rect 211798 95140 211804 95152
rect 211856 95140 211862 95192
rect 182542 93100 182548 93152
rect 182600 93140 182606 93152
rect 224218 93140 224224 93152
rect 182600 93112 224224 93140
rect 182600 93100 182606 93112
rect 224218 93100 224224 93112
rect 224276 93100 224282 93152
rect 183462 91740 183468 91792
rect 183520 91780 183526 91792
rect 221458 91780 221464 91792
rect 183520 91752 221464 91780
rect 183520 91740 183526 91752
rect 221458 91740 221464 91752
rect 221516 91740 221522 91792
rect 183370 90312 183376 90364
rect 183428 90352 183434 90364
rect 220078 90352 220084 90364
rect 183428 90324 220084 90352
rect 183428 90312 183434 90324
rect 220078 90312 220084 90324
rect 220136 90312 220142 90364
rect 580166 89088 580172 89140
rect 580224 89128 580230 89140
rect 580626 89128 580632 89140
rect 580224 89100 580632 89128
rect 580224 89088 580230 89100
rect 580626 89088 580632 89100
rect 580684 89088 580690 89140
rect 183462 88952 183468 89004
rect 183520 88992 183526 89004
rect 217318 88992 217324 89004
rect 183520 88964 217324 88992
rect 183520 88952 183526 88964
rect 217318 88952 217324 88964
rect 217376 88952 217382 89004
rect 580626 88952 580632 89004
rect 580684 88992 580690 89004
rect 580902 88992 580908 89004
rect 580684 88964 580908 88992
rect 580684 88952 580690 88964
rect 580902 88952 580908 88964
rect 580960 88952 580966 89004
rect 183370 87592 183376 87644
rect 183428 87632 183434 87644
rect 215938 87632 215944 87644
rect 183428 87604 215944 87632
rect 183428 87592 183434 87604
rect 215938 87592 215944 87604
rect 215996 87592 216002 87644
rect 183462 85484 183468 85536
rect 183520 85524 183526 85536
rect 196710 85524 196716 85536
rect 183520 85496 196716 85524
rect 183520 85484 183526 85496
rect 196710 85484 196716 85496
rect 196768 85484 196774 85536
rect 3510 84192 3516 84244
rect 3568 84232 3574 84244
rect 120718 84232 120724 84244
rect 3568 84204 120724 84232
rect 3568 84192 3574 84204
rect 120718 84192 120724 84204
rect 120776 84192 120782 84244
rect 183462 84124 183468 84176
rect 183520 84164 183526 84176
rect 193858 84164 193864 84176
rect 183520 84136 193864 84164
rect 183520 84124 183526 84136
rect 193858 84124 193864 84136
rect 193916 84124 193922 84176
rect 120902 80792 120908 80844
rect 120960 80832 120966 80844
rect 580350 80832 580356 80844
rect 120960 80804 136634 80832
rect 120960 80792 120966 80804
rect 127222 80736 127526 80764
rect 122098 80588 122104 80640
rect 122156 80628 122162 80640
rect 127222 80628 127250 80736
rect 122156 80600 127250 80628
rect 122156 80588 122162 80600
rect 127498 80220 127526 80736
rect 136606 80628 136634 80804
rect 137986 80804 139394 80832
rect 137986 80628 138014 80804
rect 139366 80764 139394 80804
rect 169726 80804 174216 80832
rect 169726 80764 169754 80804
rect 139366 80736 140774 80764
rect 136606 80600 138014 80628
rect 140746 80628 140774 80736
rect 162964 80736 169754 80764
rect 169864 80736 173204 80764
rect 162964 80696 162992 80736
rect 144886 80668 162992 80696
rect 144886 80628 144914 80668
rect 169864 80628 169892 80736
rect 140746 80600 144914 80628
rect 154638 80600 169892 80628
rect 150728 80532 153976 80560
rect 150728 80492 150756 80532
rect 150406 80464 150756 80492
rect 137986 80396 139394 80424
rect 137986 80220 138014 80396
rect 139366 80356 139394 80396
rect 150406 80356 150434 80464
rect 139366 80328 140774 80356
rect 127498 80192 138014 80220
rect 140746 80220 140774 80328
rect 149026 80328 150434 80356
rect 143506 80260 144914 80288
rect 143506 80220 143534 80260
rect 140746 80192 143534 80220
rect 144886 80220 144914 80260
rect 149026 80220 149054 80328
rect 144886 80192 149054 80220
rect 125658 80124 133046 80152
rect 6914 79976 6920 80028
rect 6972 80016 6978 80028
rect 122098 80016 122104 80028
rect 6972 79988 122104 80016
rect 6972 79976 6978 79988
rect 122098 79976 122104 79988
rect 122156 79976 122162 80028
rect 125226 79908 125232 79960
rect 125284 79948 125290 79960
rect 125658 79948 125686 80124
rect 129614 79988 130286 80016
rect 125284 79920 125686 79948
rect 125284 79908 125290 79920
rect 125824 79908 125830 79960
rect 125882 79908 125888 79960
rect 126560 79908 126566 79960
rect 126618 79908 126624 79960
rect 126652 79908 126658 79960
rect 126710 79908 126716 79960
rect 126928 79948 126934 79960
rect 126900 79908 126934 79948
rect 126986 79908 126992 79960
rect 127020 79908 127026 79960
rect 127078 79908 127084 79960
rect 127388 79908 127394 79960
rect 127446 79908 127452 79960
rect 127480 79908 127486 79960
rect 127538 79908 127544 79960
rect 127664 79948 127670 79960
rect 127590 79920 127670 79948
rect 125842 79824 125870 79908
rect 126008 79840 126014 79892
rect 126066 79840 126072 79892
rect 125842 79784 125876 79824
rect 125870 79772 125876 79784
rect 125928 79772 125934 79824
rect 126026 79756 126054 79840
rect 126100 79772 126106 79824
rect 126158 79772 126164 79824
rect 82078 79704 82084 79756
rect 82136 79744 82142 79756
rect 120902 79744 120908 79756
rect 82136 79716 120908 79744
rect 82136 79704 82142 79716
rect 120902 79704 120908 79716
rect 120960 79704 120966 79756
rect 125962 79704 125968 79756
rect 126020 79716 126054 79756
rect 126020 79704 126026 79716
rect 118666 79648 123616 79676
rect 3694 79568 3700 79620
rect 3752 79608 3758 79620
rect 118666 79608 118694 79648
rect 3752 79580 118694 79608
rect 123588 79608 123616 79648
rect 125134 79636 125140 79688
rect 125192 79676 125198 79688
rect 126118 79676 126146 79772
rect 125192 79648 126146 79676
rect 125192 79636 125198 79648
rect 125778 79608 125784 79620
rect 123588 79580 125784 79608
rect 3752 79568 3758 79580
rect 125778 79568 125784 79580
rect 125836 79568 125842 79620
rect 126578 79552 126606 79908
rect 126670 79620 126698 79908
rect 126900 79824 126928 79908
rect 127038 79824 127066 79908
rect 126744 79772 126750 79824
rect 126802 79772 126808 79824
rect 126882 79772 126888 79824
rect 126940 79772 126946 79824
rect 126974 79772 126980 79824
rect 127032 79784 127066 79824
rect 127032 79772 127038 79784
rect 126762 79688 126790 79772
rect 126762 79648 126796 79688
rect 126790 79636 126796 79648
rect 126848 79636 126854 79688
rect 127406 79620 127434 79908
rect 126670 79580 126704 79620
rect 126698 79568 126704 79580
rect 126756 79568 126762 79620
rect 127342 79568 127348 79620
rect 127400 79580 127434 79620
rect 127400 79568 127406 79580
rect 127498 79552 127526 79908
rect 127590 79608 127618 79920
rect 127664 79908 127670 79920
rect 127722 79908 127728 79960
rect 127756 79908 127762 79960
rect 127814 79908 127820 79960
rect 127848 79908 127854 79960
rect 127906 79908 127912 79960
rect 128308 79948 128314 79960
rect 128096 79920 128314 79948
rect 127774 79880 127802 79908
rect 127728 79852 127802 79880
rect 127728 79744 127756 79852
rect 127866 79824 127894 79908
rect 127802 79772 127808 79824
rect 127860 79784 127894 79824
rect 127860 79772 127866 79784
rect 127894 79744 127900 79756
rect 127728 79716 127900 79744
rect 127894 79704 127900 79716
rect 127952 79704 127958 79756
rect 127590 79580 127664 79608
rect 127636 79552 127664 79580
rect 126578 79512 126612 79552
rect 126606 79500 126612 79512
rect 126664 79500 126670 79552
rect 127434 79500 127440 79552
rect 127492 79512 127526 79552
rect 127492 79500 127498 79512
rect 127618 79500 127624 79552
rect 127676 79500 127682 79552
rect 128096 79484 128124 79920
rect 128308 79908 128314 79920
rect 128366 79908 128372 79960
rect 128400 79908 128406 79960
rect 128458 79908 128464 79960
rect 129044 79908 129050 79960
rect 129102 79908 129108 79960
rect 129136 79908 129142 79960
rect 129194 79908 129200 79960
rect 129412 79908 129418 79960
rect 129470 79908 129476 79960
rect 128216 79840 128222 79892
rect 128274 79840 128280 79892
rect 128234 79484 128262 79840
rect 128418 79756 128446 79908
rect 128584 79772 128590 79824
rect 128642 79772 128648 79824
rect 128354 79704 128360 79756
rect 128412 79716 128446 79756
rect 128412 79704 128418 79716
rect 128602 79688 128630 79772
rect 129062 79756 129090 79908
rect 128998 79704 129004 79756
rect 129056 79716 129090 79756
rect 129056 79704 129062 79716
rect 128602 79648 128636 79688
rect 128630 79636 128636 79648
rect 128688 79636 128694 79688
rect 128814 79636 128820 79688
rect 128872 79676 128878 79688
rect 129154 79676 129182 79908
rect 129228 79840 129234 79892
rect 129286 79840 129292 79892
rect 128872 79648 129182 79676
rect 128872 79636 128878 79648
rect 129246 79608 129274 79840
rect 129430 79688 129458 79908
rect 129430 79648 129464 79688
rect 129458 79636 129464 79648
rect 129516 79636 129522 79688
rect 129366 79608 129372 79620
rect 129246 79580 129372 79608
rect 129366 79568 129372 79580
rect 129424 79568 129430 79620
rect 129614 79540 129642 79988
rect 130258 79960 130286 79988
rect 132098 79988 132218 80016
rect 129780 79908 129786 79960
rect 129838 79908 129844 79960
rect 129890 79920 130102 79948
rect 129798 79688 129826 79908
rect 129734 79636 129740 79688
rect 129792 79648 129826 79688
rect 129792 79636 129798 79648
rect 129890 79608 129918 79920
rect 130074 79892 130102 79920
rect 130240 79908 130246 79960
rect 130298 79908 130304 79960
rect 130516 79948 130522 79960
rect 130350 79920 130522 79948
rect 129964 79840 129970 79892
rect 130022 79840 130028 79892
rect 130056 79840 130062 79892
rect 130114 79840 130120 79892
rect 130148 79840 130154 79892
rect 130206 79840 130212 79892
rect 129982 79688 130010 79840
rect 129982 79648 130016 79688
rect 130010 79636 130016 79648
rect 130068 79636 130074 79688
rect 130166 79676 130194 79840
rect 130166 79648 130240 79676
rect 130212 79620 130240 79648
rect 130102 79608 130108 79620
rect 129890 79580 130108 79608
rect 130102 79568 130108 79580
rect 130160 79568 130166 79620
rect 130194 79568 130200 79620
rect 130252 79568 130258 79620
rect 129476 79512 129642 79540
rect 128078 79432 128084 79484
rect 128136 79432 128142 79484
rect 128170 79432 128176 79484
rect 128228 79444 128262 79484
rect 128228 79432 128234 79444
rect 128906 79432 128912 79484
rect 128964 79472 128970 79484
rect 129476 79472 129504 79512
rect 130350 79472 130378 79920
rect 130516 79908 130522 79920
rect 130574 79908 130580 79960
rect 130792 79908 130798 79960
rect 130850 79908 130856 79960
rect 130884 79908 130890 79960
rect 130942 79908 130948 79960
rect 131160 79948 131166 79960
rect 131132 79908 131166 79948
rect 131218 79908 131224 79960
rect 131252 79908 131258 79960
rect 131310 79908 131316 79960
rect 131436 79908 131442 79960
rect 131494 79908 131500 79960
rect 131528 79908 131534 79960
rect 131586 79908 131592 79960
rect 131988 79908 131994 79960
rect 132046 79908 132052 79960
rect 130608 79840 130614 79892
rect 130666 79840 130672 79892
rect 130470 79636 130476 79688
rect 130528 79676 130534 79688
rect 130626 79676 130654 79840
rect 130528 79648 130654 79676
rect 130528 79636 130534 79648
rect 130810 79608 130838 79908
rect 130902 79756 130930 79908
rect 130976 79840 130982 79892
rect 131034 79880 131040 79892
rect 131034 79840 131068 79880
rect 130902 79716 130936 79756
rect 130930 79704 130936 79716
rect 130988 79704 130994 79756
rect 131040 79676 131068 79840
rect 131132 79688 131160 79908
rect 130580 79580 130838 79608
rect 130902 79648 131068 79676
rect 130580 79552 130608 79580
rect 130562 79500 130568 79552
rect 130620 79500 130626 79552
rect 130746 79500 130752 79552
rect 130804 79540 130810 79552
rect 130902 79540 130930 79648
rect 131114 79636 131120 79688
rect 131172 79636 131178 79688
rect 130804 79512 130930 79540
rect 130804 79500 130810 79512
rect 128964 79444 129504 79472
rect 129660 79444 130378 79472
rect 128964 79432 128970 79444
rect 118666 79376 128492 79404
rect 3878 79296 3884 79348
rect 3936 79336 3942 79348
rect 118666 79336 118694 79376
rect 3936 79308 118694 79336
rect 3936 79296 3942 79308
rect 124398 79296 124404 79348
rect 124456 79336 124462 79348
rect 127710 79336 127716 79348
rect 124456 79308 127716 79336
rect 124456 79296 124462 79308
rect 127710 79296 127716 79308
rect 127768 79296 127774 79348
rect 128464 79336 128492 79376
rect 128538 79364 128544 79416
rect 128596 79404 128602 79416
rect 129660 79404 129688 79444
rect 130930 79432 130936 79484
rect 130988 79472 130994 79484
rect 131270 79472 131298 79908
rect 131454 79824 131482 79908
rect 131436 79772 131442 79824
rect 131494 79772 131500 79824
rect 131546 79744 131574 79908
rect 131804 79772 131810 79824
rect 131862 79772 131868 79824
rect 131896 79772 131902 79824
rect 131954 79772 131960 79824
rect 131408 79716 131574 79744
rect 131408 79620 131436 79716
rect 131822 79620 131850 79772
rect 131390 79568 131396 79620
rect 131448 79568 131454 79620
rect 131666 79608 131672 79620
rect 131592 79580 131672 79608
rect 131592 79552 131620 79580
rect 131666 79568 131672 79580
rect 131724 79568 131730 79620
rect 131758 79568 131764 79620
rect 131816 79580 131850 79620
rect 131816 79568 131822 79580
rect 131574 79500 131580 79552
rect 131632 79500 131638 79552
rect 130988 79444 131298 79472
rect 130988 79432 130994 79444
rect 131666 79432 131672 79484
rect 131724 79472 131730 79484
rect 131914 79472 131942 79772
rect 132006 79688 132034 79908
rect 132098 79744 132126 79988
rect 132190 79960 132218 79988
rect 133018 79960 133046 80124
rect 143874 80124 147674 80152
rect 137434 80056 142660 80084
rect 133110 79988 133874 80016
rect 132172 79908 132178 79960
rect 132230 79908 132236 79960
rect 132908 79948 132914 79960
rect 132512 79920 132914 79948
rect 132264 79840 132270 79892
rect 132322 79880 132328 79892
rect 132322 79840 132356 79880
rect 132328 79756 132356 79840
rect 132098 79716 132264 79744
rect 132006 79648 132040 79688
rect 132034 79636 132040 79648
rect 132092 79636 132098 79688
rect 132236 79552 132264 79716
rect 132310 79704 132316 79756
rect 132368 79704 132374 79756
rect 132512 79688 132540 79920
rect 132908 79908 132914 79920
rect 132966 79908 132972 79960
rect 133000 79908 133006 79960
rect 133058 79908 133064 79960
rect 132632 79880 132638 79892
rect 132604 79840 132638 79880
rect 132690 79840 132696 79892
rect 133110 79880 133138 79988
rect 133846 79960 133874 79988
rect 134536 79988 135346 80016
rect 133368 79908 133374 79960
rect 133426 79908 133432 79960
rect 133460 79908 133466 79960
rect 133518 79908 133524 79960
rect 133552 79908 133558 79960
rect 133610 79908 133616 79960
rect 133828 79908 133834 79960
rect 133886 79908 133892 79960
rect 134104 79908 134110 79960
rect 134162 79908 134168 79960
rect 134196 79908 134202 79960
rect 134254 79908 134260 79960
rect 132972 79852 133138 79880
rect 132494 79636 132500 79688
rect 132552 79636 132558 79688
rect 132218 79500 132224 79552
rect 132276 79500 132282 79552
rect 132604 79540 132632 79840
rect 132972 79824 133000 79852
rect 133276 79840 133282 79892
rect 133334 79840 133340 79892
rect 132724 79812 132730 79824
rect 132696 79772 132730 79812
rect 132782 79772 132788 79824
rect 132954 79772 132960 79824
rect 133012 79772 133018 79824
rect 132696 79688 132724 79772
rect 133294 79688 133322 79840
rect 133386 79756 133414 79908
rect 133478 79824 133506 79908
rect 133570 79880 133598 79908
rect 133570 79852 133644 79880
rect 133478 79784 133512 79824
rect 133506 79772 133512 79784
rect 133564 79772 133570 79824
rect 133386 79716 133420 79756
rect 133414 79704 133420 79716
rect 133472 79704 133478 79756
rect 132678 79636 132684 79688
rect 132736 79636 132742 79688
rect 133294 79648 133328 79688
rect 133322 79636 133328 79648
rect 133380 79636 133386 79688
rect 132770 79568 132776 79620
rect 132828 79608 132834 79620
rect 133616 79608 133644 79852
rect 133920 79840 133926 79892
rect 133978 79840 133984 79892
rect 132828 79580 133644 79608
rect 132828 79568 132834 79580
rect 133782 79568 133788 79620
rect 133840 79608 133846 79620
rect 133938 79608 133966 79840
rect 134122 79620 134150 79908
rect 133840 79580 133966 79608
rect 133840 79568 133846 79580
rect 134058 79568 134064 79620
rect 134116 79580 134150 79620
rect 134116 79568 134122 79580
rect 134214 79552 134242 79908
rect 134536 79620 134564 79988
rect 135318 79960 135346 79988
rect 136054 79988 136266 80016
rect 136054 79960 136082 79988
rect 135116 79908 135122 79960
rect 135174 79908 135180 79960
rect 135208 79908 135214 79960
rect 135266 79908 135272 79960
rect 135300 79908 135306 79960
rect 135358 79908 135364 79960
rect 135392 79908 135398 79960
rect 135450 79908 135456 79960
rect 136036 79908 136042 79960
rect 136094 79908 136100 79960
rect 136128 79908 136134 79960
rect 136186 79908 136192 79960
rect 134840 79840 134846 79892
rect 134898 79840 134904 79892
rect 134858 79812 134886 79840
rect 134812 79784 134886 79812
rect 134812 79676 134840 79784
rect 134886 79704 134892 79756
rect 134944 79744 134950 79756
rect 135134 79744 135162 79908
rect 134944 79716 135162 79744
rect 134944 79704 134950 79716
rect 135226 79688 135254 79908
rect 135410 79824 135438 79908
rect 135576 79840 135582 79892
rect 135634 79840 135640 79892
rect 135760 79840 135766 79892
rect 135818 79880 135824 79892
rect 135818 79852 135944 79880
rect 135818 79840 135824 79852
rect 135346 79772 135352 79824
rect 135404 79784 135438 79824
rect 135404 79772 135410 79784
rect 134978 79676 134984 79688
rect 134812 79648 134984 79676
rect 134978 79636 134984 79648
rect 135036 79636 135042 79688
rect 135162 79636 135168 79688
rect 135220 79648 135254 79688
rect 135594 79676 135622 79840
rect 135668 79772 135674 79824
rect 135726 79812 135732 79824
rect 135726 79772 135760 79812
rect 135732 79688 135760 79772
rect 135806 79704 135812 79756
rect 135864 79704 135870 79756
rect 135410 79648 135622 79676
rect 135220 79636 135226 79648
rect 134518 79568 134524 79620
rect 134576 79568 134582 79620
rect 135254 79568 135260 79620
rect 135312 79608 135318 79620
rect 135410 79608 135438 79648
rect 135714 79636 135720 79688
rect 135772 79636 135778 79688
rect 135312 79580 135438 79608
rect 135312 79568 135318 79580
rect 135530 79568 135536 79620
rect 135588 79608 135594 79620
rect 135824 79608 135852 79704
rect 135916 79688 135944 79852
rect 135898 79636 135904 79688
rect 135956 79636 135962 79688
rect 135990 79636 135996 79688
rect 136048 79676 136054 79688
rect 136146 79676 136174 79908
rect 136048 79648 136174 79676
rect 136048 79636 136054 79648
rect 135588 79580 135852 79608
rect 135588 79568 135594 79580
rect 136082 79568 136088 79620
rect 136140 79608 136146 79620
rect 136238 79608 136266 79988
rect 137434 79960 137462 80056
rect 137710 79988 138060 80016
rect 136312 79908 136318 79960
rect 136370 79908 136376 79960
rect 136680 79908 136686 79960
rect 136738 79908 136744 79960
rect 136772 79908 136778 79960
rect 136830 79908 136836 79960
rect 137048 79908 137054 79960
rect 137106 79908 137112 79960
rect 137140 79908 137146 79960
rect 137198 79908 137204 79960
rect 137232 79908 137238 79960
rect 137290 79908 137296 79960
rect 137324 79908 137330 79960
rect 137382 79908 137388 79960
rect 137416 79908 137422 79960
rect 137474 79908 137480 79960
rect 137600 79908 137606 79960
rect 137658 79908 137664 79960
rect 136140 79580 136266 79608
rect 136140 79568 136146 79580
rect 133138 79540 133144 79552
rect 132604 79512 133144 79540
rect 133138 79500 133144 79512
rect 133196 79500 133202 79552
rect 134150 79500 134156 79552
rect 134208 79512 134242 79552
rect 134208 79500 134214 79512
rect 135898 79500 135904 79552
rect 135956 79540 135962 79552
rect 136330 79540 136358 79908
rect 136698 79880 136726 79908
rect 135956 79512 136358 79540
rect 136652 79852 136726 79880
rect 136652 79540 136680 79852
rect 136790 79824 136818 79908
rect 136864 79840 136870 79892
rect 136922 79840 136928 79892
rect 136726 79772 136732 79824
rect 136784 79784 136818 79824
rect 136784 79772 136790 79784
rect 136882 79688 136910 79840
rect 137066 79812 137094 79908
rect 137020 79784 137094 79812
rect 136882 79648 136916 79688
rect 136910 79636 136916 79648
rect 136968 79636 136974 79688
rect 136818 79568 136824 79620
rect 136876 79608 136882 79620
rect 137020 79608 137048 79784
rect 137158 79744 137186 79908
rect 137112 79716 137186 79744
rect 137250 79744 137278 79908
rect 137342 79812 137370 79908
rect 137342 79784 137508 79812
rect 137370 79744 137376 79756
rect 137250 79716 137376 79744
rect 137112 79620 137140 79716
rect 137370 79704 137376 79716
rect 137428 79704 137434 79756
rect 136876 79580 137048 79608
rect 136876 79568 136882 79580
rect 137094 79568 137100 79620
rect 137152 79568 137158 79620
rect 137186 79568 137192 79620
rect 137244 79608 137250 79620
rect 137480 79608 137508 79784
rect 137244 79580 137508 79608
rect 137244 79568 137250 79580
rect 137002 79540 137008 79552
rect 136652 79512 137008 79540
rect 135956 79500 135962 79512
rect 137002 79500 137008 79512
rect 137060 79500 137066 79552
rect 137462 79500 137468 79552
rect 137520 79540 137526 79552
rect 137618 79540 137646 79908
rect 137710 79892 137738 79988
rect 137876 79908 137882 79960
rect 137934 79908 137940 79960
rect 137692 79840 137698 79892
rect 137750 79840 137756 79892
rect 137784 79840 137790 79892
rect 137842 79840 137848 79892
rect 137802 79688 137830 79840
rect 137894 79824 137922 79908
rect 137894 79784 137928 79824
rect 137922 79772 137928 79784
rect 137980 79772 137986 79824
rect 137738 79636 137744 79688
rect 137796 79648 137830 79688
rect 137796 79636 137802 79648
rect 137520 79512 137646 79540
rect 137520 79500 137526 79512
rect 131724 79444 131942 79472
rect 131724 79432 131730 79444
rect 135622 79432 135628 79484
rect 135680 79472 135686 79484
rect 136174 79472 136180 79484
rect 135680 79444 136180 79472
rect 135680 79432 135686 79444
rect 136174 79432 136180 79444
rect 136232 79432 136238 79484
rect 128596 79376 129688 79404
rect 128596 79364 128602 79376
rect 129918 79364 129924 79416
rect 129976 79404 129982 79416
rect 135530 79404 135536 79416
rect 129976 79376 135536 79404
rect 129976 79364 129982 79376
rect 135530 79364 135536 79376
rect 135588 79364 135594 79416
rect 136174 79336 136180 79348
rect 128464 79308 136180 79336
rect 136174 79296 136180 79308
rect 136232 79296 136238 79348
rect 138032 79336 138060 79988
rect 138124 79988 138934 80016
rect 138124 79688 138152 79988
rect 138906 79960 138934 79988
rect 139642 79988 139854 80016
rect 138336 79908 138342 79960
rect 138394 79908 138400 79960
rect 138796 79908 138802 79960
rect 138854 79908 138860 79960
rect 138888 79908 138894 79960
rect 138946 79908 138952 79960
rect 138980 79908 138986 79960
rect 139038 79908 139044 79960
rect 139348 79908 139354 79960
rect 139406 79908 139412 79960
rect 139532 79908 139538 79960
rect 139590 79908 139596 79960
rect 138244 79840 138250 79892
rect 138302 79840 138308 79892
rect 138106 79636 138112 79688
rect 138164 79636 138170 79688
rect 138262 79472 138290 79840
rect 138354 79540 138382 79908
rect 138704 79880 138710 79892
rect 138676 79840 138710 79880
rect 138762 79840 138768 79892
rect 138814 79880 138842 79908
rect 138814 79852 138934 79880
rect 138520 79772 138526 79824
rect 138578 79772 138584 79824
rect 138538 79620 138566 79772
rect 138676 79756 138704 79840
rect 138658 79704 138664 79756
rect 138716 79704 138722 79756
rect 138474 79568 138480 79620
rect 138532 79580 138566 79620
rect 138532 79568 138538 79580
rect 138566 79540 138572 79552
rect 138354 79512 138572 79540
rect 138566 79500 138572 79512
rect 138624 79500 138630 79552
rect 138906 79540 138934 79852
rect 138998 79676 139026 79908
rect 139256 79840 139262 79892
rect 139314 79840 139320 79892
rect 139118 79676 139124 79688
rect 138998 79648 139124 79676
rect 139118 79636 139124 79648
rect 139176 79636 139182 79688
rect 139274 79620 139302 79840
rect 139366 79688 139394 79908
rect 139550 79824 139578 79908
rect 139486 79772 139492 79824
rect 139544 79784 139578 79824
rect 139544 79772 139550 79784
rect 139642 79688 139670 79988
rect 139826 79960 139854 79988
rect 139716 79908 139722 79960
rect 139774 79908 139780 79960
rect 139808 79908 139814 79960
rect 139866 79908 139872 79960
rect 140176 79908 140182 79960
rect 140234 79948 140240 79960
rect 140234 79920 140498 79948
rect 140234 79908 140240 79920
rect 139366 79648 139400 79688
rect 139394 79636 139400 79648
rect 139452 79636 139458 79688
rect 139578 79636 139584 79688
rect 139636 79648 139670 79688
rect 139636 79636 139642 79648
rect 139274 79580 139308 79620
rect 139302 79568 139308 79580
rect 139360 79568 139366 79620
rect 139734 79608 139762 79908
rect 140268 79880 140274 79892
rect 140240 79840 140274 79880
rect 140326 79840 140332 79892
rect 140360 79840 140366 79892
rect 140418 79840 140424 79892
rect 140240 79688 140268 79840
rect 140222 79636 140228 79688
rect 140280 79636 140286 79688
rect 140038 79608 140044 79620
rect 139734 79580 140044 79608
rect 140038 79568 140044 79580
rect 140096 79568 140102 79620
rect 140378 79608 140406 79840
rect 140240 79580 140406 79608
rect 139118 79540 139124 79552
rect 138906 79512 139124 79540
rect 139118 79500 139124 79512
rect 139176 79500 139182 79552
rect 138382 79472 138388 79484
rect 138262 79444 138388 79472
rect 138382 79432 138388 79444
rect 138440 79432 138446 79484
rect 140240 79472 140268 79580
rect 140314 79500 140320 79552
rect 140372 79540 140378 79552
rect 140470 79540 140498 79920
rect 140636 79908 140642 79960
rect 140694 79908 140700 79960
rect 141004 79908 141010 79960
rect 141062 79908 141068 79960
rect 141740 79948 141746 79960
rect 141712 79908 141746 79948
rect 141798 79908 141804 79960
rect 141832 79908 141838 79960
rect 141890 79908 141896 79960
rect 141924 79908 141930 79960
rect 141982 79908 141988 79960
rect 142384 79908 142390 79960
rect 142442 79908 142448 79960
rect 140654 79688 140682 79908
rect 140820 79880 140826 79892
rect 140792 79840 140826 79880
rect 140878 79840 140884 79892
rect 140792 79756 140820 79840
rect 141022 79824 141050 79908
rect 141188 79840 141194 79892
rect 141246 79840 141252 79892
rect 141556 79840 141562 79892
rect 141614 79880 141620 79892
rect 141614 79840 141648 79880
rect 140958 79772 140964 79824
rect 141016 79784 141050 79824
rect 141016 79772 141022 79784
rect 140774 79704 140780 79756
rect 140832 79704 140838 79756
rect 140866 79704 140872 79756
rect 140924 79744 140930 79756
rect 141206 79744 141234 79840
rect 140924 79716 141234 79744
rect 140924 79704 140930 79716
rect 140590 79636 140596 79688
rect 140648 79648 140682 79688
rect 140648 79636 140654 79648
rect 140372 79512 140498 79540
rect 140372 79500 140378 79512
rect 141326 79500 141332 79552
rect 141384 79540 141390 79552
rect 141620 79540 141648 79840
rect 141712 79620 141740 79908
rect 141850 79824 141878 79908
rect 141786 79772 141792 79824
rect 141844 79784 141878 79824
rect 141844 79772 141850 79784
rect 141942 79620 141970 79908
rect 141694 79568 141700 79620
rect 141752 79568 141758 79620
rect 141942 79580 141976 79620
rect 141970 79568 141976 79580
rect 142028 79568 142034 79620
rect 142154 79568 142160 79620
rect 142212 79608 142218 79620
rect 142402 79608 142430 79908
rect 142476 79840 142482 79892
rect 142534 79840 142540 79892
rect 142212 79580 142430 79608
rect 142212 79568 142218 79580
rect 142494 79552 142522 79840
rect 142632 79552 142660 80056
rect 143230 79988 143534 80016
rect 143120 79948 143126 79960
rect 143092 79908 143126 79948
rect 143178 79908 143184 79960
rect 142936 79840 142942 79892
rect 142994 79840 143000 79892
rect 141384 79512 141648 79540
rect 141384 79500 141390 79512
rect 142430 79500 142436 79552
rect 142488 79512 142522 79552
rect 142488 79500 142494 79512
rect 142614 79500 142620 79552
rect 142672 79500 142678 79552
rect 142954 79540 142982 79840
rect 143092 79688 143120 79908
rect 143230 79824 143258 79988
rect 143506 79960 143534 79988
rect 143874 79960 143902 80124
rect 147646 80084 147674 80124
rect 147646 80056 151768 80084
rect 143966 79988 144914 80016
rect 143304 79908 143310 79960
rect 143362 79908 143368 79960
rect 143488 79908 143494 79960
rect 143546 79908 143552 79960
rect 143856 79908 143862 79960
rect 143914 79908 143920 79960
rect 143166 79772 143172 79824
rect 143224 79784 143258 79824
rect 143322 79824 143350 79908
rect 143580 79840 143586 79892
rect 143638 79880 143644 79892
rect 143966 79880 143994 79988
rect 144040 79908 144046 79960
rect 144098 79908 144104 79960
rect 144224 79908 144230 79960
rect 144282 79908 144288 79960
rect 144316 79908 144322 79960
rect 144374 79908 144380 79960
rect 144500 79908 144506 79960
rect 144558 79908 144564 79960
rect 144684 79908 144690 79960
rect 144742 79908 144748 79960
rect 144776 79908 144782 79960
rect 144834 79908 144840 79960
rect 143638 79852 143994 79880
rect 143638 79840 143644 79852
rect 143322 79784 143356 79824
rect 143224 79772 143230 79784
rect 143350 79772 143356 79784
rect 143408 79772 143414 79824
rect 143672 79772 143678 79824
rect 143730 79772 143736 79824
rect 143074 79636 143080 79688
rect 143132 79636 143138 79688
rect 143690 79676 143718 79772
rect 143460 79648 143718 79676
rect 143258 79540 143264 79552
rect 142954 79512 143264 79540
rect 143258 79500 143264 79512
rect 143316 79500 143322 79552
rect 143460 79540 143488 79648
rect 143534 79568 143540 79620
rect 143592 79608 143598 79620
rect 144058 79608 144086 79908
rect 144242 79880 144270 79908
rect 143592 79580 144086 79608
rect 144196 79852 144270 79880
rect 143592 79568 143598 79580
rect 143994 79540 144000 79552
rect 143460 79512 144000 79540
rect 143994 79500 144000 79512
rect 144052 79500 144058 79552
rect 144196 79540 144224 79852
rect 144334 79824 144362 79908
rect 144518 79824 144546 79908
rect 144270 79772 144276 79824
rect 144328 79784 144362 79824
rect 144328 79772 144334 79784
rect 144500 79772 144506 79824
rect 144558 79772 144564 79824
rect 144454 79568 144460 79620
rect 144512 79608 144518 79620
rect 144702 79608 144730 79908
rect 144512 79580 144730 79608
rect 144794 79608 144822 79908
rect 144886 79756 144914 79988
rect 144978 79988 148962 80016
rect 144978 79892 145006 79988
rect 145420 79908 145426 79960
rect 145478 79908 145484 79960
rect 145512 79908 145518 79960
rect 145570 79908 145576 79960
rect 145696 79908 145702 79960
rect 145754 79908 145760 79960
rect 145788 79908 145794 79960
rect 145846 79908 145852 79960
rect 146524 79908 146530 79960
rect 146582 79908 146588 79960
rect 146616 79908 146622 79960
rect 146674 79948 146680 79960
rect 146674 79920 146846 79948
rect 146674 79908 146680 79920
rect 144960 79840 144966 79892
rect 145018 79840 145024 79892
rect 145144 79840 145150 79892
rect 145202 79840 145208 79892
rect 145328 79880 145334 79892
rect 145254 79852 145334 79880
rect 144886 79716 144920 79756
rect 144914 79704 144920 79716
rect 144972 79704 144978 79756
rect 145162 79744 145190 79840
rect 145024 79716 145190 79744
rect 145024 79688 145052 79716
rect 145254 79688 145282 79852
rect 145328 79840 145334 79852
rect 145386 79840 145392 79892
rect 145438 79688 145466 79908
rect 145530 79756 145558 79908
rect 145714 79756 145742 79908
rect 145530 79716 145564 79756
rect 145558 79704 145564 79716
rect 145616 79704 145622 79756
rect 145650 79704 145656 79756
rect 145708 79716 145742 79756
rect 145708 79704 145714 79716
rect 145006 79636 145012 79688
rect 145064 79636 145070 79688
rect 145190 79636 145196 79688
rect 145248 79648 145282 79688
rect 145248 79636 145254 79648
rect 145374 79636 145380 79688
rect 145432 79648 145466 79688
rect 145806 79688 145834 79908
rect 145972 79840 145978 79892
rect 146030 79840 146036 79892
rect 145990 79688 146018 79840
rect 146432 79772 146438 79824
rect 146490 79772 146496 79824
rect 145806 79648 145840 79688
rect 145432 79636 145438 79648
rect 145834 79636 145840 79648
rect 145892 79636 145898 79688
rect 145926 79636 145932 79688
rect 145984 79648 146018 79688
rect 146450 79688 146478 79772
rect 146542 79744 146570 79908
rect 146708 79880 146714 79892
rect 146680 79840 146714 79880
rect 146766 79840 146772 79892
rect 146542 79716 146616 79744
rect 146450 79648 146484 79688
rect 145984 79636 145990 79648
rect 146478 79636 146484 79648
rect 146536 79636 146542 79688
rect 146588 79620 146616 79716
rect 146680 79620 146708 79840
rect 146818 79688 146846 79920
rect 146892 79908 146898 79960
rect 146950 79908 146956 79960
rect 147352 79908 147358 79960
rect 147410 79908 147416 79960
rect 146754 79636 146760 79688
rect 146812 79648 146846 79688
rect 146812 79636 146818 79648
rect 146386 79608 146392 79620
rect 144794 79580 146392 79608
rect 144512 79568 144518 79580
rect 146386 79568 146392 79580
rect 146444 79568 146450 79620
rect 146570 79568 146576 79620
rect 146628 79568 146634 79620
rect 146662 79568 146668 79620
rect 146720 79568 146726 79620
rect 146910 79608 146938 79908
rect 147168 79840 147174 79892
rect 147226 79840 147232 79892
rect 147260 79840 147266 79892
rect 147318 79840 147324 79892
rect 147186 79676 147214 79840
rect 147278 79744 147306 79840
rect 147370 79812 147398 79908
rect 147720 79840 147726 79892
rect 147778 79880 147784 79892
rect 147778 79852 148318 79880
rect 147778 79840 147784 79852
rect 147370 79784 147628 79812
rect 147278 79716 147536 79744
rect 147186 79648 147260 79676
rect 147122 79608 147128 79620
rect 146910 79580 147128 79608
rect 147122 79568 147128 79580
rect 147180 79568 147186 79620
rect 146202 79540 146208 79552
rect 144196 79512 146208 79540
rect 146202 79500 146208 79512
rect 146260 79500 146266 79552
rect 147030 79500 147036 79552
rect 147088 79540 147094 79552
rect 147232 79540 147260 79648
rect 147508 79620 147536 79716
rect 147600 79620 147628 79784
rect 147904 79772 147910 79824
rect 147962 79772 147968 79824
rect 147996 79772 148002 79824
rect 148054 79772 148060 79824
rect 148088 79772 148094 79824
rect 148146 79772 148152 79824
rect 147490 79568 147496 79620
rect 147548 79568 147554 79620
rect 147582 79568 147588 79620
rect 147640 79568 147646 79620
rect 147088 79512 147260 79540
rect 147088 79500 147094 79512
rect 147766 79500 147772 79552
rect 147824 79540 147830 79552
rect 147922 79540 147950 79772
rect 148014 79620 148042 79772
rect 148106 79744 148134 79772
rect 148106 79716 148180 79744
rect 148014 79580 148048 79620
rect 148042 79568 148048 79580
rect 148100 79568 148106 79620
rect 147824 79512 147950 79540
rect 147824 79500 147830 79512
rect 143166 79472 143172 79484
rect 140240 79444 143172 79472
rect 143166 79432 143172 79444
rect 143224 79432 143230 79484
rect 147858 79432 147864 79484
rect 147916 79472 147922 79484
rect 148152 79472 148180 79716
rect 148290 79540 148318 79852
rect 148364 79840 148370 79892
rect 148422 79840 148428 79892
rect 148548 79840 148554 79892
rect 148606 79840 148612 79892
rect 148382 79676 148410 79840
rect 148566 79744 148594 79840
rect 148566 79716 148732 79744
rect 148704 79688 148732 79716
rect 148382 79648 148502 79676
rect 148474 79608 148502 79648
rect 148686 79636 148692 79688
rect 148744 79636 148750 79688
rect 148934 79620 148962 79988
rect 149008 79908 149014 79960
rect 149066 79908 149072 79960
rect 150296 79908 150302 79960
rect 150354 79908 150360 79960
rect 150572 79908 150578 79960
rect 150630 79908 150636 79960
rect 150756 79908 150762 79960
rect 150814 79908 150820 79960
rect 150848 79908 150854 79960
rect 150906 79908 150912 79960
rect 150940 79908 150946 79960
rect 150998 79908 151004 79960
rect 151216 79908 151222 79960
rect 151274 79908 151280 79960
rect 151492 79908 151498 79960
rect 151550 79908 151556 79960
rect 149026 79676 149054 79908
rect 149376 79840 149382 79892
rect 149434 79840 149440 79892
rect 149468 79840 149474 79892
rect 149526 79880 149532 79892
rect 149526 79840 149560 79880
rect 149836 79840 149842 79892
rect 149894 79840 149900 79892
rect 149928 79840 149934 79892
rect 149986 79880 149992 79892
rect 149986 79852 150204 79880
rect 149986 79840 149992 79852
rect 149100 79772 149106 79824
rect 149158 79812 149164 79824
rect 149158 79772 149192 79812
rect 149026 79648 149100 79676
rect 149072 79620 149100 79648
rect 149164 79620 149192 79772
rect 149394 79744 149422 79840
rect 149256 79716 149422 79744
rect 148594 79608 148600 79620
rect 148474 79580 148600 79608
rect 148594 79568 148600 79580
rect 148652 79568 148658 79620
rect 148934 79580 148968 79620
rect 148962 79568 148968 79580
rect 149020 79568 149026 79620
rect 149054 79568 149060 79620
rect 149112 79568 149118 79620
rect 149146 79568 149152 79620
rect 149204 79568 149210 79620
rect 148410 79540 148416 79552
rect 148290 79512 148416 79540
rect 148410 79500 148416 79512
rect 148468 79500 148474 79552
rect 149256 79540 149284 79716
rect 149532 79688 149560 79840
rect 149514 79636 149520 79688
rect 149572 79636 149578 79688
rect 149330 79568 149336 79620
rect 149388 79608 149394 79620
rect 149854 79608 149882 79840
rect 150020 79772 150026 79824
rect 150078 79772 150084 79824
rect 150038 79744 150066 79772
rect 149388 79580 149882 79608
rect 149992 79716 150066 79744
rect 149388 79568 149394 79580
rect 149992 79552 150020 79716
rect 150176 79688 150204 79852
rect 150158 79636 150164 79688
rect 150216 79636 150222 79688
rect 150314 79620 150342 79908
rect 150388 79840 150394 79892
rect 150446 79840 150452 79892
rect 150406 79756 150434 79840
rect 150406 79716 150440 79756
rect 150434 79704 150440 79716
rect 150492 79704 150498 79756
rect 150590 79688 150618 79908
rect 150664 79840 150670 79892
rect 150722 79840 150728 79892
rect 150526 79636 150532 79688
rect 150584 79648 150618 79688
rect 150584 79636 150590 79648
rect 150250 79568 150256 79620
rect 150308 79580 150342 79620
rect 150308 79568 150314 79580
rect 149606 79540 149612 79552
rect 149256 79512 149612 79540
rect 149606 79500 149612 79512
rect 149664 79500 149670 79552
rect 149974 79500 149980 79552
rect 150032 79500 150038 79552
rect 150342 79500 150348 79552
rect 150400 79540 150406 79552
rect 150682 79540 150710 79840
rect 150774 79608 150802 79908
rect 150866 79824 150894 79908
rect 150848 79772 150854 79824
rect 150906 79772 150912 79824
rect 150958 79744 150986 79908
rect 150958 79716 151124 79744
rect 150986 79608 150992 79620
rect 150774 79580 150992 79608
rect 150986 79568 150992 79580
rect 151044 79568 151050 79620
rect 150400 79512 150710 79540
rect 150400 79500 150406 79512
rect 150802 79500 150808 79552
rect 150860 79540 150866 79552
rect 151096 79540 151124 79716
rect 151234 79620 151262 79908
rect 151308 79840 151314 79892
rect 151366 79840 151372 79892
rect 151400 79840 151406 79892
rect 151458 79840 151464 79892
rect 151510 79880 151538 79908
rect 151510 79852 151584 79880
rect 151326 79744 151354 79840
rect 151418 79812 151446 79840
rect 151418 79784 151492 79812
rect 151326 79716 151400 79744
rect 151372 79620 151400 79716
rect 151464 79688 151492 79784
rect 151556 79688 151584 79852
rect 151740 79688 151768 80056
rect 151860 79908 151866 79960
rect 151918 79908 151924 79960
rect 151952 79908 151958 79960
rect 152010 79908 152016 79960
rect 152504 79908 152510 79960
rect 152562 79908 152568 79960
rect 152688 79908 152694 79960
rect 152746 79948 152752 79960
rect 152746 79920 152918 79948
rect 152746 79908 152752 79920
rect 151878 79880 151906 79908
rect 151832 79852 151906 79880
rect 151446 79636 151452 79688
rect 151504 79636 151510 79688
rect 151538 79636 151544 79688
rect 151596 79636 151602 79688
rect 151722 79636 151728 79688
rect 151780 79636 151786 79688
rect 151234 79580 151268 79620
rect 151262 79568 151268 79580
rect 151320 79568 151326 79620
rect 151354 79568 151360 79620
rect 151412 79568 151418 79620
rect 150860 79512 151124 79540
rect 151832 79540 151860 79852
rect 151970 79812 151998 79908
rect 152228 79840 152234 79892
rect 152286 79840 152292 79892
rect 151924 79784 151998 79812
rect 151924 79620 151952 79784
rect 152136 79772 152142 79824
rect 152194 79772 152200 79824
rect 152154 79744 152182 79772
rect 152016 79716 152182 79744
rect 152016 79688 152044 79716
rect 151998 79636 152004 79688
rect 152056 79636 152062 79688
rect 152090 79636 152096 79688
rect 152148 79676 152154 79688
rect 152246 79676 152274 79840
rect 152522 79756 152550 79908
rect 152596 79840 152602 79892
rect 152654 79880 152660 79892
rect 152654 79852 152826 79880
rect 152654 79840 152660 79852
rect 152522 79716 152556 79756
rect 152550 79704 152556 79716
rect 152608 79704 152614 79756
rect 152148 79648 152274 79676
rect 152148 79636 152154 79648
rect 151906 79568 151912 79620
rect 151964 79568 151970 79620
rect 152798 79552 152826 79852
rect 152890 79676 152918 79920
rect 152964 79908 152970 79960
rect 153022 79908 153028 79960
rect 153148 79908 153154 79960
rect 153206 79908 153212 79960
rect 153240 79908 153246 79960
rect 153298 79908 153304 79960
rect 153332 79908 153338 79960
rect 153390 79908 153396 79960
rect 153424 79908 153430 79960
rect 153482 79908 153488 79960
rect 152982 79756 153010 79908
rect 153166 79812 153194 79908
rect 153120 79784 153194 79812
rect 153120 79756 153148 79784
rect 153258 79756 153286 79908
rect 152982 79716 153016 79756
rect 153010 79704 153016 79716
rect 153068 79704 153074 79756
rect 153102 79704 153108 79756
rect 153160 79704 153166 79756
rect 153194 79704 153200 79756
rect 153252 79716 153286 79756
rect 153252 79704 153258 79716
rect 153350 79688 153378 79908
rect 152890 79648 152964 79676
rect 152936 79552 152964 79648
rect 153286 79636 153292 79688
rect 153344 79648 153378 79688
rect 153344 79636 153350 79648
rect 152550 79540 152556 79552
rect 151832 79512 152556 79540
rect 150860 79500 150866 79512
rect 152550 79500 152556 79512
rect 152608 79500 152614 79552
rect 152798 79512 152832 79552
rect 152826 79500 152832 79512
rect 152884 79500 152890 79552
rect 152918 79500 152924 79552
rect 152976 79500 152982 79552
rect 153442 79540 153470 79908
rect 153562 79540 153568 79552
rect 153442 79512 153568 79540
rect 153562 79500 153568 79512
rect 153620 79500 153626 79552
rect 147916 79444 148180 79472
rect 153948 79472 153976 80532
rect 154638 79960 154666 80600
rect 161446 80464 173112 80492
rect 161446 80288 161474 80464
rect 173084 80356 173112 80464
rect 173176 80424 173204 80736
rect 174188 80696 174216 80804
rect 178006 80804 580356 80832
rect 178006 80696 178034 80804
rect 580350 80792 580356 80804
rect 580408 80792 580414 80844
rect 178586 80724 178592 80776
rect 178644 80764 178650 80776
rect 580718 80764 580724 80776
rect 178644 80736 580724 80764
rect 178644 80724 178650 80736
rect 580718 80724 580724 80736
rect 580776 80724 580782 80776
rect 580810 80696 580816 80708
rect 174188 80668 174492 80696
rect 174464 80628 174492 80668
rect 174832 80668 178034 80696
rect 180766 80668 580816 80696
rect 174832 80640 174860 80668
rect 174722 80628 174728 80640
rect 174464 80600 174728 80628
rect 174722 80588 174728 80600
rect 174780 80588 174786 80640
rect 174814 80588 174820 80640
rect 174872 80588 174878 80640
rect 174998 80588 175004 80640
rect 175056 80628 175062 80640
rect 180766 80628 180794 80668
rect 580810 80656 580816 80668
rect 580868 80656 580874 80708
rect 175056 80600 180794 80628
rect 175056 80588 175062 80600
rect 176102 80452 176108 80504
rect 176160 80492 176166 80504
rect 181346 80492 181352 80504
rect 176160 80464 181352 80492
rect 176160 80452 176166 80464
rect 181346 80452 181352 80464
rect 181404 80452 181410 80504
rect 174446 80424 174452 80436
rect 173176 80396 174452 80424
rect 174446 80384 174452 80396
rect 174504 80384 174510 80436
rect 174906 80356 174912 80368
rect 173084 80328 174912 80356
rect 174906 80316 174912 80328
rect 174964 80316 174970 80368
rect 174538 80288 174544 80300
rect 158364 80260 161474 80288
rect 163194 80260 174544 80288
rect 154068 79908 154074 79960
rect 154126 79908 154132 79960
rect 154620 79908 154626 79960
rect 154678 79908 154684 79960
rect 156000 79908 156006 79960
rect 156058 79908 156064 79960
rect 156184 79908 156190 79960
rect 156242 79908 156248 79960
rect 156736 79948 156742 79960
rect 156616 79920 156742 79948
rect 154086 79756 154114 79908
rect 154896 79840 154902 79892
rect 154954 79880 154960 79892
rect 154954 79852 155724 79880
rect 154954 79840 154960 79852
rect 154436 79812 154442 79824
rect 154408 79772 154442 79812
rect 154494 79772 154500 79824
rect 155080 79772 155086 79824
rect 155138 79772 155144 79824
rect 155264 79772 155270 79824
rect 155322 79772 155328 79824
rect 155356 79772 155362 79824
rect 155414 79772 155420 79824
rect 155448 79772 155454 79824
rect 155506 79772 155512 79824
rect 154086 79716 154120 79756
rect 154114 79704 154120 79716
rect 154172 79704 154178 79756
rect 154206 79636 154212 79688
rect 154264 79676 154270 79688
rect 154408 79676 154436 79772
rect 155098 79744 155126 79772
rect 155052 79716 155126 79744
rect 155052 79688 155080 79716
rect 154264 79648 154436 79676
rect 154264 79636 154270 79648
rect 155034 79636 155040 79688
rect 155092 79636 155098 79688
rect 155282 79620 155310 79772
rect 155374 79688 155402 79772
rect 155466 79744 155494 79772
rect 155466 79716 155540 79744
rect 155374 79648 155408 79688
rect 155402 79636 155408 79648
rect 155460 79636 155466 79688
rect 155512 79620 155540 79716
rect 154850 79608 154856 79620
rect 154546 79580 154856 79608
rect 154206 79500 154212 79552
rect 154264 79540 154270 79552
rect 154546 79540 154574 79580
rect 154850 79568 154856 79580
rect 154908 79568 154914 79620
rect 155282 79580 155316 79620
rect 155310 79568 155316 79580
rect 155368 79568 155374 79620
rect 155494 79568 155500 79620
rect 155552 79568 155558 79620
rect 155696 79552 155724 79852
rect 155816 79840 155822 79892
rect 155874 79840 155880 79892
rect 155834 79688 155862 79840
rect 156018 79824 156046 79908
rect 156018 79784 156052 79824
rect 156046 79772 156052 79784
rect 156104 79772 156110 79824
rect 156202 79756 156230 79908
rect 156368 79772 156374 79824
rect 156426 79772 156432 79824
rect 156138 79704 156144 79756
rect 156196 79716 156230 79756
rect 156196 79704 156202 79716
rect 155834 79648 155868 79688
rect 155862 79636 155868 79648
rect 155920 79636 155926 79688
rect 156386 79552 156414 79772
rect 154264 79512 154574 79540
rect 154264 79500 154270 79512
rect 155678 79500 155684 79552
rect 155736 79500 155742 79552
rect 156322 79500 156328 79552
rect 156380 79512 156414 79552
rect 156616 79540 156644 79920
rect 156736 79908 156742 79920
rect 156794 79908 156800 79960
rect 156828 79908 156834 79960
rect 156886 79908 156892 79960
rect 157196 79908 157202 79960
rect 157254 79908 157260 79960
rect 157288 79908 157294 79960
rect 157346 79908 157352 79960
rect 157380 79908 157386 79960
rect 157438 79948 157444 79960
rect 157438 79920 157978 79948
rect 157438 79908 157444 79920
rect 156846 79880 156874 79908
rect 156708 79852 156874 79880
rect 156708 79744 156736 79852
rect 157214 79824 157242 79908
rect 157150 79772 157156 79824
rect 157208 79784 157242 79824
rect 157208 79772 157214 79784
rect 156874 79744 156880 79756
rect 156708 79716 156880 79744
rect 156874 79704 156880 79716
rect 156932 79704 156938 79756
rect 157306 79744 157334 79908
rect 157472 79840 157478 79892
rect 157530 79840 157536 79892
rect 157306 79716 157380 79744
rect 156782 79636 156788 79688
rect 156840 79676 156846 79688
rect 157242 79676 157248 79688
rect 156840 79648 157248 79676
rect 156840 79636 156846 79648
rect 157242 79636 157248 79648
rect 157300 79636 157306 79688
rect 156690 79568 156696 79620
rect 156748 79608 156754 79620
rect 157352 79608 157380 79716
rect 157490 79688 157518 79840
rect 157564 79772 157570 79824
rect 157622 79812 157628 79824
rect 157622 79772 157656 79812
rect 157490 79648 157524 79688
rect 157518 79636 157524 79648
rect 157576 79636 157582 79688
rect 157628 79620 157656 79772
rect 157950 79620 157978 79920
rect 158024 79908 158030 79960
rect 158082 79908 158088 79960
rect 158116 79908 158122 79960
rect 158174 79908 158180 79960
rect 158042 79756 158070 79908
rect 158134 79812 158162 79908
rect 158134 79784 158208 79812
rect 158042 79716 158076 79756
rect 158070 79704 158076 79716
rect 158128 79704 158134 79756
rect 156748 79580 157380 79608
rect 156748 79568 156754 79580
rect 157610 79568 157616 79620
rect 157668 79568 157674 79620
rect 157950 79580 157984 79620
rect 157978 79568 157984 79580
rect 158036 79568 158042 79620
rect 156782 79540 156788 79552
rect 156616 79512 156788 79540
rect 156380 79500 156386 79512
rect 156782 79500 156788 79512
rect 156840 79500 156846 79552
rect 157794 79500 157800 79552
rect 157852 79540 157858 79552
rect 158180 79540 158208 79784
rect 158254 79568 158260 79620
rect 158312 79608 158318 79620
rect 158364 79608 158392 80260
rect 163194 80220 163222 80260
rect 174538 80248 174544 80260
rect 174596 80248 174602 80300
rect 176378 80248 176384 80300
rect 176436 80288 176442 80300
rect 200114 80288 200120 80300
rect 176436 80260 200120 80288
rect 176436 80248 176442 80260
rect 200114 80248 200120 80260
rect 200172 80248 200178 80300
rect 159054 80192 163222 80220
rect 159054 79960 159082 80192
rect 174630 80180 174636 80232
rect 174688 80220 174694 80232
rect 231854 80220 231860 80232
rect 174688 80192 231860 80220
rect 174688 80180 174694 80192
rect 231854 80180 231860 80192
rect 231912 80180 231918 80232
rect 174814 80152 174820 80164
rect 167932 80124 170444 80152
rect 162964 80056 165200 80084
rect 158852 79908 158858 79960
rect 158910 79948 158916 79960
rect 158910 79908 158944 79948
rect 159036 79908 159042 79960
rect 159094 79908 159100 79960
rect 159312 79908 159318 79960
rect 159370 79908 159376 79960
rect 160048 79908 160054 79960
rect 160106 79908 160112 79960
rect 160140 79908 160146 79960
rect 160198 79908 160204 79960
rect 160416 79908 160422 79960
rect 160474 79908 160480 79960
rect 160600 79908 160606 79960
rect 160658 79908 160664 79960
rect 160784 79908 160790 79960
rect 160842 79908 160848 79960
rect 160876 79908 160882 79960
rect 160934 79908 160940 79960
rect 161520 79908 161526 79960
rect 161578 79908 161584 79960
rect 161888 79908 161894 79960
rect 161946 79908 161952 79960
rect 162440 79908 162446 79960
rect 162498 79908 162504 79960
rect 162964 79948 162992 80056
rect 165172 80016 165200 80056
rect 167932 80016 167960 80124
rect 163102 79988 165108 80016
rect 165172 79988 167960 80016
rect 163102 79960 163130 79988
rect 162688 79920 162992 79948
rect 158576 79840 158582 79892
rect 158634 79840 158640 79892
rect 158760 79880 158766 79892
rect 158686 79852 158766 79880
rect 158594 79688 158622 79840
rect 158530 79636 158536 79688
rect 158588 79648 158622 79688
rect 158588 79636 158594 79648
rect 158686 79620 158714 79852
rect 158760 79840 158766 79852
rect 158818 79840 158824 79892
rect 158916 79824 158944 79908
rect 159220 79840 159226 79892
rect 159278 79840 159284 79892
rect 159330 79880 159358 79908
rect 159496 79880 159502 79892
rect 159330 79852 159404 79880
rect 158898 79772 158904 79824
rect 158956 79772 158962 79824
rect 158312 79580 158392 79608
rect 158312 79568 158318 79580
rect 158622 79568 158628 79620
rect 158680 79580 158714 79620
rect 159238 79608 159266 79840
rect 159192 79580 159266 79608
rect 158680 79568 158686 79580
rect 157852 79512 158208 79540
rect 157852 79500 157858 79512
rect 153948 79444 155816 79472
rect 147916 79432 147922 79444
rect 139946 79364 139952 79416
rect 140004 79404 140010 79416
rect 152642 79404 152648 79416
rect 140004 79376 152648 79404
rect 140004 79364 140010 79376
rect 152642 79364 152648 79376
rect 152700 79364 152706 79416
rect 153470 79364 153476 79416
rect 153528 79404 153534 79416
rect 153654 79404 153660 79416
rect 153528 79376 153660 79404
rect 153528 79364 153534 79376
rect 153654 79364 153660 79376
rect 153712 79364 153718 79416
rect 155126 79404 155132 79416
rect 153856 79376 155132 79404
rect 144546 79336 144552 79348
rect 138032 79308 144552 79336
rect 144546 79296 144552 79308
rect 144604 79296 144610 79348
rect 153856 79336 153884 79376
rect 155126 79364 155132 79376
rect 155184 79364 155190 79416
rect 144886 79308 153884 79336
rect 155788 79336 155816 79444
rect 158162 79364 158168 79416
rect 158220 79404 158226 79416
rect 158346 79404 158352 79416
rect 158220 79376 158352 79404
rect 158220 79364 158226 79376
rect 158346 79364 158352 79376
rect 158404 79364 158410 79416
rect 159192 79404 159220 79580
rect 159376 79540 159404 79852
rect 159468 79840 159502 79880
rect 159554 79840 159560 79892
rect 159588 79840 159594 79892
rect 159646 79880 159652 79892
rect 159646 79852 159956 79880
rect 159646 79840 159652 79852
rect 159468 79688 159496 79840
rect 159928 79688 159956 79852
rect 159450 79636 159456 79688
rect 159508 79636 159514 79688
rect 159910 79636 159916 79688
rect 159968 79636 159974 79688
rect 160066 79552 160094 79908
rect 160158 79824 160186 79908
rect 160324 79880 160330 79892
rect 160296 79840 160330 79880
rect 160382 79840 160388 79892
rect 160140 79772 160146 79824
rect 160198 79772 160204 79824
rect 159450 79540 159456 79552
rect 159376 79512 159456 79540
rect 159450 79500 159456 79512
rect 159508 79500 159514 79552
rect 160002 79500 160008 79552
rect 160060 79512 160094 79552
rect 160060 79500 160066 79512
rect 159726 79404 159732 79416
rect 159192 79376 159732 79404
rect 159726 79364 159732 79376
rect 159784 79364 159790 79416
rect 160002 79364 160008 79416
rect 160060 79404 160066 79416
rect 160296 79404 160324 79840
rect 160434 79688 160462 79908
rect 160434 79648 160468 79688
rect 160462 79636 160468 79648
rect 160520 79636 160526 79688
rect 160618 79540 160646 79908
rect 160802 79688 160830 79908
rect 160894 79824 160922 79908
rect 161152 79880 161158 79892
rect 161032 79852 161158 79880
rect 160876 79772 160882 79824
rect 160934 79772 160940 79824
rect 160738 79636 160744 79688
rect 160796 79648 160830 79688
rect 160796 79636 160802 79648
rect 161032 79608 161060 79852
rect 161152 79840 161158 79852
rect 161210 79840 161216 79892
rect 161244 79840 161250 79892
rect 161302 79840 161308 79892
rect 161336 79840 161342 79892
rect 161394 79840 161400 79892
rect 161106 79704 161112 79756
rect 161164 79744 161170 79756
rect 161262 79744 161290 79840
rect 161164 79716 161290 79744
rect 161164 79704 161170 79716
rect 161198 79636 161204 79688
rect 161256 79676 161262 79688
rect 161354 79676 161382 79840
rect 161538 79824 161566 79908
rect 161704 79840 161710 79892
rect 161762 79840 161768 79892
rect 161520 79772 161526 79824
rect 161578 79772 161584 79824
rect 161256 79648 161382 79676
rect 161256 79636 161262 79648
rect 161566 79636 161572 79688
rect 161624 79676 161630 79688
rect 161722 79676 161750 79840
rect 161906 79756 161934 79908
rect 161980 79840 161986 79892
rect 162038 79880 162044 79892
rect 162348 79880 162354 79892
rect 162038 79840 162072 79880
rect 161906 79716 161940 79756
rect 161934 79704 161940 79716
rect 161992 79704 161998 79756
rect 162044 79688 162072 79840
rect 162228 79852 162354 79880
rect 161624 79648 161750 79676
rect 161624 79636 161630 79648
rect 162026 79636 162032 79688
rect 162084 79636 162090 79688
rect 162228 79676 162256 79852
rect 162348 79840 162354 79852
rect 162406 79840 162412 79892
rect 162458 79880 162486 79908
rect 162458 79852 162624 79880
rect 162302 79704 162308 79756
rect 162360 79744 162366 79756
rect 162360 79716 162532 79744
rect 162360 79704 162366 79716
rect 162504 79688 162532 79716
rect 162394 79676 162400 79688
rect 162228 79648 162400 79676
rect 162394 79636 162400 79648
rect 162452 79636 162458 79688
rect 162486 79636 162492 79688
rect 162544 79636 162550 79688
rect 161750 79608 161756 79620
rect 161032 79580 161756 79608
rect 161750 79568 161756 79580
rect 161808 79568 161814 79620
rect 162302 79568 162308 79620
rect 162360 79608 162366 79620
rect 162596 79608 162624 79852
rect 162360 79580 162624 79608
rect 162360 79568 162366 79580
rect 160922 79540 160928 79552
rect 160618 79512 160928 79540
rect 160922 79500 160928 79512
rect 160980 79500 160986 79552
rect 162578 79500 162584 79552
rect 162636 79540 162642 79552
rect 162688 79540 162716 79920
rect 163084 79908 163090 79960
rect 163142 79908 163148 79960
rect 164188 79908 164194 79960
rect 164246 79908 164252 79960
rect 164280 79908 164286 79960
rect 164338 79908 164344 79960
rect 164832 79948 164838 79960
rect 164804 79908 164838 79948
rect 164890 79908 164896 79960
rect 164924 79908 164930 79960
rect 164982 79948 164988 79960
rect 164982 79908 165016 79948
rect 162992 79840 162998 79892
rect 163050 79840 163056 79892
rect 163452 79840 163458 79892
rect 163510 79840 163516 79892
rect 163544 79840 163550 79892
rect 163602 79840 163608 79892
rect 163728 79840 163734 79892
rect 163786 79880 163792 79892
rect 163786 79852 163866 79880
rect 163786 79840 163792 79852
rect 163010 79676 163038 79840
rect 162636 79512 162716 79540
rect 162780 79648 163038 79676
rect 162780 79540 162808 79648
rect 162854 79568 162860 79620
rect 162912 79608 162918 79620
rect 163470 79608 163498 79840
rect 163562 79744 163590 79840
rect 163682 79744 163688 79756
rect 163562 79716 163688 79744
rect 163682 79704 163688 79716
rect 163740 79704 163746 79756
rect 162912 79580 163498 79608
rect 162912 79568 162918 79580
rect 162946 79540 162952 79552
rect 162780 79512 162952 79540
rect 162636 79500 162642 79512
rect 162946 79500 162952 79512
rect 163004 79500 163010 79552
rect 163038 79500 163044 79552
rect 163096 79540 163102 79552
rect 163222 79540 163228 79552
rect 163096 79512 163228 79540
rect 163096 79500 163102 79512
rect 163222 79500 163228 79512
rect 163280 79500 163286 79552
rect 160830 79432 160836 79484
rect 160888 79472 160894 79484
rect 160888 79444 162808 79472
rect 160888 79432 160894 79444
rect 160060 79376 160324 79404
rect 160060 79364 160066 79376
rect 160554 79364 160560 79416
rect 160612 79404 160618 79416
rect 161382 79404 161388 79416
rect 160612 79376 161388 79404
rect 160612 79364 160618 79376
rect 161382 79364 161388 79376
rect 161440 79364 161446 79416
rect 161566 79364 161572 79416
rect 161624 79404 161630 79416
rect 162302 79404 162308 79416
rect 161624 79376 162308 79404
rect 161624 79364 161630 79376
rect 162302 79364 162308 79376
rect 162360 79364 162366 79416
rect 162670 79336 162676 79348
rect 155788 79308 162676 79336
rect 120718 79228 120724 79280
rect 120776 79268 120782 79280
rect 144886 79268 144914 79308
rect 162670 79296 162676 79308
rect 162728 79296 162734 79348
rect 162780 79336 162808 79444
rect 163038 79364 163044 79416
rect 163096 79404 163102 79416
rect 163498 79404 163504 79416
rect 163096 79376 163504 79404
rect 163096 79364 163102 79376
rect 163498 79364 163504 79376
rect 163556 79364 163562 79416
rect 163838 79404 163866 79852
rect 164004 79840 164010 79892
rect 164062 79880 164068 79892
rect 164062 79840 164096 79880
rect 164068 79472 164096 79840
rect 164206 79688 164234 79908
rect 164142 79636 164148 79688
rect 164200 79648 164234 79688
rect 164200 79636 164206 79648
rect 164298 79540 164326 79908
rect 164464 79840 164470 79892
rect 164522 79840 164528 79892
rect 164482 79744 164510 79840
rect 164482 79716 164648 79744
rect 164620 79620 164648 79716
rect 164602 79568 164608 79620
rect 164660 79568 164666 79620
rect 164804 79552 164832 79908
rect 164988 79688 165016 79908
rect 164970 79636 164976 79688
rect 165028 79636 165034 79688
rect 164510 79540 164516 79552
rect 164298 79512 164516 79540
rect 164510 79500 164516 79512
rect 164568 79500 164574 79552
rect 164786 79500 164792 79552
rect 164844 79500 164850 79552
rect 165080 79540 165108 79988
rect 165660 79908 165666 79960
rect 165718 79908 165724 79960
rect 165752 79908 165758 79960
rect 165810 79908 165816 79960
rect 166488 79908 166494 79960
rect 166546 79908 166552 79960
rect 166856 79908 166862 79960
rect 166914 79908 166920 79960
rect 168420 79908 168426 79960
rect 168478 79908 168484 79960
rect 168604 79908 168610 79960
rect 168662 79908 168668 79960
rect 168788 79908 168794 79960
rect 168846 79948 168852 79960
rect 168846 79920 169616 79948
rect 168846 79908 168852 79920
rect 165384 79840 165390 79892
rect 165442 79840 165448 79892
rect 165476 79840 165482 79892
rect 165534 79840 165540 79892
rect 165568 79840 165574 79892
rect 165626 79840 165632 79892
rect 165402 79812 165430 79840
rect 165264 79784 165430 79812
rect 165264 79620 165292 79784
rect 165494 79756 165522 79840
rect 165430 79704 165436 79756
rect 165488 79716 165522 79756
rect 165488 79704 165494 79716
rect 165586 79688 165614 79840
rect 165522 79636 165528 79688
rect 165580 79648 165614 79688
rect 165580 79636 165586 79648
rect 165678 79620 165706 79908
rect 165246 79568 165252 79620
rect 165304 79568 165310 79620
rect 165614 79568 165620 79620
rect 165672 79580 165706 79620
rect 165672 79568 165678 79580
rect 165430 79540 165436 79552
rect 165080 79512 165436 79540
rect 165430 79500 165436 79512
rect 165488 79500 165494 79552
rect 165770 79540 165798 79908
rect 166120 79772 166126 79824
rect 166178 79772 166184 79824
rect 166212 79772 166218 79824
rect 166270 79772 166276 79824
rect 166138 79552 166166 79772
rect 166230 79620 166258 79772
rect 166506 79756 166534 79908
rect 166442 79704 166448 79756
rect 166500 79716 166534 79756
rect 166500 79704 166506 79716
rect 166874 79620 166902 79908
rect 167684 79840 167690 79892
rect 167742 79880 167748 79892
rect 167742 79840 167776 79880
rect 167960 79840 167966 79892
rect 168018 79840 168024 79892
rect 167748 79620 167776 79840
rect 167868 79772 167874 79824
rect 167926 79772 167932 79824
rect 167886 79744 167914 79772
rect 167840 79716 167914 79744
rect 167840 79620 167868 79716
rect 167978 79688 168006 79840
rect 168052 79772 168058 79824
rect 168110 79772 168116 79824
rect 167914 79636 167920 79688
rect 167972 79648 168006 79688
rect 168070 79688 168098 79772
rect 168438 79756 168466 79908
rect 168512 79840 168518 79892
rect 168570 79840 168576 79892
rect 168374 79704 168380 79756
rect 168432 79716 168466 79756
rect 168432 79704 168438 79716
rect 168530 79688 168558 79840
rect 168070 79648 168104 79688
rect 167972 79636 167978 79648
rect 168098 79636 168104 79648
rect 168156 79636 168162 79688
rect 168466 79636 168472 79688
rect 168524 79648 168558 79688
rect 168524 79636 168530 79648
rect 168622 79620 168650 79908
rect 169248 79840 169254 79892
rect 169306 79840 169312 79892
rect 169156 79772 169162 79824
rect 169214 79772 169220 79824
rect 166230 79580 166264 79620
rect 166258 79568 166264 79580
rect 166316 79568 166322 79620
rect 166350 79568 166356 79620
rect 166408 79608 166414 79620
rect 166534 79608 166540 79620
rect 166408 79580 166540 79608
rect 166408 79568 166414 79580
rect 166534 79568 166540 79580
rect 166592 79568 166598 79620
rect 166810 79568 166816 79620
rect 166868 79580 166902 79620
rect 166868 79568 166874 79580
rect 167086 79568 167092 79620
rect 167144 79608 167150 79620
rect 167638 79608 167644 79620
rect 167144 79580 167644 79608
rect 167144 79568 167150 79580
rect 167638 79568 167644 79580
rect 167696 79568 167702 79620
rect 167730 79568 167736 79620
rect 167788 79568 167794 79620
rect 167822 79568 167828 79620
rect 167880 79568 167886 79620
rect 168558 79568 168564 79620
rect 168616 79580 168650 79620
rect 169174 79620 169202 79772
rect 169266 79688 169294 79840
rect 169266 79648 169300 79688
rect 169294 79636 169300 79648
rect 169352 79636 169358 79688
rect 169588 79620 169616 79920
rect 169892 79908 169898 79960
rect 169950 79908 169956 79960
rect 169984 79908 169990 79960
rect 170042 79908 170048 79960
rect 170260 79908 170266 79960
rect 170318 79908 170324 79960
rect 169800 79880 169806 79892
rect 169772 79840 169806 79880
rect 169858 79840 169864 79892
rect 169772 79756 169800 79840
rect 169754 79704 169760 79756
rect 169812 79704 169818 79756
rect 169910 79688 169938 79908
rect 170002 79744 170030 79908
rect 170168 79840 170174 79892
rect 170226 79840 170232 79892
rect 170186 79756 170214 79840
rect 170002 79716 170076 79744
rect 169910 79648 169944 79688
rect 169938 79636 169944 79648
rect 169996 79636 170002 79688
rect 169174 79580 169208 79620
rect 168616 79568 168622 79580
rect 169202 79568 169208 79580
rect 169260 79568 169266 79620
rect 169570 79568 169576 79620
rect 169628 79568 169634 79620
rect 169846 79568 169852 79620
rect 169904 79608 169910 79620
rect 170048 79608 170076 79716
rect 170122 79704 170128 79756
rect 170180 79716 170214 79756
rect 170180 79704 170186 79716
rect 170278 79688 170306 79908
rect 170416 79688 170444 80124
rect 172302 80124 174820 80152
rect 172008 79908 172014 79960
rect 172066 79948 172072 79960
rect 172302 79948 172330 80124
rect 174814 80112 174820 80124
rect 174872 80112 174878 80164
rect 174906 80112 174912 80164
rect 174964 80152 174970 80164
rect 252554 80152 252560 80164
rect 174964 80124 252560 80152
rect 174964 80112 174970 80124
rect 252554 80112 252560 80124
rect 252612 80112 252618 80164
rect 175458 80084 175464 80096
rect 172394 80056 175464 80084
rect 172394 79960 172422 80056
rect 175458 80044 175464 80056
rect 175516 80044 175522 80096
rect 175550 80044 175556 80096
rect 175608 80084 175614 80096
rect 430574 80084 430580 80096
rect 175608 80056 430580 80084
rect 175608 80044 175614 80056
rect 430574 80044 430580 80056
rect 430632 80044 430638 80096
rect 178586 80016 178592 80028
rect 172578 79988 178592 80016
rect 172066 79920 172330 79948
rect 172066 79908 172072 79920
rect 172376 79908 172382 79960
rect 172434 79908 172440 79960
rect 170536 79840 170542 79892
rect 170594 79840 170600 79892
rect 172578 79880 172606 79988
rect 178586 79976 178592 79988
rect 178644 79976 178650 80028
rect 172652 79908 172658 79960
rect 172710 79908 172716 79960
rect 172744 79908 172750 79960
rect 172802 79908 172808 79960
rect 172928 79908 172934 79960
rect 172986 79908 172992 79960
rect 173112 79908 173118 79960
rect 173170 79948 173176 79960
rect 173170 79920 173480 79948
rect 173170 79908 173176 79920
rect 171336 79852 172606 79880
rect 170214 79636 170220 79688
rect 170272 79648 170306 79688
rect 170272 79636 170278 79648
rect 170398 79636 170404 79688
rect 170456 79636 170462 79688
rect 169904 79580 170076 79608
rect 169904 79568 169910 79580
rect 170306 79568 170312 79620
rect 170364 79608 170370 79620
rect 170554 79608 170582 79840
rect 170720 79772 170726 79824
rect 170778 79772 170784 79824
rect 171088 79772 171094 79824
rect 171146 79772 171152 79824
rect 170738 79744 170766 79772
rect 170738 79716 170996 79744
rect 170364 79580 170582 79608
rect 170968 79608 170996 79716
rect 171106 79688 171134 79772
rect 171336 79756 171364 79852
rect 171456 79772 171462 79824
rect 171514 79772 171520 79824
rect 171318 79704 171324 79756
rect 171376 79704 171382 79756
rect 171474 79744 171502 79772
rect 171474 79716 172376 79744
rect 171106 79648 171140 79688
rect 171134 79636 171140 79648
rect 171192 79636 171198 79688
rect 171226 79636 171232 79688
rect 171284 79676 171290 79688
rect 172146 79676 172152 79688
rect 171284 79648 172152 79676
rect 171284 79636 171290 79648
rect 172146 79636 172152 79648
rect 172204 79636 172210 79688
rect 172348 79620 172376 79716
rect 172670 79688 172698 79908
rect 172606 79636 172612 79688
rect 172664 79648 172698 79688
rect 172664 79636 172670 79648
rect 171318 79608 171324 79620
rect 170968 79580 171324 79608
rect 170364 79568 170370 79580
rect 171318 79568 171324 79580
rect 171376 79568 171382 79620
rect 172330 79568 172336 79620
rect 172388 79568 172394 79620
rect 172762 79608 172790 79908
rect 172946 79756 172974 79908
rect 173296 79880 173302 79892
rect 173268 79840 173302 79880
rect 173354 79840 173360 79892
rect 173268 79756 173296 79840
rect 172882 79704 172888 79756
rect 172940 79716 172974 79756
rect 172940 79704 172946 79716
rect 173250 79704 173256 79756
rect 173308 79704 173314 79756
rect 173452 79688 173480 79920
rect 173572 79908 173578 79960
rect 173630 79908 173636 79960
rect 173664 79908 173670 79960
rect 173722 79908 173728 79960
rect 173756 79908 173762 79960
rect 173814 79908 173820 79960
rect 173848 79908 173854 79960
rect 173906 79948 173912 79960
rect 174722 79948 174728 79960
rect 173906 79920 174728 79948
rect 173906 79908 173912 79920
rect 174722 79908 174728 79920
rect 174780 79908 174786 79960
rect 173590 79756 173618 79908
rect 173682 79812 173710 79908
rect 173774 79880 173802 79908
rect 173774 79852 173848 79880
rect 173820 79824 173848 79852
rect 174538 79840 174544 79892
rect 174596 79880 174602 79892
rect 175550 79880 175556 79892
rect 174596 79852 175556 79880
rect 174596 79840 174602 79852
rect 175550 79840 175556 79852
rect 175608 79840 175614 79892
rect 173682 79784 173756 79812
rect 173728 79756 173756 79784
rect 173802 79772 173808 79824
rect 173860 79772 173866 79824
rect 179386 79784 183554 79812
rect 173590 79716 173624 79756
rect 173618 79704 173624 79716
rect 173676 79704 173682 79756
rect 173710 79704 173716 79756
rect 173768 79704 173774 79756
rect 173434 79636 173440 79688
rect 173492 79636 173498 79688
rect 179386 79608 179414 79784
rect 172762 79580 179414 79608
rect 183526 79608 183554 79784
rect 201494 79608 201500 79620
rect 183526 79580 201500 79608
rect 201494 79568 201500 79580
rect 201552 79568 201558 79620
rect 165982 79540 165988 79552
rect 165770 79512 165988 79540
rect 165982 79500 165988 79512
rect 166040 79500 166046 79552
rect 166138 79512 166172 79552
rect 166166 79500 166172 79512
rect 166224 79500 166230 79552
rect 171870 79540 171876 79552
rect 166276 79512 171876 79540
rect 164418 79472 164424 79484
rect 164068 79444 164424 79472
rect 164418 79432 164424 79444
rect 164476 79432 164482 79484
rect 166276 79472 166304 79512
rect 171870 79500 171876 79512
rect 171928 79500 171934 79552
rect 172422 79500 172428 79552
rect 172480 79540 172486 79552
rect 180058 79540 180064 79552
rect 172480 79512 180064 79540
rect 172480 79500 172486 79512
rect 180058 79500 180064 79512
rect 180116 79500 180122 79552
rect 166092 79444 166304 79472
rect 164050 79404 164056 79416
rect 163838 79376 164056 79404
rect 164050 79364 164056 79376
rect 164108 79364 164114 79416
rect 166092 79336 166120 79444
rect 167362 79432 167368 79484
rect 167420 79472 167426 79484
rect 171778 79472 171784 79484
rect 167420 79444 171784 79472
rect 167420 79432 167426 79444
rect 171778 79432 171784 79444
rect 171836 79432 171842 79484
rect 172238 79432 172244 79484
rect 172296 79472 172302 79484
rect 527174 79472 527180 79484
rect 172296 79444 527180 79472
rect 172296 79432 172302 79444
rect 527174 79432 527180 79444
rect 527232 79432 527238 79484
rect 171226 79404 171232 79416
rect 162780 79308 166120 79336
rect 166184 79376 171232 79404
rect 157334 79268 157340 79280
rect 120776 79240 126100 79268
rect 120776 79228 120782 79240
rect 121086 79160 121092 79212
rect 121144 79200 121150 79212
rect 126072 79200 126100 79240
rect 131592 79240 144914 79268
rect 147646 79240 157340 79268
rect 121144 79172 126008 79200
rect 126072 79172 126192 79200
rect 121144 79160 121150 79172
rect 125318 79024 125324 79076
rect 125376 79064 125382 79076
rect 125376 79036 125686 79064
rect 125376 79024 125382 79036
rect 125410 78956 125416 79008
rect 125468 78996 125474 79008
rect 125468 78968 125594 78996
rect 125468 78956 125474 78968
rect 125566 78860 125594 78968
rect 125658 78928 125686 79036
rect 125980 78996 126008 79172
rect 126164 79064 126192 79172
rect 131592 79064 131620 79240
rect 147646 79200 147674 79240
rect 157334 79228 157340 79240
rect 157392 79228 157398 79280
rect 157426 79228 157432 79280
rect 157484 79268 157490 79280
rect 157886 79268 157892 79280
rect 157484 79240 157892 79268
rect 157484 79228 157490 79240
rect 157886 79228 157892 79240
rect 157944 79228 157950 79280
rect 157978 79228 157984 79280
rect 158036 79268 158042 79280
rect 166184 79268 166212 79376
rect 171226 79364 171232 79376
rect 171284 79364 171290 79416
rect 173526 79404 173532 79416
rect 171336 79376 173532 79404
rect 166626 79296 166632 79348
rect 166684 79336 166690 79348
rect 171042 79336 171048 79348
rect 166684 79308 171048 79336
rect 166684 79296 166690 79308
rect 171042 79296 171048 79308
rect 171100 79296 171106 79348
rect 171336 79268 171364 79376
rect 173526 79364 173532 79376
rect 173584 79364 173590 79416
rect 176286 79364 176292 79416
rect 176344 79404 176350 79416
rect 580534 79404 580540 79416
rect 176344 79376 580540 79404
rect 176344 79364 176350 79376
rect 580534 79364 580540 79376
rect 580592 79364 580598 79416
rect 171870 79296 171876 79348
rect 171928 79336 171934 79348
rect 173986 79336 173992 79348
rect 171928 79308 173992 79336
rect 171928 79296 171934 79308
rect 173986 79296 173992 79308
rect 174044 79296 174050 79348
rect 176194 79296 176200 79348
rect 176252 79336 176258 79348
rect 580166 79336 580172 79348
rect 176252 79308 580172 79336
rect 176252 79296 176258 79308
rect 580166 79296 580172 79308
rect 580224 79296 580230 79348
rect 158036 79240 166212 79268
rect 166276 79240 171364 79268
rect 158036 79228 158042 79240
rect 161566 79200 161572 79212
rect 126164 79036 131620 79064
rect 135226 79172 147674 79200
rect 152476 79172 161572 79200
rect 135226 78996 135254 79172
rect 136174 79092 136180 79144
rect 136232 79132 136238 79144
rect 152476 79132 152504 79172
rect 161566 79160 161572 79172
rect 161624 79160 161630 79212
rect 165798 79160 165804 79212
rect 165856 79200 165862 79212
rect 166276 79200 166304 79240
rect 172330 79228 172336 79280
rect 172388 79268 172394 79280
rect 183094 79268 183100 79280
rect 172388 79240 183100 79268
rect 172388 79228 172394 79240
rect 183094 79228 183100 79240
rect 183152 79228 183158 79280
rect 165856 79172 166304 79200
rect 165856 79160 165862 79172
rect 167086 79160 167092 79212
rect 167144 79200 167150 79212
rect 167270 79200 167276 79212
rect 167144 79172 167276 79200
rect 167144 79160 167150 79172
rect 167270 79160 167276 79172
rect 167328 79160 167334 79212
rect 168006 79160 168012 79212
rect 168064 79200 168070 79212
rect 168064 79172 169340 79200
rect 168064 79160 168070 79172
rect 136232 79104 152504 79132
rect 136232 79092 136238 79104
rect 152642 79092 152648 79144
rect 152700 79132 152706 79144
rect 154206 79132 154212 79144
rect 152700 79104 154212 79132
rect 152700 79092 152706 79104
rect 154206 79092 154212 79104
rect 154264 79092 154270 79144
rect 155126 79092 155132 79144
rect 155184 79132 155190 79144
rect 167362 79132 167368 79144
rect 155184 79104 167368 79132
rect 155184 79092 155190 79104
rect 167362 79092 167368 79104
rect 167420 79092 167426 79144
rect 168374 79092 168380 79144
rect 168432 79132 168438 79144
rect 168650 79132 168656 79144
rect 168432 79104 168656 79132
rect 168432 79092 168438 79104
rect 168650 79092 168656 79104
rect 168708 79092 168714 79144
rect 169312 79132 169340 79172
rect 171042 79160 171048 79212
rect 171100 79200 171106 79212
rect 174630 79200 174636 79212
rect 171100 79172 174636 79200
rect 171100 79160 171106 79172
rect 174630 79160 174636 79172
rect 174688 79160 174694 79212
rect 174722 79160 174728 79212
rect 174780 79200 174786 79212
rect 183186 79200 183192 79212
rect 174780 79172 183192 79200
rect 174780 79160 174786 79172
rect 183186 79160 183192 79172
rect 183244 79160 183250 79212
rect 249794 79132 249800 79144
rect 169312 79104 249800 79132
rect 249794 79092 249800 79104
rect 249852 79092 249858 79144
rect 135530 79024 135536 79076
rect 135588 79064 135594 79076
rect 139946 79064 139952 79076
rect 135588 79036 139952 79064
rect 135588 79024 135594 79036
rect 139946 79024 139952 79036
rect 140004 79024 140010 79076
rect 145282 79024 145288 79076
rect 145340 79064 145346 79076
rect 152366 79064 152372 79076
rect 145340 79036 152372 79064
rect 145340 79024 145346 79036
rect 152366 79024 152372 79036
rect 152424 79024 152430 79076
rect 153194 79024 153200 79076
rect 153252 79064 153258 79076
rect 160094 79064 160100 79076
rect 153252 79036 160100 79064
rect 153252 79024 153258 79036
rect 160094 79024 160100 79036
rect 160152 79024 160158 79076
rect 161474 79024 161480 79076
rect 161532 79064 161538 79076
rect 165798 79064 165804 79076
rect 161532 79036 165804 79064
rect 161532 79024 161538 79036
rect 165798 79024 165804 79036
rect 165856 79024 165862 79076
rect 167178 79024 167184 79076
rect 167236 79064 167242 79076
rect 167546 79064 167552 79076
rect 167236 79036 167552 79064
rect 167236 79024 167242 79036
rect 167546 79024 167552 79036
rect 167604 79024 167610 79076
rect 168282 79024 168288 79076
rect 168340 79064 168346 79076
rect 195974 79064 195980 79076
rect 168340 79036 195980 79064
rect 168340 79024 168346 79036
rect 195974 79024 195980 79036
rect 196032 79024 196038 79076
rect 125980 78968 135254 78996
rect 151722 78956 151728 79008
rect 151780 78996 151786 79008
rect 152642 78996 152648 79008
rect 151780 78968 152648 78996
rect 151780 78956 151786 78968
rect 152642 78956 152648 78968
rect 152700 78956 152706 79008
rect 153378 78956 153384 79008
rect 153436 78996 153442 79008
rect 153838 78996 153844 79008
rect 153436 78968 153844 78996
rect 153436 78956 153442 78968
rect 153838 78956 153844 78968
rect 153896 78956 153902 79008
rect 154850 78956 154856 79008
rect 154908 78996 154914 79008
rect 154908 78968 159404 78996
rect 154908 78956 154914 78968
rect 132770 78928 132776 78940
rect 125658 78900 132776 78928
rect 132770 78888 132776 78900
rect 132828 78888 132834 78940
rect 148410 78888 148416 78940
rect 148468 78928 148474 78940
rect 157426 78928 157432 78940
rect 148468 78900 157432 78928
rect 148468 78888 148474 78900
rect 157426 78888 157432 78900
rect 157484 78888 157490 78940
rect 157794 78888 157800 78940
rect 157852 78928 157858 78940
rect 159174 78928 159180 78940
rect 157852 78900 159180 78928
rect 157852 78888 157858 78900
rect 159174 78888 159180 78900
rect 159232 78888 159238 78940
rect 159376 78928 159404 78968
rect 160646 78956 160652 79008
rect 160704 78996 160710 79008
rect 161014 78996 161020 79008
rect 160704 78968 161020 78996
rect 160704 78956 160710 78968
rect 161014 78956 161020 78968
rect 161072 78956 161078 79008
rect 162210 78956 162216 79008
rect 162268 78996 162274 79008
rect 267826 78996 267832 79008
rect 162268 78968 267832 78996
rect 162268 78956 162274 78968
rect 267826 78956 267832 78968
rect 267884 78956 267890 79008
rect 167178 78928 167184 78940
rect 159376 78900 167184 78928
rect 167178 78888 167184 78900
rect 167236 78888 167242 78940
rect 167270 78888 167276 78940
rect 167328 78928 167334 78940
rect 213914 78928 213920 78940
rect 167328 78900 213920 78928
rect 167328 78888 167334 78900
rect 213914 78888 213920 78900
rect 213972 78888 213978 78940
rect 131022 78860 131028 78872
rect 125566 78832 131028 78860
rect 131022 78820 131028 78832
rect 131080 78820 131086 78872
rect 137370 78820 137376 78872
rect 137428 78860 137434 78872
rect 137830 78860 137836 78872
rect 137428 78832 137836 78860
rect 137428 78820 137434 78832
rect 137830 78820 137836 78832
rect 137888 78820 137894 78872
rect 150986 78820 150992 78872
rect 151044 78860 151050 78872
rect 151722 78860 151728 78872
rect 151044 78832 151728 78860
rect 151044 78820 151050 78832
rect 151722 78820 151728 78832
rect 151780 78820 151786 78872
rect 157334 78820 157340 78872
rect 157392 78860 157398 78872
rect 160830 78860 160836 78872
rect 157392 78832 160836 78860
rect 157392 78820 157398 78832
rect 160830 78820 160836 78832
rect 160888 78820 160894 78872
rect 161014 78820 161020 78872
rect 161072 78860 161078 78872
rect 172146 78860 172152 78872
rect 161072 78832 172152 78860
rect 161072 78820 161078 78832
rect 172146 78820 172152 78832
rect 172204 78820 172210 78872
rect 172238 78820 172244 78872
rect 172296 78860 172302 78872
rect 174722 78860 174728 78872
rect 172296 78832 174728 78860
rect 172296 78820 172302 78832
rect 174722 78820 174728 78832
rect 174780 78820 174786 78872
rect 176746 78820 176752 78872
rect 176804 78860 176810 78872
rect 266354 78860 266360 78872
rect 176804 78832 266360 78860
rect 176804 78820 176810 78832
rect 266354 78820 266360 78832
rect 266412 78820 266418 78872
rect 129642 78752 129648 78804
rect 129700 78792 129706 78804
rect 130102 78792 130108 78804
rect 129700 78764 130108 78792
rect 129700 78752 129706 78764
rect 130102 78752 130108 78764
rect 130160 78752 130166 78804
rect 132586 78752 132592 78804
rect 132644 78792 132650 78804
rect 133046 78792 133052 78804
rect 132644 78764 133052 78792
rect 132644 78752 132650 78764
rect 133046 78752 133052 78764
rect 133104 78752 133110 78804
rect 140958 78752 140964 78804
rect 141016 78792 141022 78804
rect 141418 78792 141424 78804
rect 141016 78764 141424 78792
rect 141016 78752 141022 78764
rect 141418 78752 141424 78764
rect 141476 78752 141482 78804
rect 148042 78752 148048 78804
rect 148100 78792 148106 78804
rect 148100 78764 154574 78792
rect 148100 78752 148106 78764
rect 127158 78684 127164 78736
rect 127216 78724 127222 78736
rect 127986 78724 127992 78736
rect 127216 78696 127992 78724
rect 127216 78684 127222 78696
rect 127986 78684 127992 78696
rect 128044 78684 128050 78736
rect 128998 78684 129004 78736
rect 129056 78724 129062 78736
rect 129182 78724 129188 78736
rect 129056 78696 129188 78724
rect 129056 78684 129062 78696
rect 129182 78684 129188 78696
rect 129240 78684 129246 78736
rect 132770 78684 132776 78736
rect 132828 78724 132834 78736
rect 133230 78724 133236 78736
rect 132828 78696 133236 78724
rect 132828 78684 132834 78696
rect 133230 78684 133236 78696
rect 133288 78684 133294 78736
rect 152274 78684 152280 78736
rect 152332 78724 152338 78736
rect 152458 78724 152464 78736
rect 152332 78696 152464 78724
rect 152332 78684 152338 78696
rect 152458 78684 152464 78696
rect 152516 78684 152522 78736
rect 154546 78724 154574 78764
rect 158622 78752 158628 78804
rect 158680 78792 158686 78804
rect 158680 78764 159036 78792
rect 158680 78752 158686 78764
rect 159008 78724 159036 78764
rect 159082 78752 159088 78804
rect 159140 78792 159146 78804
rect 159634 78792 159640 78804
rect 159140 78764 159640 78792
rect 159140 78752 159146 78764
rect 159634 78752 159640 78764
rect 159692 78752 159698 78804
rect 160094 78752 160100 78804
rect 160152 78792 160158 78804
rect 171502 78792 171508 78804
rect 160152 78764 171508 78792
rect 160152 78752 160158 78764
rect 171502 78752 171508 78764
rect 171560 78752 171566 78804
rect 171962 78752 171968 78804
rect 172020 78792 172026 78804
rect 172422 78792 172428 78804
rect 172020 78764 172428 78792
rect 172020 78752 172026 78764
rect 172422 78752 172428 78764
rect 172480 78752 172486 78804
rect 172514 78752 172520 78804
rect 172572 78792 172578 78804
rect 397454 78792 397460 78804
rect 172572 78764 397460 78792
rect 172572 78752 172578 78764
rect 397454 78752 397460 78764
rect 397512 78752 397518 78804
rect 426434 78724 426440 78736
rect 154546 78696 158852 78724
rect 159008 78696 426440 78724
rect 125778 78616 125784 78668
rect 125836 78656 125842 78668
rect 129918 78656 129924 78668
rect 125836 78628 129924 78656
rect 125836 78616 125842 78628
rect 129918 78616 129924 78628
rect 129976 78616 129982 78668
rect 132862 78616 132868 78668
rect 132920 78656 132926 78668
rect 133046 78656 133052 78668
rect 132920 78628 133052 78656
rect 132920 78616 132926 78628
rect 133046 78616 133052 78628
rect 133104 78616 133110 78668
rect 144454 78616 144460 78668
rect 144512 78656 144518 78668
rect 144822 78656 144828 78668
rect 144512 78628 144828 78656
rect 144512 78616 144518 78628
rect 144822 78616 144828 78628
rect 144880 78616 144886 78668
rect 147766 78616 147772 78668
rect 147824 78656 147830 78668
rect 148134 78656 148140 78668
rect 147824 78628 148140 78656
rect 147824 78616 147830 78628
rect 148134 78616 148140 78628
rect 148192 78616 148198 78668
rect 150434 78616 150440 78668
rect 150492 78656 150498 78668
rect 154298 78656 154304 78668
rect 150492 78628 154304 78656
rect 150492 78616 150498 78628
rect 154298 78616 154304 78628
rect 154356 78616 154362 78668
rect 158824 78656 158852 78696
rect 426434 78684 426440 78696
rect 426492 78684 426498 78736
rect 162578 78656 162584 78668
rect 158824 78628 162584 78656
rect 162578 78616 162584 78628
rect 162636 78616 162642 78668
rect 162946 78616 162952 78668
rect 163004 78656 163010 78668
rect 163314 78656 163320 78668
rect 163004 78628 163320 78656
rect 163004 78616 163010 78628
rect 163314 78616 163320 78628
rect 163372 78616 163378 78668
rect 166258 78616 166264 78668
rect 166316 78656 166322 78668
rect 168006 78656 168012 78668
rect 166316 78628 168012 78656
rect 166316 78616 166322 78628
rect 168006 78616 168012 78628
rect 168064 78616 168070 78668
rect 168374 78616 168380 78668
rect 168432 78656 168438 78668
rect 173802 78656 173808 78668
rect 168432 78628 173808 78656
rect 168432 78616 168438 78628
rect 173802 78616 173808 78628
rect 173860 78616 173866 78668
rect 122190 78548 122196 78600
rect 122248 78588 122254 78600
rect 128630 78588 128636 78600
rect 122248 78560 128636 78588
rect 122248 78548 122254 78560
rect 128630 78548 128636 78560
rect 128688 78548 128694 78600
rect 141142 78548 141148 78600
rect 141200 78588 141206 78600
rect 141970 78588 141976 78600
rect 141200 78560 141976 78588
rect 141200 78548 141206 78560
rect 141970 78548 141976 78560
rect 142028 78548 142034 78600
rect 146294 78548 146300 78600
rect 146352 78588 146358 78600
rect 162210 78588 162216 78600
rect 146352 78560 162216 78588
rect 146352 78548 146358 78560
rect 162210 78548 162216 78560
rect 162268 78548 162274 78600
rect 166902 78548 166908 78600
rect 166960 78588 166966 78600
rect 171962 78588 171968 78600
rect 166960 78560 171968 78588
rect 166960 78548 166966 78560
rect 171962 78548 171968 78560
rect 172020 78548 172026 78600
rect 172606 78548 172612 78600
rect 172664 78588 172670 78600
rect 176746 78588 176752 78600
rect 172664 78560 176752 78588
rect 172664 78548 172670 78560
rect 176746 78548 176752 78560
rect 176804 78548 176810 78600
rect 125778 78480 125784 78532
rect 125836 78520 125842 78532
rect 127066 78520 127072 78532
rect 125836 78492 127072 78520
rect 125836 78480 125842 78492
rect 127066 78480 127072 78492
rect 127124 78480 127130 78532
rect 146754 78480 146760 78532
rect 146812 78520 146818 78532
rect 146812 78492 154574 78520
rect 146812 78480 146818 78492
rect 154546 78452 154574 78492
rect 155862 78480 155868 78532
rect 155920 78520 155926 78532
rect 156690 78520 156696 78532
rect 155920 78492 156696 78520
rect 155920 78480 155926 78492
rect 156690 78480 156696 78492
rect 156748 78480 156754 78532
rect 157426 78480 157432 78532
rect 157484 78520 157490 78532
rect 161014 78520 161020 78532
rect 157484 78492 161020 78520
rect 157484 78480 157490 78492
rect 161014 78480 161020 78492
rect 161072 78480 161078 78532
rect 167178 78480 167184 78532
rect 167236 78520 167242 78532
rect 170858 78520 170864 78532
rect 167236 78492 170864 78520
rect 167236 78480 167242 78492
rect 170858 78480 170864 78492
rect 170916 78480 170922 78532
rect 171870 78480 171876 78532
rect 171928 78520 171934 78532
rect 255958 78520 255964 78532
rect 171928 78492 255964 78520
rect 171928 78480 171934 78492
rect 255958 78480 255964 78492
rect 256016 78480 256022 78532
rect 160094 78452 160100 78464
rect 154546 78424 160100 78452
rect 160094 78412 160100 78424
rect 160152 78412 160158 78464
rect 160370 78412 160376 78464
rect 160428 78452 160434 78464
rect 160738 78452 160744 78464
rect 160428 78424 160744 78452
rect 160428 78412 160434 78424
rect 160738 78412 160744 78424
rect 160796 78412 160802 78464
rect 162302 78412 162308 78464
rect 162360 78452 162366 78464
rect 315298 78452 315304 78464
rect 162360 78424 315304 78452
rect 162360 78412 162366 78424
rect 315298 78412 315304 78424
rect 315356 78412 315362 78464
rect 126974 78344 126980 78396
rect 127032 78384 127038 78396
rect 128354 78384 128360 78396
rect 127032 78356 128360 78384
rect 127032 78344 127038 78356
rect 128354 78344 128360 78356
rect 128412 78344 128418 78396
rect 150342 78344 150348 78396
rect 150400 78384 150406 78396
rect 150710 78384 150716 78396
rect 150400 78356 150716 78384
rect 150400 78344 150406 78356
rect 150710 78344 150716 78356
rect 150768 78344 150774 78396
rect 162762 78344 162768 78396
rect 162820 78384 162826 78396
rect 436738 78384 436744 78396
rect 162820 78356 436744 78384
rect 162820 78344 162826 78356
rect 436738 78344 436744 78356
rect 436796 78344 436802 78396
rect 120718 78276 120724 78328
rect 120776 78316 120782 78328
rect 128262 78316 128268 78328
rect 120776 78288 128268 78316
rect 120776 78276 120782 78288
rect 128262 78276 128268 78288
rect 128320 78276 128326 78328
rect 148962 78276 148968 78328
rect 149020 78316 149026 78328
rect 166258 78316 166264 78328
rect 149020 78288 166264 78316
rect 149020 78276 149026 78288
rect 166258 78276 166264 78288
rect 166316 78276 166322 78328
rect 171870 78316 171876 78328
rect 166966 78288 171876 78316
rect 116578 78208 116584 78260
rect 116636 78248 116642 78260
rect 128814 78248 128820 78260
rect 116636 78220 128820 78248
rect 116636 78208 116642 78220
rect 128814 78208 128820 78220
rect 128872 78208 128878 78260
rect 142430 78208 142436 78260
rect 142488 78248 142494 78260
rect 142706 78248 142712 78260
rect 142488 78220 142712 78248
rect 142488 78208 142494 78220
rect 142706 78208 142712 78220
rect 142764 78208 142770 78260
rect 145006 78208 145012 78260
rect 145064 78248 145070 78260
rect 145742 78248 145748 78260
rect 145064 78220 145748 78248
rect 145064 78208 145070 78220
rect 145742 78208 145748 78220
rect 145800 78208 145806 78260
rect 155402 78208 155408 78260
rect 155460 78248 155466 78260
rect 159634 78248 159640 78260
rect 155460 78220 159640 78248
rect 155460 78208 155466 78220
rect 159634 78208 159640 78220
rect 159692 78208 159698 78260
rect 161750 78208 161756 78260
rect 161808 78248 161814 78260
rect 166966 78248 166994 78288
rect 171870 78276 171876 78288
rect 171928 78276 171934 78328
rect 172054 78276 172060 78328
rect 172112 78316 172118 78328
rect 178770 78316 178776 78328
rect 172112 78288 178776 78316
rect 172112 78276 172118 78288
rect 178770 78276 178776 78288
rect 178828 78276 178834 78328
rect 161808 78220 166994 78248
rect 161808 78208 161814 78220
rect 167362 78208 167368 78260
rect 167420 78248 167426 78260
rect 167546 78248 167552 78260
rect 167420 78220 167552 78248
rect 167420 78208 167426 78220
rect 167546 78208 167552 78220
rect 167604 78208 167610 78260
rect 169018 78208 169024 78260
rect 169076 78248 169082 78260
rect 169202 78248 169208 78260
rect 169076 78220 169208 78248
rect 169076 78208 169082 78220
rect 169202 78208 169208 78220
rect 169260 78208 169266 78260
rect 483014 78248 483020 78260
rect 171796 78220 483020 78248
rect 113818 78140 113824 78192
rect 113876 78180 113882 78192
rect 126790 78180 126796 78192
rect 113876 78152 126796 78180
rect 113876 78140 113882 78152
rect 126790 78140 126796 78152
rect 126848 78140 126854 78192
rect 139394 78140 139400 78192
rect 139452 78180 139458 78192
rect 140130 78180 140136 78192
rect 139452 78152 140136 78180
rect 139452 78140 139458 78152
rect 140130 78140 140136 78152
rect 140188 78140 140194 78192
rect 142062 78140 142068 78192
rect 142120 78180 142126 78192
rect 142120 78152 151676 78180
rect 142120 78140 142126 78152
rect 128262 78072 128268 78124
rect 128320 78112 128326 78124
rect 150618 78112 150624 78124
rect 128320 78084 150624 78112
rect 128320 78072 128326 78084
rect 150618 78072 150624 78084
rect 150676 78072 150682 78124
rect 151648 78056 151676 78152
rect 152366 78140 152372 78192
rect 152424 78180 152430 78192
rect 158254 78180 158260 78192
rect 152424 78152 158260 78180
rect 152424 78140 152430 78152
rect 158254 78140 158260 78152
rect 158312 78140 158318 78192
rect 158714 78140 158720 78192
rect 158772 78180 158778 78192
rect 162302 78180 162308 78192
rect 158772 78152 162308 78180
rect 158772 78140 158778 78152
rect 162302 78140 162308 78152
rect 162360 78140 162366 78192
rect 163130 78140 163136 78192
rect 163188 78180 163194 78192
rect 171796 78180 171824 78220
rect 483014 78208 483020 78220
rect 483072 78208 483078 78260
rect 498194 78180 498200 78192
rect 163188 78152 171824 78180
rect 171888 78152 498200 78180
rect 163188 78140 163194 78152
rect 153378 78072 153384 78124
rect 153436 78112 153442 78124
rect 154114 78112 154120 78124
rect 153436 78084 154120 78112
rect 153436 78072 153442 78084
rect 154114 78072 154120 78084
rect 154172 78072 154178 78124
rect 155494 78072 155500 78124
rect 155552 78112 155558 78124
rect 155862 78112 155868 78124
rect 155552 78084 155868 78112
rect 155552 78072 155558 78084
rect 155862 78072 155868 78084
rect 155920 78072 155926 78124
rect 156138 78072 156144 78124
rect 156196 78112 156202 78124
rect 156414 78112 156420 78124
rect 156196 78084 156420 78112
rect 156196 78072 156202 78084
rect 156414 78072 156420 78084
rect 156472 78072 156478 78124
rect 160094 78072 160100 78124
rect 160152 78112 160158 78124
rect 161290 78112 161296 78124
rect 160152 78084 161296 78112
rect 160152 78072 160158 78084
rect 161290 78072 161296 78084
rect 161348 78072 161354 78124
rect 163222 78072 163228 78124
rect 163280 78112 163286 78124
rect 171778 78112 171784 78124
rect 163280 78084 171784 78112
rect 163280 78072 163286 78084
rect 171778 78072 171784 78084
rect 171836 78072 171842 78124
rect 93118 78004 93124 78056
rect 93176 78044 93182 78056
rect 127434 78044 127440 78056
rect 93176 78016 127440 78044
rect 93176 78004 93182 78016
rect 127434 78004 127440 78016
rect 127492 78004 127498 78056
rect 140498 78004 140504 78056
rect 140556 78044 140562 78056
rect 146294 78044 146300 78056
rect 140556 78016 146300 78044
rect 140556 78004 140562 78016
rect 146294 78004 146300 78016
rect 146352 78004 146358 78056
rect 150986 78004 150992 78056
rect 151044 78044 151050 78056
rect 151170 78044 151176 78056
rect 151044 78016 151176 78044
rect 151044 78004 151050 78016
rect 151170 78004 151176 78016
rect 151228 78004 151234 78056
rect 151630 78004 151636 78056
rect 151688 78004 151694 78056
rect 154482 78004 154488 78056
rect 154540 78044 154546 78056
rect 158622 78044 158628 78056
rect 154540 78016 158628 78044
rect 154540 78004 154546 78016
rect 158622 78004 158628 78016
rect 158680 78004 158686 78056
rect 159174 78004 159180 78056
rect 159232 78044 159238 78056
rect 159232 78016 164234 78044
rect 159232 78004 159238 78016
rect 10318 77936 10324 77988
rect 10376 77976 10382 77988
rect 125962 77976 125968 77988
rect 10376 77948 125968 77976
rect 10376 77936 10382 77948
rect 125962 77936 125968 77948
rect 126020 77936 126026 77988
rect 126790 77936 126796 77988
rect 126848 77976 126854 77988
rect 128538 77976 128544 77988
rect 126848 77948 128544 77976
rect 126848 77936 126854 77948
rect 128538 77936 128544 77948
rect 128596 77936 128602 77988
rect 131758 77936 131764 77988
rect 131816 77976 131822 77988
rect 132218 77976 132224 77988
rect 131816 77948 132224 77976
rect 131816 77936 131822 77948
rect 132218 77936 132224 77948
rect 132276 77936 132282 77988
rect 133230 77936 133236 77988
rect 133288 77976 133294 77988
rect 133414 77976 133420 77988
rect 133288 77948 133420 77976
rect 133288 77936 133294 77948
rect 133414 77936 133420 77948
rect 133472 77936 133478 77988
rect 141602 77936 141608 77988
rect 141660 77976 141666 77988
rect 141786 77976 141792 77988
rect 141660 77948 141792 77976
rect 141660 77936 141666 77948
rect 141786 77936 141792 77948
rect 141844 77936 141850 77988
rect 142246 77936 142252 77988
rect 142304 77976 142310 77988
rect 152366 77976 152372 77988
rect 142304 77948 152372 77976
rect 142304 77936 142310 77948
rect 152366 77936 152372 77948
rect 152424 77936 152430 77988
rect 152642 77936 152648 77988
rect 152700 77976 152706 77988
rect 152700 77948 159818 77976
rect 152700 77936 152706 77948
rect 154114 77868 154120 77920
rect 154172 77908 154178 77920
rect 155494 77908 155500 77920
rect 154172 77880 155500 77908
rect 154172 77868 154178 77880
rect 155494 77868 155500 77880
rect 155552 77868 155558 77920
rect 157610 77868 157616 77920
rect 157668 77908 157674 77920
rect 159790 77908 159818 77948
rect 161566 77936 161572 77988
rect 161624 77976 161630 77988
rect 162118 77976 162124 77988
rect 161624 77948 162124 77976
rect 161624 77936 161630 77948
rect 162118 77936 162124 77948
rect 162176 77936 162182 77988
rect 162210 77908 162216 77920
rect 157668 77880 158392 77908
rect 159790 77880 162216 77908
rect 157668 77868 157674 77880
rect 145006 77800 145012 77852
rect 145064 77840 145070 77852
rect 145374 77840 145380 77852
rect 145064 77812 145380 77840
rect 145064 77800 145070 77812
rect 145374 77800 145380 77812
rect 145432 77800 145438 77852
rect 154666 77800 154672 77852
rect 154724 77840 154730 77852
rect 158254 77840 158260 77852
rect 154724 77812 158260 77840
rect 154724 77800 154730 77812
rect 158254 77800 158260 77812
rect 158312 77800 158318 77852
rect 158364 77840 158392 77880
rect 162210 77868 162216 77880
rect 162268 77868 162274 77920
rect 164206 77908 164234 78016
rect 164510 78004 164516 78056
rect 164568 78044 164574 78056
rect 171888 78044 171916 78152
rect 498194 78140 498200 78152
rect 498252 78140 498258 78192
rect 171962 78072 171968 78124
rect 172020 78112 172026 78124
rect 532694 78112 532700 78124
rect 172020 78084 532700 78112
rect 172020 78072 172026 78084
rect 532694 78072 532700 78084
rect 532752 78072 532758 78124
rect 574738 78044 574744 78056
rect 164568 78016 171916 78044
rect 172532 78016 574744 78044
rect 164568 78004 164574 78016
rect 165614 77936 165620 77988
rect 165672 77976 165678 77988
rect 170582 77976 170588 77988
rect 165672 77948 170588 77976
rect 165672 77936 165678 77948
rect 170582 77936 170588 77948
rect 170640 77936 170646 77988
rect 170674 77936 170680 77988
rect 170732 77976 170738 77988
rect 172532 77976 172560 78016
rect 574738 78004 574744 78016
rect 574796 78004 574802 78056
rect 581086 77976 581092 77988
rect 170732 77948 172560 77976
rect 172624 77948 581092 77976
rect 170732 77936 170738 77948
rect 164206 77880 169570 77908
rect 158364 77812 169340 77840
rect 143166 77732 143172 77784
rect 143224 77772 143230 77784
rect 148410 77772 148416 77784
rect 143224 77744 148416 77772
rect 143224 77732 143230 77744
rect 148410 77732 148416 77744
rect 148468 77732 148474 77784
rect 151446 77732 151452 77784
rect 151504 77772 151510 77784
rect 153838 77772 153844 77784
rect 151504 77744 153844 77772
rect 151504 77732 151510 77744
rect 153838 77732 153844 77744
rect 153896 77732 153902 77784
rect 159174 77732 159180 77784
rect 159232 77772 159238 77784
rect 168282 77772 168288 77784
rect 159232 77744 168288 77772
rect 159232 77732 159238 77744
rect 168282 77732 168288 77744
rect 168340 77732 168346 77784
rect 123478 77664 123484 77716
rect 123536 77704 123542 77716
rect 134794 77704 134800 77716
rect 123536 77676 134800 77704
rect 123536 77664 123542 77676
rect 134794 77664 134800 77676
rect 134852 77664 134858 77716
rect 155954 77664 155960 77716
rect 156012 77704 156018 77716
rect 162118 77704 162124 77716
rect 156012 77676 162124 77704
rect 156012 77664 156018 77676
rect 162118 77664 162124 77676
rect 162176 77664 162182 77716
rect 162302 77664 162308 77716
rect 162360 77704 162366 77716
rect 167178 77704 167184 77716
rect 162360 77676 167184 77704
rect 162360 77664 162366 77676
rect 167178 77664 167184 77676
rect 167236 77664 167242 77716
rect 168466 77664 168472 77716
rect 168524 77704 168530 77716
rect 168742 77704 168748 77716
rect 168524 77676 168748 77704
rect 168524 77664 168530 77676
rect 168742 77664 168748 77676
rect 168800 77664 168806 77716
rect 169312 77704 169340 77812
rect 169542 77772 169570 77880
rect 171318 77868 171324 77920
rect 171376 77908 171382 77920
rect 172624 77908 172652 77948
rect 581086 77936 581092 77948
rect 581144 77936 581150 77988
rect 171376 77880 172652 77908
rect 171376 77868 171382 77880
rect 172698 77868 172704 77920
rect 172756 77908 172762 77920
rect 331214 77908 331220 77920
rect 172756 77880 331220 77908
rect 172756 77868 172762 77880
rect 331214 77868 331220 77880
rect 331272 77868 331278 77920
rect 171594 77800 171600 77852
rect 171652 77840 171658 77852
rect 176286 77840 176292 77852
rect 171652 77812 176292 77840
rect 171652 77800 171658 77812
rect 176286 77800 176292 77812
rect 176344 77800 176350 77852
rect 172146 77772 172152 77784
rect 169542 77744 172152 77772
rect 172146 77732 172152 77744
rect 172204 77732 172210 77784
rect 171594 77704 171600 77716
rect 169312 77676 171600 77704
rect 171594 77664 171600 77676
rect 171652 77664 171658 77716
rect 176194 77664 176200 77716
rect 176252 77704 176258 77716
rect 182910 77704 182916 77716
rect 176252 77676 182916 77704
rect 176252 77664 176258 77676
rect 182910 77664 182916 77676
rect 182968 77664 182974 77716
rect 144914 77596 144920 77648
rect 144972 77636 144978 77648
rect 145834 77636 145840 77648
rect 144972 77608 145840 77636
rect 144972 77596 144978 77608
rect 145834 77596 145840 77608
rect 145892 77596 145898 77648
rect 160922 77596 160928 77648
rect 160980 77636 160986 77648
rect 242158 77636 242164 77648
rect 160980 77608 242164 77636
rect 160980 77596 160986 77608
rect 242158 77596 242164 77608
rect 242216 77596 242222 77648
rect 139670 77528 139676 77580
rect 139728 77568 139734 77580
rect 172054 77568 172060 77580
rect 139728 77540 160692 77568
rect 139728 77528 139734 77540
rect 122098 77460 122104 77512
rect 122156 77500 122162 77512
rect 127342 77500 127348 77512
rect 122156 77472 127348 77500
rect 122156 77460 122162 77472
rect 127342 77460 127348 77472
rect 127400 77460 127406 77512
rect 128814 77460 128820 77512
rect 128872 77500 128878 77512
rect 129826 77500 129832 77512
rect 128872 77472 129832 77500
rect 128872 77460 128878 77472
rect 129826 77460 129832 77472
rect 129884 77460 129890 77512
rect 140774 77460 140780 77512
rect 140832 77500 140838 77512
rect 159174 77500 159180 77512
rect 140832 77472 159180 77500
rect 140832 77460 140838 77472
rect 159174 77460 159180 77472
rect 159232 77460 159238 77512
rect 160664 77500 160692 77540
rect 164206 77540 172060 77568
rect 164206 77500 164234 77540
rect 172054 77528 172060 77540
rect 172112 77528 172118 77580
rect 160664 77472 164234 77500
rect 165614 77460 165620 77512
rect 165672 77500 165678 77512
rect 166166 77500 166172 77512
rect 165672 77472 166172 77500
rect 165672 77460 165678 77472
rect 166166 77460 166172 77472
rect 166224 77460 166230 77512
rect 166258 77460 166264 77512
rect 166316 77500 166322 77512
rect 166442 77500 166448 77512
rect 166316 77472 166448 77500
rect 166316 77460 166322 77472
rect 166442 77460 166448 77472
rect 166500 77460 166506 77512
rect 167178 77460 167184 77512
rect 167236 77500 167242 77512
rect 167730 77500 167736 77512
rect 167236 77472 167736 77500
rect 167236 77460 167242 77472
rect 167730 77460 167736 77472
rect 167788 77460 167794 77512
rect 169662 77460 169668 77512
rect 169720 77500 169726 77512
rect 170214 77500 170220 77512
rect 169720 77472 170220 77500
rect 169720 77460 169726 77472
rect 170214 77460 170220 77472
rect 170272 77460 170278 77512
rect 170398 77460 170404 77512
rect 170456 77500 170462 77512
rect 172330 77500 172336 77512
rect 170456 77472 172336 77500
rect 170456 77460 170462 77472
rect 172330 77460 172336 77472
rect 172388 77460 172394 77512
rect 132862 77392 132868 77444
rect 132920 77432 132926 77444
rect 133690 77432 133696 77444
rect 132920 77404 133696 77432
rect 132920 77392 132926 77404
rect 133690 77392 133696 77404
rect 133748 77392 133754 77444
rect 141970 77392 141976 77444
rect 142028 77432 142034 77444
rect 176378 77432 176384 77444
rect 142028 77404 176384 77432
rect 142028 77392 142034 77404
rect 176378 77392 176384 77404
rect 176436 77392 176442 77444
rect 152366 77324 152372 77376
rect 152424 77364 152430 77376
rect 167270 77364 167276 77376
rect 152424 77336 167276 77364
rect 152424 77324 152430 77336
rect 167270 77324 167276 77336
rect 167328 77324 167334 77376
rect 168558 77324 168564 77376
rect 168616 77364 168622 77376
rect 168834 77364 168840 77376
rect 168616 77336 168840 77364
rect 168616 77324 168622 77336
rect 168834 77324 168840 77336
rect 168892 77324 168898 77376
rect 168926 77324 168932 77376
rect 168984 77364 168990 77376
rect 169110 77364 169116 77376
rect 168984 77336 169116 77364
rect 168984 77324 168990 77336
rect 169110 77324 169116 77336
rect 169168 77324 169174 77376
rect 125042 77256 125048 77308
rect 125100 77296 125106 77308
rect 126698 77296 126704 77308
rect 125100 77268 126704 77296
rect 125100 77256 125106 77268
rect 126698 77256 126704 77268
rect 126756 77256 126762 77308
rect 144822 77256 144828 77308
rect 144880 77296 144886 77308
rect 166626 77296 166632 77308
rect 144880 77268 166632 77296
rect 144880 77256 144886 77268
rect 166626 77256 166632 77268
rect 166684 77256 166690 77308
rect 171778 77256 171784 77308
rect 171836 77296 171842 77308
rect 480254 77296 480260 77308
rect 171836 77268 480260 77296
rect 171836 77256 171842 77268
rect 480254 77256 480260 77268
rect 480312 77256 480318 77308
rect 124858 77188 124864 77240
rect 124916 77228 124922 77240
rect 131206 77228 131212 77240
rect 124916 77200 131212 77228
rect 124916 77188 124922 77200
rect 131206 77188 131212 77200
rect 131264 77188 131270 77240
rect 137002 77188 137008 77240
rect 137060 77228 137066 77240
rect 138934 77228 138940 77240
rect 137060 77200 138940 77228
rect 137060 77188 137066 77200
rect 138934 77188 138940 77200
rect 138992 77188 138998 77240
rect 149330 77188 149336 77240
rect 149388 77228 149394 77240
rect 150066 77228 150072 77240
rect 149388 77200 150072 77228
rect 149388 77188 149394 77200
rect 150066 77188 150072 77200
rect 150124 77188 150130 77240
rect 152366 77188 152372 77240
rect 152424 77228 152430 77240
rect 226334 77228 226340 77240
rect 152424 77200 226340 77228
rect 152424 77188 152430 77200
rect 226334 77188 226340 77200
rect 226392 77188 226398 77240
rect 130286 77120 130292 77172
rect 130344 77160 130350 77172
rect 130562 77160 130568 77172
rect 130344 77132 130568 77160
rect 130344 77120 130350 77132
rect 130562 77120 130568 77132
rect 130620 77120 130626 77172
rect 146202 77120 146208 77172
rect 146260 77160 146266 77172
rect 240134 77160 240140 77172
rect 146260 77132 240140 77160
rect 146260 77120 146266 77132
rect 240134 77120 240140 77132
rect 240192 77120 240198 77172
rect 139302 77052 139308 77104
rect 139360 77092 139366 77104
rect 140498 77092 140504 77104
rect 139360 77064 140504 77092
rect 139360 77052 139366 77064
rect 140498 77052 140504 77064
rect 140556 77052 140562 77104
rect 147306 77052 147312 77104
rect 147364 77092 147370 77104
rect 260834 77092 260840 77104
rect 147364 77064 260840 77092
rect 147364 77052 147370 77064
rect 260834 77052 260840 77064
rect 260892 77052 260898 77104
rect 122834 76984 122840 77036
rect 122892 77024 122898 77036
rect 134886 77024 134892 77036
rect 122892 76996 134892 77024
rect 122892 76984 122898 76996
rect 134886 76984 134892 76996
rect 134944 76984 134950 77036
rect 147950 76984 147956 77036
rect 148008 77024 148014 77036
rect 296714 77024 296720 77036
rect 148008 76996 296720 77024
rect 148008 76984 148014 76996
rect 296714 76984 296720 76996
rect 296772 76984 296778 77036
rect 156046 76916 156052 76968
rect 156104 76956 156110 76968
rect 331122 76956 331128 76968
rect 156104 76928 331128 76956
rect 156104 76916 156110 76928
rect 331122 76916 331128 76928
rect 331180 76916 331186 76968
rect 118694 76848 118700 76900
rect 118752 76888 118758 76900
rect 134978 76888 134984 76900
rect 118752 76860 134984 76888
rect 118752 76848 118758 76860
rect 134978 76848 134984 76860
rect 135036 76848 135042 76900
rect 143074 76848 143080 76900
rect 143132 76888 143138 76900
rect 152366 76888 152372 76900
rect 143132 76860 152372 76888
rect 143132 76848 143138 76860
rect 152366 76848 152372 76860
rect 152424 76848 152430 76900
rect 157426 76848 157432 76900
rect 157484 76888 157490 76900
rect 158346 76888 158352 76900
rect 157484 76860 158352 76888
rect 157484 76848 157490 76860
rect 158346 76848 158352 76860
rect 158404 76848 158410 76900
rect 346394 76888 346400 76900
rect 166966 76860 346400 76888
rect 102134 76780 102140 76832
rect 102192 76820 102198 76832
rect 133506 76820 133512 76832
rect 102192 76792 133512 76820
rect 102192 76780 102198 76792
rect 133506 76780 133512 76792
rect 133564 76780 133570 76832
rect 70394 76712 70400 76764
rect 70452 76752 70458 76764
rect 125410 76752 125416 76764
rect 70452 76724 125416 76752
rect 70452 76712 70458 76724
rect 125410 76712 125416 76724
rect 125468 76712 125474 76764
rect 155034 76712 155040 76764
rect 155092 76752 155098 76764
rect 166966 76752 166994 76860
rect 346394 76848 346400 76860
rect 346452 76848 346458 76900
rect 167270 76780 167276 76832
rect 167328 76820 167334 76832
rect 167914 76820 167920 76832
rect 167328 76792 167920 76820
rect 167328 76780 167334 76792
rect 167914 76780 167920 76792
rect 167972 76780 167978 76832
rect 168834 76780 168840 76832
rect 168892 76820 168898 76832
rect 169386 76820 169392 76832
rect 168892 76792 169392 76820
rect 168892 76780 168898 76792
rect 169386 76780 169392 76792
rect 169444 76780 169450 76832
rect 173986 76780 173992 76832
rect 174044 76820 174050 76832
rect 174354 76820 174360 76832
rect 174044 76792 174360 76820
rect 174044 76780 174050 76792
rect 174354 76780 174360 76792
rect 174412 76780 174418 76832
rect 174446 76780 174452 76832
rect 174504 76820 174510 76832
rect 373994 76820 374000 76832
rect 174504 76792 374000 76820
rect 174504 76780 174510 76792
rect 373994 76780 374000 76792
rect 374052 76780 374058 76832
rect 155092 76724 166994 76752
rect 155092 76712 155098 76724
rect 171226 76712 171232 76764
rect 171284 76752 171290 76764
rect 408494 76752 408500 76764
rect 171284 76724 408500 76752
rect 171284 76712 171290 76724
rect 408494 76712 408500 76724
rect 408552 76712 408558 76764
rect 93854 76644 93860 76696
rect 93912 76684 93918 76696
rect 132494 76684 132500 76696
rect 93912 76656 132500 76684
rect 93912 76644 93918 76656
rect 132494 76644 132500 76656
rect 132552 76644 132558 76696
rect 142614 76644 142620 76696
rect 142672 76684 142678 76696
rect 144546 76684 144552 76696
rect 142672 76656 144552 76684
rect 142672 76644 142678 76656
rect 144546 76644 144552 76656
rect 144604 76644 144610 76696
rect 159450 76644 159456 76696
rect 159508 76684 159514 76696
rect 433334 76684 433340 76696
rect 159508 76656 433340 76684
rect 159508 76644 159514 76656
rect 433334 76644 433340 76656
rect 433392 76644 433398 76696
rect 69014 76576 69020 76628
rect 69072 76616 69078 76628
rect 130746 76616 130752 76628
rect 69072 76588 130752 76616
rect 69072 76576 69078 76588
rect 130746 76576 130752 76588
rect 130804 76576 130810 76628
rect 165798 76576 165804 76628
rect 165856 76616 165862 76628
rect 166074 76616 166080 76628
rect 165856 76588 166080 76616
rect 165856 76576 165862 76588
rect 166074 76576 166080 76588
rect 166132 76576 166138 76628
rect 169110 76576 169116 76628
rect 169168 76616 169174 76628
rect 169478 76616 169484 76628
rect 169168 76588 169484 76616
rect 169168 76576 169174 76588
rect 169478 76576 169484 76588
rect 169536 76576 169542 76628
rect 171778 76576 171784 76628
rect 171836 76616 171842 76628
rect 471974 76616 471980 76628
rect 171836 76588 471980 76616
rect 171836 76576 171842 76588
rect 471974 76576 471980 76588
rect 472032 76576 472038 76628
rect 6914 76508 6920 76560
rect 6972 76548 6978 76560
rect 125134 76548 125140 76560
rect 6972 76520 125140 76548
rect 6972 76508 6978 76520
rect 125134 76508 125140 76520
rect 125192 76508 125198 76560
rect 169202 76508 169208 76560
rect 169260 76548 169266 76560
rect 558914 76548 558920 76560
rect 169260 76520 558920 76548
rect 169260 76508 169266 76520
rect 558914 76508 558920 76520
rect 558972 76508 558978 76560
rect 155218 76440 155224 76492
rect 155276 76480 155282 76492
rect 208394 76480 208400 76492
rect 155276 76452 208400 76480
rect 155276 76440 155282 76452
rect 208394 76440 208400 76452
rect 208452 76440 208458 76492
rect 149054 76372 149060 76424
rect 149112 76412 149118 76424
rect 149514 76412 149520 76424
rect 149112 76384 149520 76412
rect 149112 76372 149118 76384
rect 149514 76372 149520 76384
rect 149572 76372 149578 76424
rect 151630 76372 151636 76424
rect 151688 76412 151694 76424
rect 197354 76412 197360 76424
rect 151688 76384 197360 76412
rect 151688 76372 151694 76384
rect 197354 76372 197360 76384
rect 197412 76372 197418 76424
rect 127434 76304 127440 76356
rect 127492 76344 127498 76356
rect 128078 76344 128084 76356
rect 127492 76316 128084 76344
rect 127492 76304 127498 76316
rect 128078 76304 128084 76316
rect 128136 76304 128142 76356
rect 149422 76304 149428 76356
rect 149480 76344 149486 76356
rect 149974 76344 149980 76356
rect 149480 76316 149980 76344
rect 149480 76304 149486 76316
rect 149974 76304 149980 76316
rect 150032 76304 150038 76356
rect 155678 76304 155684 76356
rect 155736 76344 155742 76356
rect 172514 76344 172520 76356
rect 155736 76316 172520 76344
rect 155736 76304 155742 76316
rect 172514 76304 172520 76316
rect 172572 76304 172578 76356
rect 162486 76236 162492 76288
rect 162544 76276 162550 76288
rect 171778 76276 171784 76288
rect 162544 76248 171784 76276
rect 162544 76236 162550 76248
rect 171778 76236 171784 76248
rect 171836 76236 171842 76288
rect 165890 76168 165896 76220
rect 165948 76208 165954 76220
rect 166166 76208 166172 76220
rect 165948 76180 166172 76208
rect 165948 76168 165954 76180
rect 166166 76168 166172 76180
rect 166224 76168 166230 76220
rect 125134 76032 125140 76084
rect 125192 76072 125198 76084
rect 132402 76072 132408 76084
rect 125192 76044 132408 76072
rect 125192 76032 125198 76044
rect 132402 76032 132408 76044
rect 132460 76032 132466 76084
rect 136082 76032 136088 76084
rect 136140 76072 136146 76084
rect 136450 76072 136456 76084
rect 136140 76044 136456 76072
rect 136140 76032 136146 76044
rect 136450 76032 136456 76044
rect 136508 76032 136514 76084
rect 165890 76032 165896 76084
rect 165948 76072 165954 76084
rect 166534 76072 166540 76084
rect 165948 76044 166540 76072
rect 165948 76032 165954 76044
rect 166534 76032 166540 76044
rect 166592 76032 166598 76084
rect 128538 75964 128544 76016
rect 128596 76004 128602 76016
rect 129090 76004 129096 76016
rect 128596 75976 129096 76004
rect 128596 75964 128602 75976
rect 129090 75964 129096 75976
rect 129148 75964 129154 76016
rect 133874 75964 133880 76016
rect 133932 76004 133938 76016
rect 135530 76004 135536 76016
rect 133932 75976 135536 76004
rect 133932 75964 133938 75976
rect 135530 75964 135536 75976
rect 135588 75964 135594 76016
rect 151722 75896 151728 75948
rect 151780 75936 151786 75948
rect 154850 75936 154856 75948
rect 151780 75908 154856 75936
rect 151780 75896 151786 75908
rect 154850 75896 154856 75908
rect 154908 75896 154914 75948
rect 173250 75936 173256 75948
rect 172440 75908 173256 75936
rect 139946 75828 139952 75880
rect 140004 75868 140010 75880
rect 172440 75868 172468 75908
rect 173250 75896 173256 75908
rect 173308 75896 173314 75948
rect 140004 75840 172468 75868
rect 140004 75828 140010 75840
rect 172514 75828 172520 75880
rect 172572 75868 172578 75880
rect 243722 75868 243728 75880
rect 172572 75840 243728 75868
rect 172572 75828 172578 75840
rect 243722 75828 243728 75840
rect 243780 75828 243786 75880
rect 156782 75760 156788 75812
rect 156840 75800 156846 75812
rect 229186 75800 229192 75812
rect 156840 75772 229192 75800
rect 156840 75760 156846 75772
rect 229186 75760 229192 75772
rect 229244 75760 229250 75812
rect 130470 75692 130476 75744
rect 130528 75732 130534 75744
rect 135254 75732 135260 75744
rect 130528 75704 135260 75732
rect 130528 75692 130534 75704
rect 135254 75692 135260 75704
rect 135312 75692 135318 75744
rect 150618 75692 150624 75744
rect 150676 75732 150682 75744
rect 258074 75732 258080 75744
rect 150676 75704 258080 75732
rect 150676 75692 150682 75704
rect 258074 75692 258080 75704
rect 258132 75692 258138 75744
rect 128630 75624 128636 75676
rect 128688 75664 128694 75676
rect 129550 75664 129556 75676
rect 128688 75636 129556 75664
rect 128688 75624 128694 75636
rect 129550 75624 129556 75636
rect 129608 75624 129614 75676
rect 151078 75624 151084 75676
rect 151136 75664 151142 75676
rect 259454 75664 259460 75676
rect 151136 75636 259460 75664
rect 151136 75624 151142 75636
rect 259454 75624 259460 75636
rect 259512 75624 259518 75676
rect 154574 75556 154580 75608
rect 154632 75596 154638 75608
rect 288526 75596 288532 75608
rect 154632 75568 288532 75596
rect 154632 75556 154638 75568
rect 288526 75556 288532 75568
rect 288584 75556 288590 75608
rect 121454 75488 121460 75540
rect 121512 75528 121518 75540
rect 135070 75528 135076 75540
rect 121512 75500 135076 75528
rect 121512 75488 121518 75500
rect 135070 75488 135076 75500
rect 135128 75488 135134 75540
rect 151354 75488 151360 75540
rect 151412 75528 151418 75540
rect 288434 75528 288440 75540
rect 151412 75500 288440 75528
rect 151412 75488 151418 75500
rect 288434 75488 288440 75500
rect 288492 75488 288498 75540
rect 51074 75420 51080 75472
rect 51132 75460 51138 75472
rect 129366 75460 129372 75472
rect 51132 75432 129372 75460
rect 51132 75420 51138 75432
rect 129366 75420 129372 75432
rect 129424 75420 129430 75472
rect 129734 75420 129740 75472
rect 129792 75460 129798 75472
rect 135714 75460 135720 75472
rect 129792 75432 135720 75460
rect 129792 75420 129798 75432
rect 135714 75420 135720 75432
rect 135772 75420 135778 75472
rect 156138 75420 156144 75472
rect 156196 75460 156202 75472
rect 340138 75460 340144 75472
rect 156196 75432 340144 75460
rect 156196 75420 156202 75432
rect 340138 75420 340144 75432
rect 340196 75420 340202 75472
rect 107654 75352 107660 75404
rect 107712 75392 107718 75404
rect 133782 75392 133788 75404
rect 107712 75364 133788 75392
rect 107712 75352 107718 75364
rect 133782 75352 133788 75364
rect 133840 75352 133846 75404
rect 134150 75352 134156 75404
rect 134208 75392 134214 75404
rect 134610 75392 134616 75404
rect 134208 75364 134616 75392
rect 134208 75352 134214 75364
rect 134610 75352 134616 75364
rect 134668 75352 134674 75404
rect 155678 75352 155684 75404
rect 155736 75392 155742 75404
rect 359366 75392 359372 75404
rect 155736 75364 359372 75392
rect 155736 75352 155742 75364
rect 359366 75352 359372 75364
rect 359424 75352 359430 75404
rect 49694 75284 49700 75336
rect 49752 75324 49758 75336
rect 129458 75324 129464 75336
rect 49752 75296 129464 75324
rect 49752 75284 49758 75296
rect 129458 75284 129464 75296
rect 129516 75284 129522 75336
rect 131206 75284 131212 75336
rect 131264 75324 131270 75336
rect 132310 75324 132316 75336
rect 131264 75296 132316 75324
rect 131264 75284 131270 75296
rect 132310 75284 132316 75296
rect 132368 75284 132374 75336
rect 135530 75284 135536 75336
rect 135588 75324 135594 75336
rect 136266 75324 136272 75336
rect 135588 75296 136272 75324
rect 135588 75284 135594 75296
rect 136266 75284 136272 75296
rect 136324 75284 136330 75336
rect 143810 75284 143816 75336
rect 143868 75324 143874 75336
rect 144270 75324 144276 75336
rect 143868 75296 144276 75324
rect 143868 75284 143874 75296
rect 144270 75284 144276 75296
rect 144328 75284 144334 75336
rect 149238 75284 149244 75336
rect 149296 75324 149302 75336
rect 150158 75324 150164 75336
rect 149296 75296 150164 75324
rect 149296 75284 149302 75296
rect 150158 75284 150164 75296
rect 150216 75284 150222 75336
rect 157426 75284 157432 75336
rect 157484 75324 157490 75336
rect 158162 75324 158168 75336
rect 157484 75296 158168 75324
rect 157484 75284 157490 75296
rect 158162 75284 158168 75296
rect 158220 75284 158226 75336
rect 163590 75284 163596 75336
rect 163648 75324 163654 75336
rect 163648 75296 165108 75324
rect 163648 75284 163654 75296
rect 46934 75216 46940 75268
rect 46992 75256 46998 75268
rect 124674 75256 124680 75268
rect 46992 75228 124680 75256
rect 46992 75216 46998 75228
rect 124674 75216 124680 75228
rect 124732 75216 124738 75268
rect 129918 75216 129924 75268
rect 129976 75256 129982 75268
rect 130378 75256 130384 75268
rect 129976 75228 130384 75256
rect 129976 75216 129982 75228
rect 130378 75216 130384 75228
rect 130436 75216 130442 75268
rect 131482 75216 131488 75268
rect 131540 75256 131546 75268
rect 131850 75256 131856 75268
rect 131540 75228 131856 75256
rect 131540 75216 131546 75228
rect 131850 75216 131856 75228
rect 131908 75216 131914 75268
rect 132678 75216 132684 75268
rect 132736 75256 132742 75268
rect 133598 75256 133604 75268
rect 132736 75228 133604 75256
rect 132736 75216 132742 75228
rect 133598 75216 133604 75228
rect 133656 75216 133662 75268
rect 134610 75216 134616 75268
rect 134668 75256 134674 75268
rect 135162 75256 135168 75268
rect 134668 75228 135168 75256
rect 134668 75216 134674 75228
rect 135162 75216 135168 75228
rect 135220 75216 135226 75268
rect 135990 75216 135996 75268
rect 136048 75256 136054 75268
rect 136542 75256 136548 75268
rect 136048 75228 136548 75256
rect 136048 75216 136054 75228
rect 136542 75216 136548 75228
rect 136600 75216 136606 75268
rect 137094 75216 137100 75268
rect 137152 75256 137158 75268
rect 137278 75256 137284 75268
rect 137152 75228 137284 75256
rect 137152 75216 137158 75228
rect 137278 75216 137284 75228
rect 137336 75216 137342 75268
rect 138106 75216 138112 75268
rect 138164 75256 138170 75268
rect 138290 75256 138296 75268
rect 138164 75228 138296 75256
rect 138164 75216 138170 75228
rect 138290 75216 138296 75228
rect 138348 75216 138354 75268
rect 138842 75216 138848 75268
rect 138900 75256 138906 75268
rect 139026 75256 139032 75268
rect 138900 75228 139032 75256
rect 138900 75216 138906 75228
rect 139026 75216 139032 75228
rect 139084 75216 139090 75268
rect 139946 75216 139952 75268
rect 140004 75256 140010 75268
rect 140222 75256 140228 75268
rect 140004 75228 140228 75256
rect 140004 75216 140010 75228
rect 140222 75216 140228 75228
rect 140280 75216 140286 75268
rect 141050 75216 141056 75268
rect 141108 75256 141114 75268
rect 141326 75256 141332 75268
rect 141108 75228 141332 75256
rect 141108 75216 141114 75228
rect 141326 75216 141332 75228
rect 141384 75216 141390 75268
rect 142614 75216 142620 75268
rect 142672 75256 142678 75268
rect 142982 75256 142988 75268
rect 142672 75228 142988 75256
rect 142672 75216 142678 75228
rect 142982 75216 142988 75228
rect 143040 75216 143046 75268
rect 145098 75216 145104 75268
rect 145156 75256 145162 75268
rect 145282 75256 145288 75268
rect 145156 75228 145288 75256
rect 145156 75216 145162 75228
rect 145282 75216 145288 75228
rect 145340 75216 145346 75268
rect 145466 75216 145472 75268
rect 145524 75256 145530 75268
rect 145650 75256 145656 75268
rect 145524 75228 145656 75256
rect 145524 75216 145530 75228
rect 145650 75216 145656 75228
rect 145708 75216 145714 75268
rect 146386 75216 146392 75268
rect 146444 75256 146450 75268
rect 146662 75256 146668 75268
rect 146444 75228 146668 75256
rect 146444 75216 146450 75228
rect 146662 75216 146668 75228
rect 146720 75216 146726 75268
rect 146754 75216 146760 75268
rect 146812 75256 146818 75268
rect 146938 75256 146944 75268
rect 146812 75228 146944 75256
rect 146812 75216 146818 75228
rect 146938 75216 146944 75228
rect 146996 75216 147002 75268
rect 147950 75216 147956 75268
rect 148008 75256 148014 75268
rect 148594 75256 148600 75268
rect 148008 75228 148600 75256
rect 148008 75216 148014 75228
rect 148594 75216 148600 75228
rect 148652 75216 148658 75268
rect 149330 75216 149336 75268
rect 149388 75256 149394 75268
rect 149790 75256 149796 75268
rect 149388 75228 149796 75256
rect 149388 75216 149394 75228
rect 149790 75216 149796 75228
rect 149848 75216 149854 75268
rect 151998 75216 152004 75268
rect 152056 75256 152062 75268
rect 152458 75256 152464 75268
rect 152056 75228 152464 75256
rect 152056 75216 152062 75228
rect 152458 75216 152464 75228
rect 152516 75216 152522 75268
rect 157518 75216 157524 75268
rect 157576 75256 157582 75268
rect 157794 75256 157800 75268
rect 157576 75228 157800 75256
rect 157576 75216 157582 75228
rect 157794 75216 157800 75228
rect 157852 75216 157858 75268
rect 158898 75216 158904 75268
rect 158956 75256 158962 75268
rect 159082 75256 159088 75268
rect 158956 75228 159088 75256
rect 158956 75216 158962 75228
rect 159082 75216 159088 75228
rect 159140 75216 159146 75268
rect 160002 75216 160008 75268
rect 160060 75256 160066 75268
rect 160830 75256 160836 75268
rect 160060 75228 160836 75256
rect 160060 75216 160066 75228
rect 160830 75216 160836 75228
rect 160888 75216 160894 75268
rect 163222 75216 163228 75268
rect 163280 75256 163286 75268
rect 163682 75256 163688 75268
rect 163280 75228 163688 75256
rect 163280 75216 163286 75228
rect 163682 75216 163688 75228
rect 163740 75216 163746 75268
rect 164418 75216 164424 75268
rect 164476 75256 164482 75268
rect 164970 75256 164976 75268
rect 164476 75228 164976 75256
rect 164476 75216 164482 75228
rect 164970 75216 164976 75228
rect 165028 75216 165034 75268
rect 165080 75256 165108 75296
rect 165430 75284 165436 75336
rect 165488 75324 165494 75336
rect 481634 75324 481640 75336
rect 165488 75296 481640 75324
rect 165488 75284 165494 75296
rect 481634 75284 481640 75296
rect 481692 75284 481698 75336
rect 489914 75256 489920 75268
rect 165080 75228 489920 75256
rect 489914 75216 489920 75228
rect 489972 75216 489978 75268
rect 26234 75148 26240 75200
rect 26292 75188 26298 75200
rect 26292 75160 118694 75188
rect 26292 75148 26298 75160
rect 118666 74984 118694 75160
rect 125962 75148 125968 75200
rect 126020 75188 126026 75200
rect 126606 75188 126612 75200
rect 126020 75160 126612 75188
rect 126020 75148 126026 75160
rect 126606 75148 126612 75160
rect 126664 75148 126670 75200
rect 130010 75148 130016 75200
rect 130068 75188 130074 75200
rect 130654 75188 130660 75200
rect 130068 75160 130660 75188
rect 130068 75148 130074 75160
rect 130654 75148 130660 75160
rect 130712 75148 130718 75200
rect 131298 75148 131304 75200
rect 131356 75188 131362 75200
rect 131574 75188 131580 75200
rect 131356 75160 131580 75188
rect 131356 75148 131362 75160
rect 131574 75148 131580 75160
rect 131632 75148 131638 75200
rect 135714 75148 135720 75200
rect 135772 75188 135778 75200
rect 136358 75188 136364 75200
rect 135772 75160 136364 75188
rect 135772 75148 135778 75160
rect 136358 75148 136364 75160
rect 136416 75148 136422 75200
rect 139670 75148 139676 75200
rect 139728 75188 139734 75200
rect 140314 75188 140320 75200
rect 139728 75160 140320 75188
rect 139728 75148 139734 75160
rect 140314 75148 140320 75160
rect 140372 75148 140378 75200
rect 142246 75148 142252 75200
rect 142304 75188 142310 75200
rect 142890 75188 142896 75200
rect 142304 75160 142896 75188
rect 142304 75148 142310 75160
rect 142890 75148 142896 75160
rect 142948 75148 142954 75200
rect 143994 75148 144000 75200
rect 144052 75188 144058 75200
rect 144454 75188 144460 75200
rect 144052 75160 144460 75188
rect 144052 75148 144058 75160
rect 144454 75148 144460 75160
rect 144512 75148 144518 75200
rect 147766 75148 147772 75200
rect 147824 75188 147830 75200
rect 148686 75188 148692 75200
rect 147824 75160 148692 75188
rect 147824 75148 147830 75160
rect 148686 75148 148692 75160
rect 148744 75148 148750 75200
rect 149422 75148 149428 75200
rect 149480 75188 149486 75200
rect 149882 75188 149888 75200
rect 149480 75160 149888 75188
rect 149480 75148 149486 75160
rect 149882 75148 149888 75160
rect 149940 75148 149946 75200
rect 151906 75148 151912 75200
rect 151964 75188 151970 75200
rect 152366 75188 152372 75200
rect 151964 75160 152372 75188
rect 151964 75148 151970 75160
rect 152366 75148 152372 75160
rect 152424 75148 152430 75200
rect 152476 75160 157472 75188
rect 126054 75080 126060 75132
rect 126112 75120 126118 75132
rect 126882 75120 126888 75132
rect 126112 75092 126888 75120
rect 126112 75080 126118 75092
rect 126882 75080 126888 75092
rect 126940 75080 126946 75132
rect 132954 75080 132960 75132
rect 133012 75120 133018 75132
rect 133322 75120 133328 75132
rect 133012 75092 133328 75120
rect 133012 75080 133018 75092
rect 133322 75080 133328 75092
rect 133380 75080 133386 75132
rect 138290 75080 138296 75132
rect 138348 75120 138354 75132
rect 138750 75120 138756 75132
rect 138348 75092 138756 75120
rect 138348 75080 138354 75092
rect 138750 75080 138756 75092
rect 138808 75080 138814 75132
rect 141050 75080 141056 75132
rect 141108 75120 141114 75132
rect 141786 75120 141792 75132
rect 141108 75092 141792 75120
rect 141108 75080 141114 75092
rect 141786 75080 141792 75092
rect 141844 75080 141850 75132
rect 145098 75080 145104 75132
rect 145156 75120 145162 75132
rect 145926 75120 145932 75132
rect 145156 75092 145932 75120
rect 145156 75080 145162 75092
rect 145926 75080 145932 75092
rect 145984 75080 145990 75132
rect 146570 75080 146576 75132
rect 146628 75120 146634 75132
rect 146938 75120 146944 75132
rect 146628 75092 146944 75120
rect 146628 75080 146634 75092
rect 146938 75080 146944 75092
rect 146996 75080 147002 75132
rect 149146 75080 149152 75132
rect 149204 75120 149210 75132
rect 152476 75120 152504 75160
rect 149204 75092 152504 75120
rect 149204 75080 149210 75092
rect 156690 75080 156696 75132
rect 156748 75120 156754 75132
rect 156748 75092 157334 75120
rect 156748 75080 156754 75092
rect 131574 75012 131580 75064
rect 131632 75052 131638 75064
rect 132126 75052 132132 75064
rect 131632 75024 132132 75052
rect 131632 75012 131638 75024
rect 132126 75012 132132 75024
rect 132184 75012 132190 75064
rect 136910 75012 136916 75064
rect 136968 75052 136974 75064
rect 137554 75052 137560 75064
rect 136968 75024 137560 75052
rect 136968 75012 136974 75024
rect 137554 75012 137560 75024
rect 137612 75012 137618 75064
rect 143534 75012 143540 75064
rect 143592 75052 143598 75064
rect 144362 75052 144368 75064
rect 143592 75024 144368 75052
rect 143592 75012 143598 75024
rect 144362 75012 144368 75024
rect 144420 75012 144426 75064
rect 146662 75012 146668 75064
rect 146720 75052 146726 75064
rect 147490 75052 147496 75064
rect 146720 75024 147496 75052
rect 146720 75012 146726 75024
rect 147490 75012 147496 75024
rect 147548 75012 147554 75064
rect 124398 74984 124404 74996
rect 118666 74956 124404 74984
rect 124398 74944 124404 74956
rect 124456 74944 124462 74996
rect 127250 74944 127256 74996
rect 127308 74984 127314 74996
rect 127618 74984 127624 74996
rect 127308 74956 127624 74984
rect 127308 74944 127314 74956
rect 127618 74944 127624 74956
rect 127676 74944 127682 74996
rect 128446 74944 128452 74996
rect 128504 74984 128510 74996
rect 128906 74984 128912 74996
rect 128504 74956 128912 74984
rect 128504 74944 128510 74956
rect 128906 74944 128912 74956
rect 128964 74944 128970 74996
rect 137002 74944 137008 74996
rect 137060 74984 137066 74996
rect 137738 74984 137744 74996
rect 137060 74956 137744 74984
rect 137060 74944 137066 74956
rect 137738 74944 137744 74956
rect 137796 74944 137802 74996
rect 146570 74944 146576 74996
rect 146628 74984 146634 74996
rect 147214 74984 147220 74996
rect 146628 74956 147220 74984
rect 146628 74944 146634 74956
rect 147214 74944 147220 74956
rect 147272 74944 147278 74996
rect 151906 74876 151912 74928
rect 151964 74916 151970 74928
rect 153102 74916 153108 74928
rect 151964 74888 153108 74916
rect 151964 74876 151970 74888
rect 153102 74876 153108 74888
rect 153160 74876 153166 74928
rect 157306 74916 157334 75092
rect 157444 74984 157472 75160
rect 157610 75148 157616 75200
rect 157668 75188 157674 75200
rect 158070 75188 158076 75200
rect 157668 75160 158076 75188
rect 157668 75148 157674 75160
rect 158070 75148 158076 75160
rect 158128 75148 158134 75200
rect 162946 75148 162952 75200
rect 163004 75188 163010 75200
rect 163774 75188 163780 75200
rect 163004 75160 163780 75188
rect 163004 75148 163010 75160
rect 163774 75148 163780 75160
rect 163832 75148 163838 75200
rect 164510 75148 164516 75200
rect 164568 75188 164574 75200
rect 165154 75188 165160 75200
rect 164568 75160 165160 75188
rect 164568 75148 164574 75160
rect 165154 75148 165160 75160
rect 165212 75148 165218 75200
rect 506474 75188 506480 75200
rect 166966 75160 506480 75188
rect 157518 75080 157524 75132
rect 157576 75120 157582 75132
rect 157978 75120 157984 75132
rect 157576 75092 157984 75120
rect 157576 75080 157582 75092
rect 157978 75080 157984 75092
rect 158036 75080 158042 75132
rect 163038 75080 163044 75132
rect 163096 75120 163102 75132
rect 163866 75120 163872 75132
rect 163096 75092 163872 75120
rect 163096 75080 163102 75092
rect 163866 75080 163872 75092
rect 163924 75080 163930 75132
rect 163682 74984 163688 74996
rect 157444 74956 163688 74984
rect 163682 74944 163688 74956
rect 163740 74944 163746 74996
rect 164878 74944 164884 74996
rect 164936 74984 164942 74996
rect 166966 74984 166994 75160
rect 506474 75148 506480 75160
rect 506532 75148 506538 75200
rect 169754 75080 169760 75132
rect 169812 75120 169818 75132
rect 170122 75120 170128 75132
rect 169812 75092 170128 75120
rect 169812 75080 169818 75092
rect 170122 75080 170128 75092
rect 170180 75080 170186 75132
rect 171502 75012 171508 75064
rect 171560 75052 171566 75064
rect 172422 75052 172428 75064
rect 171560 75024 172428 75052
rect 171560 75012 171566 75024
rect 172422 75012 172428 75024
rect 172480 75012 172486 75064
rect 164936 74956 166994 74984
rect 164936 74944 164942 74956
rect 173526 74916 173532 74928
rect 157306 74888 173532 74916
rect 173526 74876 173532 74888
rect 173584 74876 173590 74928
rect 151814 74808 151820 74860
rect 151872 74848 151878 74860
rect 152642 74848 152648 74860
rect 151872 74820 152648 74848
rect 151872 74808 151878 74820
rect 152642 74808 152648 74820
rect 152700 74808 152706 74860
rect 127342 74672 127348 74724
rect 127400 74712 127406 74724
rect 128170 74712 128176 74724
rect 127400 74684 128176 74712
rect 127400 74672 127406 74684
rect 128170 74672 128176 74684
rect 128228 74672 128234 74724
rect 139118 74468 139124 74520
rect 139176 74508 139182 74520
rect 140130 74508 140136 74520
rect 139176 74480 140136 74508
rect 139176 74468 139182 74480
rect 140130 74468 140136 74480
rect 140188 74468 140194 74520
rect 143074 74468 143080 74520
rect 143132 74508 143138 74520
rect 223574 74508 223580 74520
rect 143132 74480 223580 74508
rect 143132 74468 143138 74480
rect 223574 74468 223580 74480
rect 223632 74468 223638 74520
rect 243722 74468 243728 74520
rect 243780 74508 243786 74520
rect 347498 74508 347504 74520
rect 243780 74480 347504 74508
rect 243780 74468 243786 74480
rect 347498 74468 347504 74480
rect 347556 74468 347562 74520
rect 145742 74400 145748 74452
rect 145800 74440 145806 74452
rect 251174 74440 251180 74452
rect 145800 74412 251180 74440
rect 145800 74400 145806 74412
rect 251174 74400 251180 74412
rect 251232 74400 251238 74452
rect 156230 74332 156236 74384
rect 156288 74372 156294 74384
rect 270034 74372 270040 74384
rect 156288 74344 270040 74372
rect 156288 74332 156294 74344
rect 270034 74332 270040 74344
rect 270092 74332 270098 74384
rect 151538 74264 151544 74316
rect 151596 74304 151602 74316
rect 189074 74304 189080 74316
rect 151596 74276 189080 74304
rect 151596 74264 151602 74276
rect 189074 74264 189080 74276
rect 189132 74264 189138 74316
rect 208394 74264 208400 74316
rect 208452 74304 208458 74316
rect 322934 74304 322940 74316
rect 208452 74276 322940 74304
rect 208452 74264 208458 74276
rect 322934 74264 322940 74276
rect 322992 74264 322998 74316
rect 156598 74196 156604 74248
rect 156656 74236 156662 74248
rect 301130 74236 301136 74248
rect 156656 74208 301136 74236
rect 156656 74196 156662 74208
rect 301130 74196 301136 74208
rect 301188 74196 301194 74248
rect 128262 74128 128268 74180
rect 128320 74168 128326 74180
rect 229094 74168 229100 74180
rect 128320 74140 229100 74168
rect 128320 74128 128326 74140
rect 229094 74128 229100 74140
rect 229152 74128 229158 74180
rect 229186 74128 229192 74180
rect 229244 74168 229250 74180
rect 382918 74168 382924 74180
rect 229244 74140 382924 74168
rect 229244 74128 229250 74140
rect 382918 74128 382924 74140
rect 382976 74128 382982 74180
rect 4154 74060 4160 74112
rect 4212 74100 4218 74112
rect 125594 74100 125600 74112
rect 4212 74072 125600 74100
rect 4212 74060 4218 74072
rect 125594 74060 125600 74072
rect 125652 74060 125658 74112
rect 154298 74060 154304 74112
rect 154356 74100 154362 74112
rect 318794 74100 318800 74112
rect 154356 74072 318800 74100
rect 154356 74060 154362 74072
rect 318794 74060 318800 74072
rect 318852 74060 318858 74112
rect 118786 73992 118792 74044
rect 118844 74032 118850 74044
rect 134702 74032 134708 74044
rect 118844 74004 134708 74032
rect 118844 73992 118850 74004
rect 134702 73992 134708 74004
rect 134760 73992 134766 74044
rect 157242 73992 157248 74044
rect 157300 74032 157306 74044
rect 324314 74032 324320 74044
rect 157300 74004 324320 74032
rect 157300 73992 157306 74004
rect 324314 73992 324320 74004
rect 324372 73992 324378 74044
rect 60734 73924 60740 73976
rect 60792 73964 60798 73976
rect 130194 73964 130200 73976
rect 60792 73936 130200 73964
rect 60792 73924 60798 73936
rect 130194 73924 130200 73936
rect 130252 73924 130258 73976
rect 156966 73924 156972 73976
rect 157024 73964 157030 73976
rect 331858 73964 331864 73976
rect 157024 73936 331864 73964
rect 157024 73924 157030 73936
rect 331858 73924 331864 73936
rect 331916 73924 331922 73976
rect 30374 73856 30380 73908
rect 30432 73896 30438 73908
rect 30432 73868 118694 73896
rect 30432 73856 30438 73868
rect 118666 73828 118694 73868
rect 126330 73856 126336 73908
rect 126388 73896 126394 73908
rect 126790 73896 126796 73908
rect 126388 73868 126796 73896
rect 126388 73856 126394 73868
rect 126790 73856 126796 73868
rect 126848 73856 126854 73908
rect 156414 73856 156420 73908
rect 156472 73896 156478 73908
rect 362954 73896 362960 73908
rect 156472 73868 362960 73896
rect 156472 73856 156478 73868
rect 362954 73856 362960 73868
rect 363012 73856 363018 73908
rect 127986 73828 127992 73840
rect 118666 73800 127992 73828
rect 127986 73788 127992 73800
rect 128044 73788 128050 73840
rect 158622 73788 158628 73840
rect 158680 73828 158686 73840
rect 368474 73828 368480 73840
rect 158680 73800 368480 73828
rect 158680 73788 158686 73800
rect 368474 73788 368480 73800
rect 368532 73788 368538 73840
rect 141694 73720 141700 73772
rect 141752 73760 141758 73772
rect 209774 73760 209780 73772
rect 141752 73732 209780 73760
rect 141752 73720 141758 73732
rect 209774 73720 209780 73732
rect 209832 73720 209838 73772
rect 193858 73652 193864 73704
rect 193916 73692 193922 73704
rect 214098 73692 214104 73704
rect 193916 73664 214104 73692
rect 193916 73652 193922 73664
rect 214098 73652 214104 73664
rect 214156 73652 214162 73704
rect 369118 73652 369124 73704
rect 369176 73692 369182 73704
rect 374730 73692 374736 73704
rect 369176 73664 374736 73692
rect 369176 73652 369182 73664
rect 374730 73652 374736 73664
rect 374788 73652 374794 73704
rect 137370 73380 137376 73432
rect 137428 73420 137434 73432
rect 142982 73420 142988 73432
rect 137428 73392 142988 73420
rect 137428 73380 137434 73392
rect 142982 73380 142988 73392
rect 143040 73380 143046 73432
rect 339126 73244 339132 73296
rect 339184 73284 339190 73296
rect 341058 73284 341064 73296
rect 339184 73256 341064 73284
rect 339184 73244 339190 73256
rect 341058 73244 341064 73256
rect 341116 73244 341122 73296
rect 126238 73176 126244 73228
rect 126296 73216 126302 73228
rect 130838 73216 130844 73228
rect 126296 73188 130844 73216
rect 126296 73176 126302 73188
rect 130838 73176 130844 73188
rect 130896 73176 130902 73228
rect 151262 73108 151268 73160
rect 151320 73148 151326 73160
rect 155310 73148 155316 73160
rect 151320 73120 155316 73148
rect 151320 73108 151326 73120
rect 155310 73108 155316 73120
rect 155368 73108 155374 73160
rect 170858 73108 170864 73160
rect 170916 73148 170922 73160
rect 580166 73148 580172 73160
rect 170916 73120 580172 73148
rect 170916 73108 170922 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 150710 73040 150716 73092
rect 150768 73080 150774 73092
rect 155770 73080 155776 73092
rect 150768 73052 155776 73080
rect 150768 73040 150774 73052
rect 155770 73040 155776 73052
rect 155828 73040 155834 73092
rect 258074 72836 258080 72888
rect 258132 72876 258138 72888
rect 268194 72876 268200 72888
rect 258132 72848 268200 72876
rect 258132 72836 258138 72848
rect 268194 72836 268200 72848
rect 268252 72836 268258 72888
rect 166718 72768 166724 72820
rect 166776 72808 166782 72820
rect 181438 72808 181444 72820
rect 166776 72780 181444 72808
rect 166776 72768 166782 72780
rect 181438 72768 181444 72780
rect 181496 72768 181502 72820
rect 259454 72768 259460 72820
rect 259512 72808 259518 72820
rect 275370 72808 275376 72820
rect 259512 72780 275376 72808
rect 259512 72768 259518 72780
rect 275370 72768 275376 72780
rect 275428 72768 275434 72820
rect 150894 72700 150900 72752
rect 150952 72740 150958 72752
rect 280062 72740 280068 72752
rect 150952 72712 280068 72740
rect 150952 72700 150958 72712
rect 280062 72700 280068 72712
rect 280120 72700 280126 72752
rect 149974 72632 149980 72684
rect 150032 72672 150038 72684
rect 307754 72672 307760 72684
rect 150032 72644 307760 72672
rect 150032 72632 150038 72644
rect 307754 72632 307760 72644
rect 307812 72632 307818 72684
rect 150066 72564 150072 72616
rect 150124 72604 150130 72616
rect 311894 72604 311900 72616
rect 150124 72576 311900 72604
rect 150124 72564 150130 72576
rect 311894 72564 311900 72576
rect 311952 72564 311958 72616
rect 114554 72496 114560 72548
rect 114612 72536 114618 72548
rect 134426 72536 134432 72548
rect 114612 72508 134432 72536
rect 114612 72496 114618 72508
rect 134426 72496 134432 72508
rect 134484 72496 134490 72548
rect 153194 72496 153200 72548
rect 153252 72536 153258 72548
rect 340874 72536 340880 72548
rect 153252 72508 340880 72536
rect 153252 72496 153258 72508
rect 340874 72496 340880 72508
rect 340932 72496 340938 72548
rect 96614 72428 96620 72480
rect 96672 72468 96678 72480
rect 132586 72468 132592 72480
rect 96672 72440 132592 72468
rect 96672 72428 96678 72440
rect 132586 72428 132592 72440
rect 132644 72428 132650 72480
rect 158346 72428 158352 72480
rect 158404 72468 158410 72480
rect 354674 72468 354680 72480
rect 158404 72440 354680 72468
rect 158404 72428 158410 72440
rect 354674 72428 354680 72440
rect 354732 72428 354738 72480
rect 288434 72156 288440 72208
rect 288492 72196 288498 72208
rect 296162 72196 296168 72208
rect 288492 72168 296168 72196
rect 288492 72156 288498 72168
rect 296162 72156 296168 72168
rect 296220 72156 296226 72208
rect 378410 71748 378416 71800
rect 378468 71788 378474 71800
rect 384758 71788 384764 71800
rect 378468 71760 384764 71788
rect 378468 71748 378474 71760
rect 384758 71748 384764 71760
rect 384816 71748 384822 71800
rect 150986 71680 150992 71732
rect 151044 71720 151050 71732
rect 215294 71720 215300 71732
rect 151044 71692 215300 71720
rect 151044 71680 151050 71692
rect 215294 71680 215300 71692
rect 215352 71680 215358 71732
rect 229094 71680 229100 71732
rect 229152 71720 229158 71732
rect 258718 71720 258724 71732
rect 229152 71692 258724 71720
rect 229152 71680 229158 71692
rect 258718 71680 258724 71692
rect 258776 71680 258782 71732
rect 349798 71680 349804 71732
rect 349856 71720 349862 71732
rect 355502 71720 355508 71732
rect 349856 71692 355508 71720
rect 349856 71680 349862 71692
rect 355502 71680 355508 71692
rect 355560 71680 355566 71732
rect 359366 71680 359372 71732
rect 359424 71720 359430 71732
rect 365070 71720 365076 71732
rect 359424 71692 365076 71720
rect 359424 71680 359430 71692
rect 365070 71680 365076 71692
rect 365128 71680 365134 71732
rect 3418 71612 3424 71664
rect 3476 71652 3482 71664
rect 9030 71652 9036 71664
rect 3476 71624 9036 71652
rect 3476 71612 3482 71624
rect 9030 71612 9036 71624
rect 9088 71612 9094 71664
rect 189074 71612 189080 71664
rect 189132 71652 189138 71664
rect 286318 71652 286324 71664
rect 189132 71624 286324 71652
rect 189132 71612 189138 71624
rect 286318 71612 286324 71624
rect 286376 71612 286382 71664
rect 154666 71544 154672 71596
rect 154724 71584 154730 71596
rect 255314 71584 255320 71596
rect 154724 71556 255320 71584
rect 154724 71544 154730 71556
rect 255314 71544 255320 71556
rect 255372 71544 255378 71596
rect 150802 71476 150808 71528
rect 150860 71516 150866 71528
rect 264238 71516 264244 71528
rect 150860 71488 264244 71516
rect 150860 71476 150866 71488
rect 264238 71476 264244 71488
rect 264296 71476 264302 71528
rect 154850 71408 154856 71460
rect 154908 71448 154914 71460
rect 271874 71448 271880 71460
rect 154908 71420 271880 71448
rect 154908 71408 154914 71420
rect 271874 71408 271880 71420
rect 271932 71408 271938 71460
rect 155494 71340 155500 71392
rect 155552 71380 155558 71392
rect 287606 71380 287612 71392
rect 155552 71352 287612 71380
rect 155552 71340 155558 71352
rect 287606 71340 287612 71352
rect 287664 71340 287670 71392
rect 301130 71340 301136 71392
rect 301188 71380 301194 71392
rect 311158 71380 311164 71392
rect 301188 71352 311164 71380
rect 301188 71340 301194 71352
rect 311158 71340 311164 71352
rect 311216 71340 311222 71392
rect 324314 71340 324320 71392
rect 324372 71380 324378 71392
rect 330478 71380 330484 71392
rect 324372 71352 330484 71380
rect 324372 71340 324378 71352
rect 330478 71340 330484 71352
rect 330536 71340 330542 71392
rect 155402 71272 155408 71324
rect 155460 71312 155466 71324
rect 316678 71312 316684 71324
rect 155460 71284 316684 71312
rect 155460 71272 155466 71284
rect 316678 71272 316684 71284
rect 316736 71272 316742 71324
rect 322934 71272 322940 71324
rect 322992 71312 322998 71324
rect 332594 71312 332600 71324
rect 322992 71284 332600 71312
rect 322992 71272 322998 71284
rect 332594 71272 332600 71284
rect 332652 71272 332658 71324
rect 154758 71204 154764 71256
rect 154816 71244 154822 71256
rect 339402 71244 339408 71256
rect 154816 71216 339408 71244
rect 154816 71204 154822 71216
rect 339402 71204 339408 71216
rect 339460 71204 339466 71256
rect 362954 71204 362960 71256
rect 363012 71244 363018 71256
rect 370498 71244 370504 71256
rect 363012 71216 370504 71244
rect 363012 71204 363018 71216
rect 370498 71204 370504 71216
rect 370556 71204 370562 71256
rect 165062 71136 165068 71188
rect 165120 71176 165126 71188
rect 500954 71176 500960 71188
rect 165120 71148 500960 71176
rect 165120 71136 165126 71148
rect 500954 71136 500960 71148
rect 501012 71136 501018 71188
rect 165522 71068 165528 71120
rect 165580 71108 165586 71120
rect 507854 71108 507860 71120
rect 165580 71080 507860 71108
rect 165580 71068 165586 71080
rect 507854 71068 507860 71080
rect 507912 71068 507918 71120
rect 138014 71000 138020 71052
rect 138072 71040 138078 71052
rect 165062 71040 165068 71052
rect 138072 71012 165068 71040
rect 138072 71000 138078 71012
rect 165062 71000 165068 71012
rect 165120 71000 165126 71052
rect 168006 71000 168012 71052
rect 168064 71040 168070 71052
rect 539594 71040 539600 71052
rect 168064 71012 539600 71040
rect 168064 71000 168070 71012
rect 539594 71000 539600 71012
rect 539652 71000 539658 71052
rect 148410 70932 148416 70984
rect 148468 70972 148474 70984
rect 190454 70972 190460 70984
rect 148468 70944 190460 70972
rect 148468 70932 148474 70944
rect 190454 70932 190460 70944
rect 190512 70932 190518 70984
rect 214098 70932 214104 70984
rect 214156 70972 214162 70984
rect 257338 70972 257344 70984
rect 214156 70944 257344 70972
rect 214156 70932 214162 70944
rect 257338 70932 257344 70944
rect 257396 70932 257402 70984
rect 164050 70524 164056 70576
rect 164108 70564 164114 70576
rect 170398 70564 170404 70576
rect 164108 70536 170404 70564
rect 164108 70524 164114 70536
rect 170398 70524 170404 70536
rect 170456 70524 170462 70576
rect 155310 70320 155316 70372
rect 155368 70360 155374 70372
rect 250438 70360 250444 70372
rect 155368 70332 250444 70360
rect 155368 70320 155374 70332
rect 250438 70320 250444 70332
rect 250496 70320 250502 70372
rect 155770 70252 155776 70304
rect 155828 70292 155834 70304
rect 271782 70292 271788 70304
rect 155828 70264 271788 70292
rect 155828 70252 155834 70264
rect 271782 70252 271788 70264
rect 271840 70252 271846 70304
rect 140038 70184 140044 70236
rect 140096 70224 140102 70236
rect 173434 70224 173440 70236
rect 140096 70196 173440 70224
rect 140096 70184 140102 70196
rect 173434 70184 173440 70196
rect 173492 70184 173498 70236
rect 173526 70184 173532 70236
rect 173584 70224 173590 70236
rect 327718 70224 327724 70236
rect 173584 70196 327724 70224
rect 173584 70184 173590 70196
rect 327718 70184 327724 70196
rect 327776 70184 327782 70236
rect 155954 70116 155960 70168
rect 156012 70156 156018 70168
rect 326982 70156 326988 70168
rect 156012 70128 326988 70156
rect 156012 70116 156018 70128
rect 326982 70116 326988 70128
rect 327040 70116 327046 70168
rect 154666 70048 154672 70100
rect 154724 70088 154730 70100
rect 327810 70088 327816 70100
rect 154724 70060 327816 70088
rect 154724 70048 154730 70060
rect 327810 70048 327816 70060
rect 327868 70048 327874 70100
rect 155862 69980 155868 70032
rect 155920 70020 155926 70032
rect 338758 70020 338764 70032
rect 155920 69992 338764 70020
rect 155920 69980 155926 69992
rect 338758 69980 338764 69992
rect 338816 69980 338822 70032
rect 156874 69912 156880 69964
rect 156932 69952 156938 69964
rect 361574 69952 361580 69964
rect 156932 69924 361580 69952
rect 156932 69912 156938 69924
rect 361574 69912 361580 69924
rect 361632 69912 361638 69964
rect 164786 69844 164792 69896
rect 164844 69884 164850 69896
rect 505094 69884 505100 69896
rect 164844 69856 505100 69884
rect 164844 69844 164850 69856
rect 505094 69844 505100 69856
rect 505152 69844 505158 69896
rect 166350 69776 166356 69828
rect 166408 69816 166414 69828
rect 523034 69816 523040 69828
rect 166408 69788 523040 69816
rect 166408 69776 166414 69788
rect 523034 69776 523040 69788
rect 523092 69776 523098 69828
rect 137278 69708 137284 69760
rect 137336 69748 137342 69760
rect 149146 69748 149152 69760
rect 137336 69720 149152 69748
rect 137336 69708 137342 69720
rect 149146 69708 149152 69720
rect 149204 69708 149210 69760
rect 167086 69708 167092 69760
rect 167144 69748 167150 69760
rect 536834 69748 536840 69760
rect 167144 69720 536840 69748
rect 167144 69708 167150 69720
rect 536834 69708 536840 69720
rect 536892 69708 536898 69760
rect 138566 69640 138572 69692
rect 138624 69680 138630 69692
rect 140222 69680 140228 69692
rect 138624 69652 140228 69680
rect 138624 69640 138630 69652
rect 140222 69640 140228 69652
rect 140280 69640 140286 69692
rect 169110 69640 169116 69692
rect 169168 69680 169174 69692
rect 564434 69680 564440 69692
rect 169168 69652 564440 69680
rect 169168 69640 169174 69652
rect 564434 69640 564440 69652
rect 564492 69640 564498 69692
rect 141510 69572 141516 69624
rect 141568 69612 141574 69624
rect 209866 69612 209872 69624
rect 141568 69584 209872 69612
rect 141568 69572 141574 69584
rect 209866 69572 209872 69584
rect 209924 69572 209930 69624
rect 215294 68960 215300 69012
rect 215352 69000 215358 69012
rect 218146 69000 218152 69012
rect 215352 68972 218152 69000
rect 215352 68960 215358 68972
rect 218146 68960 218152 68972
rect 218204 68960 218210 69012
rect 255314 68960 255320 69012
rect 255372 69000 255378 69012
rect 258810 69000 258816 69012
rect 255372 68972 258816 69000
rect 255372 68960 255378 68972
rect 258810 68960 258816 68972
rect 258868 68960 258874 69012
rect 288526 68960 288532 69012
rect 288584 69000 288590 69012
rect 295334 69000 295340 69012
rect 288584 68972 295340 69000
rect 288584 68960 288590 68972
rect 295334 68960 295340 68972
rect 295392 68960 295398 69012
rect 331122 68960 331128 69012
rect 331180 69000 331186 69012
rect 335998 69000 336004 69012
rect 331180 68972 336004 69000
rect 331180 68960 331186 68972
rect 335998 68960 336004 68972
rect 336056 68960 336062 69012
rect 346394 68960 346400 69012
rect 346452 69000 346458 69012
rect 349798 69000 349804 69012
rect 346452 68972 349804 69000
rect 346452 68960 346458 68972
rect 349798 68960 349804 68972
rect 349856 68960 349862 69012
rect 341058 68620 341064 68672
rect 341116 68660 341122 68672
rect 352558 68660 352564 68672
rect 341116 68632 352564 68660
rect 341116 68620 341122 68632
rect 352558 68620 352564 68632
rect 352616 68620 352622 68672
rect 355502 68620 355508 68672
rect 355560 68660 355566 68672
rect 359274 68660 359280 68672
rect 355560 68632 359280 68660
rect 355560 68620 355566 68632
rect 359274 68620 359280 68632
rect 359332 68620 359338 68672
rect 332594 68552 332600 68604
rect 332652 68592 332658 68604
rect 347222 68592 347228 68604
rect 332652 68564 347228 68592
rect 332652 68552 332658 68564
rect 347222 68552 347228 68564
rect 347280 68552 347286 68604
rect 153746 68484 153752 68536
rect 153804 68524 153810 68536
rect 358814 68524 358820 68536
rect 153804 68496 358820 68524
rect 153804 68484 153810 68496
rect 358814 68484 358820 68496
rect 358872 68484 358878 68536
rect 166258 68416 166264 68468
rect 166316 68456 166322 68468
rect 525794 68456 525800 68468
rect 166316 68428 525800 68456
rect 166316 68416 166322 68428
rect 525794 68416 525800 68428
rect 525852 68416 525858 68468
rect 169018 68348 169024 68400
rect 169076 68388 169082 68400
rect 557534 68388 557540 68400
rect 169076 68360 557540 68388
rect 169076 68348 169082 68360
rect 557534 68348 557540 68360
rect 557592 68348 557598 68400
rect 170766 68280 170772 68332
rect 170824 68320 170830 68332
rect 564526 68320 564532 68332
rect 170824 68292 564532 68320
rect 170824 68280 170830 68292
rect 564526 68280 564532 68292
rect 564584 68280 564590 68332
rect 365070 68212 365076 68264
rect 365128 68252 365134 68264
rect 369118 68252 369124 68264
rect 365128 68224 369124 68252
rect 365128 68212 365134 68224
rect 369118 68212 369124 68224
rect 369176 68212 369182 68264
rect 271874 68144 271880 68196
rect 271932 68184 271938 68196
rect 275278 68184 275284 68196
rect 271932 68156 275284 68184
rect 271932 68144 271938 68156
rect 275278 68144 275284 68156
rect 275336 68144 275342 68196
rect 137186 67532 137192 67584
rect 137244 67572 137250 67584
rect 138658 67572 138664 67584
rect 137244 67544 138664 67572
rect 137244 67532 137250 67544
rect 138658 67532 138664 67544
rect 138716 67532 138722 67584
rect 270034 67532 270040 67584
rect 270092 67572 270098 67584
rect 275186 67572 275192 67584
rect 270092 67544 275192 67572
rect 270092 67532 270098 67544
rect 275186 67532 275192 67544
rect 275244 67532 275250 67584
rect 306926 67532 306932 67584
rect 306984 67572 306990 67584
rect 309778 67572 309784 67584
rect 306984 67544 309784 67572
rect 306984 67532 306990 67544
rect 309778 67532 309784 67544
rect 309836 67532 309842 67584
rect 384758 67532 384764 67584
rect 384816 67572 384822 67584
rect 387058 67572 387064 67584
rect 384816 67544 387064 67572
rect 384816 67532 384822 67544
rect 387058 67532 387064 67544
rect 387116 67532 387122 67584
rect 326982 67464 326988 67516
rect 327040 67504 327046 67516
rect 329098 67504 329104 67516
rect 327040 67476 329104 67504
rect 327040 67464 327046 67476
rect 329098 67464 329104 67476
rect 329156 67464 329162 67516
rect 138474 67056 138480 67108
rect 138532 67096 138538 67108
rect 167086 67096 167092 67108
rect 138532 67068 167092 67096
rect 138532 67056 138538 67068
rect 167086 67056 167092 67068
rect 167144 67056 167150 67108
rect 139946 66988 139952 67040
rect 140004 67028 140010 67040
rect 189074 67028 189080 67040
rect 140004 67000 189080 67028
rect 140004 66988 140010 67000
rect 189074 66988 189080 67000
rect 189132 66988 189138 67040
rect 142798 66920 142804 66972
rect 142856 66960 142862 66972
rect 220814 66960 220820 66972
rect 142856 66932 220820 66960
rect 142856 66920 142862 66932
rect 220814 66920 220820 66932
rect 220872 66920 220878 66972
rect 145558 66852 145564 66904
rect 145616 66892 145622 66904
rect 256694 66892 256700 66904
rect 145616 66864 256700 66892
rect 145616 66852 145622 66864
rect 256694 66852 256700 66864
rect 256752 66852 256758 66904
rect 339402 66716 339408 66768
rect 339460 66756 339466 66768
rect 345658 66756 345664 66768
rect 339460 66728 345664 66756
rect 339460 66716 339466 66728
rect 345658 66716 345664 66728
rect 345716 66716 345722 66768
rect 271782 66444 271788 66496
rect 271840 66484 271846 66496
rect 278774 66484 278780 66496
rect 271840 66456 278780 66484
rect 271840 66444 271846 66456
rect 278774 66444 278780 66456
rect 278832 66444 278838 66496
rect 268194 66172 268200 66224
rect 268252 66212 268258 66224
rect 271138 66212 271144 66224
rect 268252 66184 271144 66212
rect 268252 66172 268258 66184
rect 271138 66172 271144 66184
rect 271196 66172 271202 66224
rect 287606 66172 287612 66224
rect 287664 66212 287670 66224
rect 291102 66212 291108 66224
rect 287664 66184 291108 66212
rect 287664 66172 287670 66184
rect 291102 66172 291108 66184
rect 291160 66172 291166 66224
rect 347498 66172 347504 66224
rect 347556 66212 347562 66224
rect 349982 66212 349988 66224
rect 347556 66184 349988 66212
rect 347556 66172 347562 66184
rect 349982 66172 349988 66184
rect 350040 66172 350046 66224
rect 142706 65764 142712 65816
rect 142764 65804 142770 65816
rect 218054 65804 218060 65816
rect 142764 65776 218060 65804
rect 142764 65764 142770 65776
rect 218054 65764 218060 65776
rect 218112 65764 218118 65816
rect 218146 65764 218152 65816
rect 218204 65804 218210 65816
rect 226242 65804 226248 65816
rect 218204 65776 226248 65804
rect 218204 65764 218210 65776
rect 226242 65764 226248 65776
rect 226300 65764 226306 65816
rect 144178 65696 144184 65748
rect 144236 65736 144242 65748
rect 238754 65736 238760 65748
rect 144236 65708 238760 65736
rect 144236 65696 144242 65708
rect 238754 65696 238760 65708
rect 238812 65696 238818 65748
rect 280062 65696 280068 65748
rect 280120 65736 280126 65748
rect 292850 65736 292856 65748
rect 280120 65708 292856 65736
rect 280120 65696 280126 65708
rect 292850 65696 292856 65708
rect 292908 65696 292914 65748
rect 295334 65696 295340 65748
rect 295392 65736 295398 65748
rect 303614 65736 303620 65748
rect 295392 65708 303620 65736
rect 295392 65696 295398 65708
rect 303614 65696 303620 65708
rect 303672 65696 303678 65748
rect 311158 65696 311164 65748
rect 311216 65736 311222 65748
rect 316034 65736 316040 65748
rect 311216 65708 316040 65736
rect 311216 65696 311222 65708
rect 316034 65696 316040 65708
rect 316092 65696 316098 65748
rect 330478 65696 330484 65748
rect 330536 65736 330542 65748
rect 340782 65736 340788 65748
rect 330536 65708 340788 65736
rect 330536 65696 330542 65708
rect 340782 65696 340788 65708
rect 340840 65696 340846 65748
rect 359274 65696 359280 65748
rect 359332 65736 359338 65748
rect 370958 65736 370964 65748
rect 359332 65708 370964 65736
rect 359332 65696 359338 65708
rect 370958 65696 370964 65708
rect 371016 65696 371022 65748
rect 163406 65628 163412 65680
rect 163464 65668 163470 65680
rect 484394 65668 484400 65680
rect 163464 65640 484400 65668
rect 163464 65628 163470 65640
rect 484394 65628 484400 65640
rect 484452 65628 484458 65680
rect 167730 65560 167736 65612
rect 167788 65600 167794 65612
rect 543734 65600 543740 65612
rect 167788 65572 543740 65600
rect 167788 65560 167794 65572
rect 543734 65560 543740 65572
rect 543792 65560 543798 65612
rect 170214 65492 170220 65544
rect 170272 65532 170278 65544
rect 572714 65532 572720 65544
rect 170272 65504 572720 65532
rect 170272 65492 170278 65504
rect 572714 65492 572720 65504
rect 572772 65492 572778 65544
rect 361574 64880 361580 64932
rect 361632 64920 361638 64932
rect 364978 64920 364984 64932
rect 361632 64892 364984 64920
rect 361632 64880 361638 64892
rect 364978 64880 364984 64892
rect 365036 64880 365042 64932
rect 264238 64404 264244 64456
rect 264296 64444 264302 64456
rect 269758 64444 269764 64456
rect 264296 64416 269764 64444
rect 264296 64404 264302 64416
rect 269758 64404 269764 64416
rect 269816 64404 269822 64456
rect 152550 64268 152556 64320
rect 152608 64308 152614 64320
rect 338114 64308 338120 64320
rect 152608 64280 338120 64308
rect 152608 64268 152614 64280
rect 338114 64268 338120 64280
rect 338172 64268 338178 64320
rect 157978 64200 157984 64252
rect 158036 64240 158042 64252
rect 374086 64240 374092 64252
rect 158036 64212 374092 64240
rect 158036 64200 158042 64212
rect 374086 64200 374092 64212
rect 374144 64200 374150 64252
rect 170122 64132 170128 64184
rect 170180 64172 170186 64184
rect 568574 64172 568580 64184
rect 170180 64144 568580 64172
rect 170180 64132 170186 64144
rect 568574 64132 568580 64144
rect 568632 64132 568638 64184
rect 352558 63996 352564 64048
rect 352616 64036 352622 64048
rect 357342 64036 357348 64048
rect 352616 64008 357348 64036
rect 352616 63996 352622 64008
rect 357342 63996 357348 64008
rect 357400 63996 357406 64048
rect 275370 63724 275376 63776
rect 275428 63764 275434 63776
rect 278406 63764 278412 63776
rect 275428 63736 278412 63764
rect 275428 63724 275434 63736
rect 278406 63724 278412 63736
rect 278464 63724 278470 63776
rect 278774 63588 278780 63640
rect 278832 63628 278838 63640
rect 283006 63628 283012 63640
rect 278832 63600 283012 63628
rect 278832 63588 278838 63600
rect 283006 63588 283012 63600
rect 283064 63588 283070 63640
rect 139854 63112 139860 63164
rect 139912 63152 139918 63164
rect 184934 63152 184940 63164
rect 139912 63124 184940 63152
rect 139912 63112 139918 63124
rect 184934 63112 184940 63124
rect 184992 63112 184998 63164
rect 142614 63044 142620 63096
rect 142672 63084 142678 63096
rect 224954 63084 224960 63096
rect 142672 63056 224960 63084
rect 142672 63044 142678 63056
rect 224954 63044 224960 63056
rect 225012 63044 225018 63096
rect 147122 62976 147128 63028
rect 147180 63016 147186 63028
rect 274634 63016 274640 63028
rect 147180 62988 274640 63016
rect 147180 62976 147186 62988
rect 274634 62976 274640 62988
rect 274692 62976 274698 63028
rect 152458 62908 152464 62960
rect 152516 62948 152522 62960
rect 340966 62948 340972 62960
rect 152516 62920 340972 62948
rect 152516 62908 152522 62920
rect 340966 62908 340972 62920
rect 341024 62908 341030 62960
rect 163314 62840 163320 62892
rect 163372 62880 163378 62892
rect 481726 62880 481732 62892
rect 163372 62852 481732 62880
rect 163372 62840 163378 62852
rect 481726 62840 481732 62852
rect 481784 62840 481790 62892
rect 170674 62772 170680 62824
rect 170732 62812 170738 62824
rect 514754 62812 514760 62824
rect 170732 62784 514760 62812
rect 170732 62772 170738 62784
rect 514754 62772 514760 62784
rect 514812 62772 514818 62824
rect 316034 62568 316040 62620
rect 316092 62608 316098 62620
rect 318978 62608 318984 62620
rect 316092 62580 318984 62608
rect 316092 62568 316098 62580
rect 318978 62568 318984 62580
rect 319036 62568 319042 62620
rect 138382 62024 138388 62076
rect 138440 62064 138446 62076
rect 142798 62064 142804 62076
rect 138440 62036 142804 62064
rect 138440 62024 138446 62036
rect 142798 62024 142804 62036
rect 142856 62024 142862 62076
rect 349982 61956 349988 62008
rect 350040 61996 350046 62008
rect 353938 61996 353944 62008
rect 350040 61968 353944 61996
rect 350040 61956 350046 61968
rect 353938 61956 353944 61968
rect 353996 61956 354002 62008
rect 370958 61752 370964 61804
rect 371016 61792 371022 61804
rect 376662 61792 376668 61804
rect 371016 61764 376668 61792
rect 371016 61752 371022 61764
rect 376662 61752 376668 61764
rect 376720 61752 376726 61804
rect 257338 61616 257344 61668
rect 257396 61656 257402 61668
rect 262858 61656 262864 61668
rect 257396 61628 262864 61656
rect 257396 61616 257402 61628
rect 262858 61616 262864 61628
rect 262916 61616 262922 61668
rect 275186 61616 275192 61668
rect 275244 61656 275250 61668
rect 297358 61656 297364 61668
rect 275244 61628 297364 61656
rect 275244 61616 275250 61628
rect 297358 61616 297364 61628
rect 297416 61616 297422 61668
rect 148318 61548 148324 61600
rect 148376 61588 148382 61600
rect 292574 61588 292580 61600
rect 148376 61560 292580 61588
rect 148376 61548 148382 61560
rect 292574 61548 292580 61560
rect 292632 61548 292638 61600
rect 340782 61548 340788 61600
rect 340840 61588 340846 61600
rect 354030 61588 354036 61600
rect 340840 61560 354036 61588
rect 340840 61548 340846 61560
rect 354030 61548 354036 61560
rect 354088 61548 354094 61600
rect 149698 61480 149704 61532
rect 149756 61520 149762 61532
rect 306374 61520 306380 61532
rect 149756 61492 306380 61520
rect 149756 61480 149762 61492
rect 306374 61480 306380 61492
rect 306432 61480 306438 61532
rect 347222 61480 347228 61532
rect 347280 61520 347286 61532
rect 363598 61520 363604 61532
rect 347280 61492 363604 61520
rect 347280 61480 347286 61492
rect 363598 61480 363604 61492
rect 363656 61480 363662 61532
rect 153654 61412 153660 61464
rect 153712 61452 153718 61464
rect 362954 61452 362960 61464
rect 153712 61424 362960 61452
rect 153712 61412 153718 61424
rect 362954 61412 362960 61424
rect 363012 61412 363018 61464
rect 102226 61344 102232 61396
rect 102284 61384 102290 61396
rect 125318 61384 125324 61396
rect 102284 61356 125324 61384
rect 102284 61344 102290 61356
rect 125318 61344 125324 61356
rect 125376 61344 125382 61396
rect 157886 61344 157892 61396
rect 157944 61384 157950 61396
rect 412634 61384 412640 61396
rect 157944 61356 412640 61384
rect 157944 61344 157950 61356
rect 412634 61344 412640 61356
rect 412692 61344 412698 61396
rect 292850 60936 292856 60988
rect 292908 60976 292914 60988
rect 295978 60976 295984 60988
rect 292908 60948 295984 60976
rect 292908 60936 292914 60948
rect 295978 60936 295984 60948
rect 296036 60936 296042 60988
rect 338758 60732 338764 60784
rect 338816 60772 338822 60784
rect 344278 60772 344284 60784
rect 338816 60744 344284 60772
rect 338816 60732 338822 60744
rect 344278 60732 344284 60744
rect 344336 60732 344342 60784
rect 183278 60664 183284 60716
rect 183336 60704 183342 60716
rect 580166 60704 580172 60716
rect 183336 60676 580172 60704
rect 183336 60664 183342 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 327810 60596 327816 60648
rect 327868 60636 327874 60648
rect 332594 60636 332600 60648
rect 327868 60608 332600 60636
rect 327868 60596 327874 60608
rect 332594 60596 332600 60608
rect 332652 60596 332658 60648
rect 318978 60392 318984 60444
rect 319036 60432 319042 60444
rect 327902 60432 327908 60444
rect 319036 60404 327908 60432
rect 319036 60392 319042 60404
rect 327902 60392 327908 60404
rect 327960 60392 327966 60444
rect 141418 60120 141424 60172
rect 141476 60160 141482 60172
rect 207014 60160 207020 60172
rect 141476 60132 207020 60160
rect 141476 60120 141482 60132
rect 207014 60120 207020 60132
rect 207072 60120 207078 60172
rect 226242 60120 226248 60172
rect 226300 60160 226306 60172
rect 247678 60160 247684 60172
rect 226300 60132 247684 60160
rect 226300 60120 226306 60132
rect 247678 60120 247684 60132
rect 247736 60120 247742 60172
rect 144086 60052 144092 60104
rect 144144 60092 144150 60104
rect 233234 60092 233240 60104
rect 144144 60064 233240 60092
rect 144144 60052 144150 60064
rect 233234 60052 233240 60064
rect 233292 60052 233298 60104
rect 149606 59984 149612 60036
rect 149664 60024 149670 60036
rect 304994 60024 305000 60036
rect 149664 59996 305000 60024
rect 149664 59984 149670 59996
rect 304994 59984 305000 59996
rect 305052 59984 305058 60036
rect 258810 59916 258816 59968
rect 258868 59956 258874 59968
rect 264330 59956 264336 59968
rect 258868 59928 264336 59956
rect 258868 59916 258874 59928
rect 264330 59916 264336 59928
rect 264388 59916 264394 59968
rect 120074 59576 120080 59628
rect 120132 59616 120138 59628
rect 123478 59616 123484 59628
rect 120132 59588 123484 59616
rect 120132 59576 120138 59588
rect 123478 59576 123484 59588
rect 123536 59576 123542 59628
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 181254 59344 181260 59356
rect 3108 59316 181260 59344
rect 3108 59304 3114 59316
rect 181254 59304 181260 59316
rect 181312 59304 181318 59356
rect 258718 59304 258724 59356
rect 258776 59344 258782 59356
rect 261478 59344 261484 59356
rect 258776 59316 261484 59344
rect 258776 59304 258782 59316
rect 261478 59304 261484 59316
rect 261536 59304 261542 59356
rect 303614 59304 303620 59356
rect 303672 59344 303678 59356
rect 307018 59344 307024 59356
rect 303672 59316 307024 59344
rect 303672 59304 303678 59316
rect 307018 59304 307024 59316
rect 307076 59304 307082 59356
rect 357342 59304 357348 59356
rect 357400 59344 357406 59356
rect 363690 59344 363696 59356
rect 357400 59316 363696 59344
rect 357400 59304 357406 59316
rect 363690 59304 363696 59316
rect 363748 59304 363754 59356
rect 286318 58760 286324 58812
rect 286376 58800 286382 58812
rect 298738 58800 298744 58812
rect 286376 58772 298744 58800
rect 286376 58760 286382 58772
rect 298738 58760 298744 58772
rect 298796 58760 298802 58812
rect 283006 58692 283012 58744
rect 283064 58732 283070 58744
rect 291838 58732 291844 58744
rect 283064 58704 291844 58732
rect 283064 58692 283070 58704
rect 291838 58692 291844 58704
rect 291896 58692 291902 58744
rect 296162 58692 296168 58744
rect 296220 58732 296226 58744
rect 313918 58732 313924 58744
rect 296220 58704 313924 58732
rect 296220 58692 296226 58704
rect 313918 58692 313924 58704
rect 313976 58692 313982 58744
rect 275278 58624 275284 58676
rect 275336 58664 275342 58676
rect 283650 58664 283656 58676
rect 275336 58636 283656 58664
rect 275336 58624 275342 58636
rect 283650 58624 283656 58636
rect 283708 58624 283714 58676
rect 291102 58624 291108 58676
rect 291160 58664 291166 58676
rect 311158 58664 311164 58676
rect 291160 58636 311164 58664
rect 291160 58624 291166 58636
rect 311158 58624 311164 58636
rect 311216 58624 311222 58676
rect 335998 58624 336004 58676
rect 336056 58664 336062 58676
rect 362218 58664 362224 58676
rect 336056 58636 362224 58664
rect 336056 58624 336062 58636
rect 362218 58624 362224 58636
rect 362276 58624 362282 58676
rect 95234 57196 95240 57248
rect 95292 57236 95298 57248
rect 125226 57236 125232 57248
rect 95292 57208 125232 57236
rect 95292 57196 95298 57208
rect 125226 57196 125232 57208
rect 125284 57196 125290 57248
rect 296070 57196 296076 57248
rect 296128 57236 296134 57248
rect 301590 57236 301596 57248
rect 296128 57208 301596 57236
rect 296128 57196 296134 57208
rect 301590 57196 301596 57208
rect 301648 57196 301654 57248
rect 309778 57196 309784 57248
rect 309836 57236 309842 57248
rect 323578 57236 323584 57248
rect 309836 57208 323584 57236
rect 309836 57196 309842 57208
rect 323578 57196 323584 57208
rect 323636 57196 323642 57248
rect 376662 57196 376668 57248
rect 376720 57236 376726 57248
rect 384390 57236 384396 57248
rect 376720 57208 384396 57236
rect 376720 57196 376726 57208
rect 384390 57196 384396 57208
rect 384448 57196 384454 57248
rect 332594 56584 332600 56636
rect 332652 56624 332658 56636
rect 335998 56624 336004 56636
rect 332652 56596 336004 56624
rect 332652 56584 332658 56596
rect 335998 56584 336004 56596
rect 336056 56584 336062 56636
rect 261478 56516 261484 56568
rect 261536 56556 261542 56568
rect 264238 56556 264244 56568
rect 261536 56528 264244 56556
rect 261536 56516 261542 56528
rect 264238 56516 264244 56528
rect 264296 56516 264302 56568
rect 278406 56516 278412 56568
rect 278464 56556 278470 56568
rect 280798 56556 280804 56568
rect 278464 56528 280804 56556
rect 278464 56516 278470 56528
rect 280798 56516 280804 56528
rect 280856 56516 280862 56568
rect 329098 56516 329104 56568
rect 329156 56556 329162 56568
rect 333974 56556 333980 56568
rect 329156 56528 333980 56556
rect 329156 56516 329162 56528
rect 333974 56516 333980 56528
rect 334032 56516 334038 56568
rect 369118 56516 369124 56568
rect 369176 56556 369182 56568
rect 371878 56556 371884 56568
rect 369176 56528 371884 56556
rect 369176 56516 369182 56528
rect 371878 56516 371884 56528
rect 371936 56516 371942 56568
rect 88334 55836 88340 55888
rect 88392 55876 88398 55888
rect 125134 55876 125140 55888
rect 88392 55848 125140 55876
rect 88392 55836 88398 55848
rect 125134 55836 125140 55848
rect 125192 55836 125198 55888
rect 370498 55836 370504 55888
rect 370556 55876 370562 55888
rect 387702 55876 387708 55888
rect 370556 55848 387708 55876
rect 370556 55836 370562 55848
rect 387702 55836 387708 55848
rect 387760 55836 387766 55888
rect 291838 54612 291844 54664
rect 291896 54652 291902 54664
rect 295334 54652 295340 54664
rect 291896 54624 295340 54652
rect 291896 54612 291902 54624
rect 295334 54612 295340 54624
rect 295392 54612 295398 54664
rect 283650 54476 283656 54528
rect 283708 54516 283714 54528
rect 292666 54516 292672 54528
rect 283708 54488 292672 54516
rect 283708 54476 283714 54488
rect 292666 54476 292672 54488
rect 292724 54476 292730 54528
rect 297358 54476 297364 54528
rect 297416 54516 297422 54528
rect 326338 54516 326344 54528
rect 297416 54488 326344 54516
rect 297416 54476 297422 54488
rect 326338 54476 326344 54488
rect 326396 54476 326402 54528
rect 340138 54476 340144 54528
rect 340196 54516 340202 54528
rect 343634 54516 343640 54528
rect 340196 54488 343640 54516
rect 340196 54476 340202 54488
rect 343634 54476 343640 54488
rect 343692 54476 343698 54528
rect 364978 54476 364984 54528
rect 365036 54516 365042 54528
rect 374638 54516 374644 54528
rect 365036 54488 374644 54516
rect 365036 54476 365042 54488
rect 374638 54476 374644 54488
rect 374696 54476 374702 54528
rect 262858 54408 262864 54460
rect 262916 54448 262922 54460
rect 269850 54448 269856 54460
rect 262916 54420 269856 54448
rect 262916 54408 262922 54420
rect 269850 54408 269856 54420
rect 269908 54408 269914 54460
rect 250438 54340 250444 54392
rect 250496 54380 250502 54392
rect 253014 54380 253020 54392
rect 250496 54352 253020 54380
rect 250496 54340 250502 54352
rect 253014 54340 253020 54352
rect 253072 54340 253078 54392
rect 374730 54340 374736 54392
rect 374788 54380 374794 54392
rect 380158 54380 380164 54392
rect 374788 54352 380164 54380
rect 374788 54340 374794 54352
rect 380158 54340 380164 54352
rect 380216 54340 380222 54392
rect 363598 53728 363604 53780
rect 363656 53768 363662 53780
rect 366542 53768 366548 53780
rect 363656 53740 366548 53768
rect 363656 53728 363662 53740
rect 366542 53728 366548 53740
rect 366600 53728 366606 53780
rect 313918 53456 313924 53508
rect 313976 53496 313982 53508
rect 316770 53496 316776 53508
rect 313976 53468 316776 53496
rect 313976 53456 313982 53468
rect 316770 53456 316776 53468
rect 316828 53456 316834 53508
rect 363690 53252 363696 53304
rect 363748 53292 363754 53304
rect 367002 53292 367008 53304
rect 363748 53264 367008 53292
rect 363748 53252 363754 53264
rect 367002 53252 367008 53264
rect 367060 53252 367066 53304
rect 354030 53116 354036 53168
rect 354088 53156 354094 53168
rect 356238 53156 356244 53168
rect 354088 53128 356244 53156
rect 354088 53116 354094 53128
rect 356238 53116 356244 53128
rect 356296 53116 356302 53168
rect 264330 53048 264336 53100
rect 264388 53088 264394 53100
rect 281350 53088 281356 53100
rect 264388 53060 281356 53088
rect 264388 53048 264394 53060
rect 281350 53048 281356 53060
rect 281408 53048 281414 53100
rect 311158 53048 311164 53100
rect 311216 53088 311222 53100
rect 318150 53088 318156 53100
rect 311216 53060 318156 53088
rect 311216 53048 311222 53060
rect 318150 53048 318156 53060
rect 318208 53048 318214 53100
rect 333974 53048 333980 53100
rect 334032 53088 334038 53100
rect 340138 53088 340144 53100
rect 334032 53060 340144 53088
rect 334032 53048 334038 53060
rect 340138 53048 340144 53060
rect 340196 53048 340202 53100
rect 327902 52368 327908 52420
rect 327960 52408 327966 52420
rect 332594 52408 332600 52420
rect 327960 52380 332600 52408
rect 327960 52368 327966 52380
rect 332594 52368 332600 52380
rect 332652 52368 332658 52420
rect 362218 52368 362224 52420
rect 362276 52408 362282 52420
rect 365622 52408 365628 52420
rect 362276 52380 365628 52408
rect 362276 52368 362282 52380
rect 365622 52368 365628 52380
rect 365680 52368 365686 52420
rect 13814 51688 13820 51740
rect 13872 51728 13878 51740
rect 125042 51728 125048 51740
rect 13872 51700 125048 51728
rect 13872 51688 13878 51700
rect 125042 51688 125048 51700
rect 125100 51688 125106 51740
rect 295334 51688 295340 51740
rect 295392 51728 295398 51740
rect 318058 51728 318064 51740
rect 295392 51700 318064 51728
rect 295392 51688 295398 51700
rect 318058 51688 318064 51700
rect 318116 51688 318122 51740
rect 387702 51212 387708 51264
rect 387760 51252 387766 51264
rect 391198 51252 391204 51264
rect 387760 51224 391204 51252
rect 387760 51212 387766 51224
rect 391198 51212 391204 51224
rect 391256 51212 391262 51264
rect 253014 51008 253020 51060
rect 253072 51048 253078 51060
rect 258718 51048 258724 51060
rect 253072 51020 258724 51048
rect 253072 51008 253078 51020
rect 258718 51008 258724 51020
rect 258776 51008 258782 51060
rect 353938 51008 353944 51060
rect 353996 51048 354002 51060
rect 356698 51048 356704 51060
rect 353996 51020 356704 51048
rect 353996 51008 354002 51020
rect 356698 51008 356704 51020
rect 356756 51008 356762 51060
rect 269758 50940 269764 50992
rect 269816 50980 269822 50992
rect 273162 50980 273168 50992
rect 269816 50952 273168 50980
rect 269816 50940 269822 50952
rect 273162 50940 273168 50952
rect 273220 50940 273226 50992
rect 247678 50328 247684 50380
rect 247736 50368 247742 50380
rect 274726 50368 274732 50380
rect 247736 50340 274732 50368
rect 247736 50328 247742 50340
rect 274726 50328 274732 50340
rect 274784 50328 274790 50380
rect 331858 50328 331864 50380
rect 331916 50368 331922 50380
rect 339954 50368 339960 50380
rect 331916 50340 339960 50368
rect 331916 50328 331922 50340
rect 339954 50328 339960 50340
rect 340012 50328 340018 50380
rect 343634 50328 343640 50380
rect 343692 50368 343698 50380
rect 359458 50368 359464 50380
rect 343692 50340 359464 50368
rect 343692 50328 343698 50340
rect 359458 50328 359464 50340
rect 359516 50328 359522 50380
rect 366542 49784 366548 49836
rect 366600 49824 366606 49836
rect 373258 49824 373264 49836
rect 366600 49796 373264 49824
rect 366600 49784 366606 49796
rect 373258 49784 373264 49796
rect 373316 49784 373322 49836
rect 271138 49648 271144 49700
rect 271196 49688 271202 49700
rect 277486 49688 277492 49700
rect 271196 49660 277492 49688
rect 271196 49648 271202 49660
rect 277486 49648 277492 49660
rect 277544 49648 277550 49700
rect 307018 49648 307024 49700
rect 307076 49688 307082 49700
rect 311986 49688 311992 49700
rect 307076 49660 311992 49688
rect 307076 49648 307082 49660
rect 311986 49648 311992 49660
rect 312044 49648 312050 49700
rect 332594 49648 332600 49700
rect 332652 49688 332658 49700
rect 337378 49688 337384 49700
rect 332652 49660 337384 49688
rect 332652 49648 332658 49660
rect 337378 49648 337384 49660
rect 337436 49648 337442 49700
rect 349798 48220 349804 48272
rect 349856 48260 349862 48272
rect 352006 48260 352012 48272
rect 349856 48232 352012 48260
rect 349856 48220 349862 48232
rect 352006 48220 352012 48232
rect 352064 48220 352070 48272
rect 365622 48220 365628 48272
rect 365680 48260 365686 48272
rect 370498 48260 370504 48272
rect 365680 48232 370504 48260
rect 365680 48220 365686 48232
rect 370498 48220 370504 48232
rect 370556 48220 370562 48272
rect 367002 48152 367008 48204
rect 367060 48192 367066 48204
rect 371234 48192 371240 48204
rect 367060 48164 371240 48192
rect 367060 48152 367066 48164
rect 371234 48152 371240 48164
rect 371292 48152 371298 48204
rect 356238 47608 356244 47660
rect 356296 47648 356302 47660
rect 374178 47648 374184 47660
rect 356296 47620 374184 47648
rect 356296 47608 356302 47620
rect 374178 47608 374184 47620
rect 374236 47608 374242 47660
rect 163222 47540 163228 47592
rect 163280 47580 163286 47592
rect 488534 47580 488540 47592
rect 163280 47552 488540 47580
rect 163280 47540 163286 47552
rect 488534 47540 488540 47552
rect 488592 47540 488598 47592
rect 344278 47268 344284 47320
rect 344336 47308 344342 47320
rect 346394 47308 346400 47320
rect 344336 47280 346400 47308
rect 344336 47268 344342 47280
rect 346394 47268 346400 47280
rect 346452 47268 346458 47320
rect 118510 46860 118516 46912
rect 118568 46900 118574 46912
rect 580166 46900 580172 46912
rect 118568 46872 580172 46900
rect 118568 46860 118574 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 264238 46792 264244 46844
rect 264296 46832 264302 46844
rect 266998 46832 267004 46844
rect 264296 46804 267004 46832
rect 264296 46792 264302 46804
rect 266998 46792 267004 46804
rect 267056 46792 267062 46844
rect 301590 46792 301596 46844
rect 301648 46832 301654 46844
rect 304258 46832 304264 46844
rect 301648 46804 304264 46832
rect 301648 46792 301654 46804
rect 304258 46792 304264 46804
rect 304316 46792 304322 46844
rect 274726 46520 274732 46572
rect 274784 46560 274790 46572
rect 279418 46560 279424 46572
rect 274784 46532 279424 46560
rect 274784 46520 274790 46532
rect 279418 46520 279424 46532
rect 279476 46520 279482 46572
rect 273162 46248 273168 46300
rect 273220 46288 273226 46300
rect 282178 46288 282184 46300
rect 273220 46260 282184 46288
rect 273220 46248 273226 46260
rect 282178 46248 282184 46260
rect 282236 46248 282242 46300
rect 277486 46180 277492 46232
rect 277544 46220 277550 46232
rect 288434 46220 288440 46232
rect 277544 46192 288440 46220
rect 277544 46180 277550 46192
rect 288434 46180 288440 46192
rect 288492 46180 288498 46232
rect 292666 46180 292672 46232
rect 292724 46220 292730 46232
rect 301498 46220 301504 46232
rect 292724 46192 301504 46220
rect 292724 46180 292730 46192
rect 301498 46180 301504 46192
rect 301556 46180 301562 46232
rect 339954 46180 339960 46232
rect 340012 46220 340018 46232
rect 349798 46220 349804 46232
rect 340012 46192 349804 46220
rect 340012 46180 340018 46192
rect 349798 46180 349804 46192
rect 349856 46180 349862 46232
rect 311986 46044 311992 46096
rect 312044 46084 312050 46096
rect 317414 46084 317420 46096
rect 312044 46056 317420 46084
rect 312044 46044 312050 46056
rect 317414 46044 317420 46056
rect 317472 46044 317478 46096
rect 281350 45568 281356 45620
rect 281408 45608 281414 45620
rect 287698 45608 287704 45620
rect 281408 45580 287704 45608
rect 281408 45568 281414 45580
rect 287698 45568 287704 45580
rect 287756 45568 287762 45620
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 174078 45540 174084 45552
rect 3476 45512 174084 45540
rect 3476 45500 3482 45512
rect 174078 45500 174084 45512
rect 174136 45500 174142 45552
rect 327718 45092 327724 45144
rect 327776 45132 327782 45144
rect 332594 45132 332600 45144
rect 327776 45104 332600 45132
rect 327776 45092 327782 45104
rect 332594 45092 332600 45104
rect 332652 45092 332658 45144
rect 346394 44888 346400 44940
rect 346452 44928 346458 44940
rect 359550 44928 359556 44940
rect 346452 44900 359556 44928
rect 346452 44888 346458 44900
rect 359550 44888 359556 44900
rect 359608 44888 359614 44940
rect 67634 44820 67640 44872
rect 67692 44860 67698 44872
rect 130194 44860 130200 44872
rect 67692 44832 130200 44860
rect 67692 44820 67698 44832
rect 130194 44820 130200 44832
rect 130252 44820 130258 44872
rect 139762 44820 139768 44872
rect 139820 44860 139826 44872
rect 185026 44860 185032 44872
rect 139820 44832 185032 44860
rect 139820 44820 139826 44832
rect 185026 44820 185032 44832
rect 185084 44820 185090 44872
rect 340138 44820 340144 44872
rect 340196 44860 340202 44872
rect 352098 44860 352104 44872
rect 340196 44832 352104 44860
rect 340196 44820 340202 44832
rect 352098 44820 352104 44832
rect 352156 44820 352162 44872
rect 318150 44684 318156 44736
rect 318208 44724 318214 44736
rect 324314 44724 324320 44736
rect 318208 44696 324320 44724
rect 318208 44684 318214 44696
rect 324314 44684 324320 44696
rect 324372 44684 324378 44736
rect 374178 44616 374184 44668
rect 374236 44656 374242 44668
rect 383010 44656 383016 44668
rect 374236 44628 383016 44656
rect 374236 44616 374242 44628
rect 383010 44616 383016 44628
rect 383068 44616 383074 44668
rect 335998 44140 336004 44192
rect 336056 44180 336062 44192
rect 339402 44180 339408 44192
rect 336056 44152 339408 44180
rect 336056 44140 336062 44152
rect 339402 44140 339408 44152
rect 339460 44140 339466 44192
rect 317414 43392 317420 43444
rect 317472 43432 317478 43444
rect 344278 43432 344284 43444
rect 317472 43404 344284 43432
rect 317472 43392 317478 43404
rect 344278 43392 344284 43404
rect 344336 43392 344342 43444
rect 371234 43120 371240 43172
rect 371292 43160 371298 43172
rect 376018 43160 376024 43172
rect 371292 43132 376024 43160
rect 371292 43120 371298 43132
rect 376018 43120 376024 43132
rect 376076 43120 376082 43172
rect 269850 42916 269856 42968
rect 269908 42956 269914 42968
rect 276014 42956 276020 42968
rect 269908 42928 276020 42956
rect 269908 42916 269914 42928
rect 276014 42916 276020 42928
rect 276072 42916 276078 42968
rect 316770 42780 316776 42832
rect 316828 42820 316834 42832
rect 319438 42820 319444 42832
rect 316828 42792 319444 42820
rect 316828 42780 316834 42792
rect 319438 42780 319444 42792
rect 319496 42780 319502 42832
rect 352006 42712 352012 42764
rect 352064 42752 352070 42764
rect 355318 42752 355324 42764
rect 352064 42724 355324 42752
rect 352064 42712 352070 42724
rect 355318 42712 355324 42724
rect 355376 42712 355382 42764
rect 280798 42236 280804 42288
rect 280856 42276 280862 42288
rect 284294 42276 284300 42288
rect 280856 42248 284300 42276
rect 280856 42236 280862 42248
rect 284294 42236 284300 42248
rect 284352 42236 284358 42288
rect 316678 41828 316684 41880
rect 316736 41868 316742 41880
rect 319806 41868 319812 41880
rect 316736 41840 319812 41868
rect 316736 41828 316742 41840
rect 319806 41828 319812 41840
rect 319864 41828 319870 41880
rect 324314 40672 324320 40724
rect 324372 40712 324378 40724
rect 330478 40712 330484 40724
rect 324372 40684 330484 40712
rect 324372 40672 324378 40684
rect 330478 40672 330484 40684
rect 330536 40672 330542 40724
rect 339402 40672 339408 40724
rect 339460 40712 339466 40724
rect 341058 40712 341064 40724
rect 339460 40684 341064 40712
rect 339460 40672 339466 40684
rect 341058 40672 341064 40684
rect 341116 40672 341122 40724
rect 352098 40672 352104 40724
rect 352156 40712 352162 40724
rect 375282 40712 375288 40724
rect 352156 40684 375288 40712
rect 352156 40672 352162 40684
rect 375282 40672 375288 40684
rect 375340 40672 375346 40724
rect 288434 39992 288440 40044
rect 288492 40032 288498 40044
rect 291838 40032 291844 40044
rect 288492 40004 291844 40032
rect 288492 39992 288498 40004
rect 291838 39992 291844 40004
rect 291896 39992 291902 40044
rect 323578 39992 323584 40044
rect 323636 40032 323642 40044
rect 326430 40032 326436 40044
rect 323636 40004 326436 40032
rect 323636 39992 323642 40004
rect 326430 39992 326436 40004
rect 326488 39992 326494 40044
rect 276014 39380 276020 39432
rect 276072 39420 276078 39432
rect 284938 39420 284944 39432
rect 276072 39392 284944 39420
rect 276072 39380 276078 39392
rect 284938 39380 284944 39392
rect 284996 39380 285002 39432
rect 332594 39380 332600 39432
rect 332652 39420 332658 39432
rect 340138 39420 340144 39432
rect 332652 39392 340144 39420
rect 332652 39380 332658 39392
rect 340138 39380 340144 39392
rect 340196 39380 340202 39432
rect 258718 39312 258724 39364
rect 258776 39352 258782 39364
rect 278038 39352 278044 39364
rect 258776 39324 278044 39352
rect 258776 39312 258782 39324
rect 278038 39312 278044 39324
rect 278096 39312 278102 39364
rect 326338 39312 326344 39364
rect 326396 39352 326402 39364
rect 337930 39352 337936 39364
rect 326396 39324 337936 39352
rect 326396 39312 326402 39324
rect 337930 39312 337936 39324
rect 337988 39312 337994 39364
rect 345658 39312 345664 39364
rect 345716 39352 345722 39364
rect 362218 39352 362224 39364
rect 345716 39324 362224 39352
rect 345716 39312 345722 39324
rect 362218 39312 362224 39324
rect 362276 39312 362282 39364
rect 45554 37884 45560 37936
rect 45612 37924 45618 37936
rect 116578 37924 116584 37936
rect 45612 37896 116584 37924
rect 45612 37884 45618 37896
rect 116578 37884 116584 37896
rect 116636 37884 116642 37936
rect 282178 37884 282184 37936
rect 282236 37924 282242 37936
rect 298278 37924 298284 37936
rect 282236 37896 298284 37924
rect 282236 37884 282242 37896
rect 298278 37884 298284 37896
rect 298336 37884 298342 37936
rect 375282 37884 375288 37936
rect 375340 37924 375346 37936
rect 388438 37924 388444 37936
rect 375340 37896 388444 37924
rect 375340 37884 375346 37896
rect 388438 37884 388444 37896
rect 388496 37884 388502 37936
rect 284294 37476 284300 37528
rect 284352 37516 284358 37528
rect 287422 37516 287428 37528
rect 284352 37488 287428 37516
rect 284352 37476 284358 37488
rect 287422 37476 287428 37488
rect 287480 37476 287486 37528
rect 380158 37272 380164 37324
rect 380216 37312 380222 37324
rect 384298 37312 384304 37324
rect 380216 37284 384304 37312
rect 380216 37272 380222 37284
rect 384298 37272 384304 37284
rect 384356 37272 384362 37324
rect 319806 37204 319812 37256
rect 319864 37244 319870 37256
rect 322842 37244 322848 37256
rect 319864 37216 322848 37244
rect 319864 37204 319870 37216
rect 322842 37204 322848 37216
rect 322900 37204 322906 37256
rect 337930 37204 337936 37256
rect 337988 37244 337994 37256
rect 342898 37244 342904 37256
rect 337988 37216 342904 37244
rect 337988 37204 337994 37216
rect 342898 37204 342904 37216
rect 342956 37204 342962 37256
rect 355318 37204 355324 37256
rect 355376 37244 355382 37256
rect 360838 37244 360844 37256
rect 355376 37216 360844 37244
rect 355376 37204 355382 37216
rect 360838 37204 360844 37216
rect 360896 37204 360902 37256
rect 341058 37136 341064 37188
rect 341116 37176 341122 37188
rect 344370 37176 344376 37188
rect 341116 37148 344376 37176
rect 341116 37136 341122 37148
rect 344370 37136 344376 37148
rect 344428 37136 344434 37188
rect 340138 36592 340144 36644
rect 340196 36632 340202 36644
rect 362126 36632 362132 36644
rect 340196 36604 362132 36632
rect 340196 36592 340202 36604
rect 362126 36592 362132 36604
rect 362184 36592 362190 36644
rect 7558 36524 7564 36576
rect 7616 36564 7622 36576
rect 124214 36564 124220 36576
rect 7616 36536 124220 36564
rect 7616 36524 7622 36536
rect 124214 36524 124220 36536
rect 124272 36524 124278 36576
rect 172146 36524 172152 36576
rect 172204 36564 172210 36576
rect 418154 36564 418160 36576
rect 172204 36536 418160 36564
rect 172204 36524 172210 36536
rect 418154 36524 418160 36536
rect 418212 36524 418218 36576
rect 382918 35912 382924 35964
rect 382976 35952 382982 35964
rect 385678 35952 385684 35964
rect 382976 35924 385684 35952
rect 382976 35912 382982 35924
rect 385678 35912 385684 35924
rect 385736 35912 385742 35964
rect 148134 35300 148140 35352
rect 148192 35340 148198 35352
rect 287054 35340 287060 35352
rect 148192 35312 287060 35340
rect 148192 35300 148198 35312
rect 287054 35300 287060 35312
rect 287112 35300 287118 35352
rect 287422 35300 287428 35352
rect 287480 35340 287486 35352
rect 299198 35340 299204 35352
rect 287480 35312 299204 35340
rect 287480 35300 287486 35312
rect 299198 35300 299204 35312
rect 299256 35300 299262 35352
rect 356698 35300 356704 35352
rect 356756 35340 356762 35352
rect 361574 35340 361580 35352
rect 356756 35312 361580 35340
rect 356756 35300 356762 35312
rect 361574 35300 361580 35312
rect 361632 35300 361638 35352
rect 148226 35232 148232 35284
rect 148284 35272 148290 35284
rect 291194 35272 291200 35284
rect 148284 35244 291200 35272
rect 148284 35232 148290 35244
rect 291194 35232 291200 35244
rect 291252 35232 291258 35284
rect 38654 35164 38660 35216
rect 38712 35204 38718 35216
rect 122190 35204 122196 35216
rect 38712 35176 122196 35204
rect 38712 35164 38718 35176
rect 122190 35164 122196 35176
rect 122248 35164 122254 35216
rect 153562 35164 153568 35216
rect 153620 35204 153626 35216
rect 357434 35204 357440 35216
rect 153620 35176 357440 35204
rect 153620 35164 153626 35176
rect 357434 35164 357440 35176
rect 357492 35164 357498 35216
rect 278038 34552 278044 34604
rect 278096 34592 278102 34604
rect 285674 34592 285680 34604
rect 278096 34564 285680 34592
rect 278096 34552 278102 34564
rect 285674 34552 285680 34564
rect 285732 34552 285738 34604
rect 141326 33940 141332 33992
rect 141384 33980 141390 33992
rect 198734 33980 198740 33992
rect 141384 33952 198740 33980
rect 141384 33940 141390 33952
rect 198734 33940 198740 33952
rect 198792 33940 198798 33992
rect 344278 33940 344284 33992
rect 344336 33980 344342 33992
rect 347590 33980 347596 33992
rect 344336 33952 347596 33980
rect 344336 33940 344342 33952
rect 347590 33940 347596 33952
rect 347648 33940 347654 33992
rect 141234 33872 141240 33924
rect 141292 33912 141298 33924
rect 205634 33912 205640 33924
rect 141292 33884 205640 33912
rect 141292 33872 141298 33884
rect 205634 33872 205640 33884
rect 205692 33872 205698 33924
rect 142522 33804 142528 33856
rect 142580 33844 142586 33856
rect 219434 33844 219440 33856
rect 142580 33816 219440 33844
rect 142580 33804 142586 33816
rect 219434 33804 219440 33816
rect 219492 33804 219498 33856
rect 376018 33804 376024 33856
rect 376076 33844 376082 33856
rect 384482 33844 384488 33856
rect 376076 33816 384488 33844
rect 376076 33804 376082 33816
rect 384482 33804 384488 33816
rect 384540 33804 384546 33856
rect 145466 33736 145472 33788
rect 145524 33776 145530 33788
rect 259454 33776 259460 33788
rect 145524 33748 259460 33776
rect 145524 33736 145530 33748
rect 259454 33736 259460 33748
rect 259512 33736 259518 33788
rect 322842 33736 322848 33788
rect 322900 33776 322906 33788
rect 329098 33776 329104 33788
rect 322900 33748 329104 33776
rect 322900 33736 322906 33748
rect 329098 33736 329104 33748
rect 329156 33736 329162 33788
rect 383010 33736 383016 33788
rect 383068 33776 383074 33788
rect 396718 33776 396724 33788
rect 383068 33748 396724 33776
rect 383068 33736 383074 33748
rect 396718 33736 396724 33748
rect 396776 33736 396782 33788
rect 171962 33056 171968 33108
rect 172020 33096 172026 33108
rect 580166 33096 580172 33108
rect 172020 33068 580172 33096
rect 172020 33056 172026 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 361574 32988 361580 33040
rect 361632 33028 361638 33040
rect 364978 33028 364984 33040
rect 361632 33000 364984 33028
rect 361632 32988 361638 33000
rect 364978 32988 364984 33000
rect 365036 32988 365042 33040
rect 384390 32784 384396 32836
rect 384448 32824 384454 32836
rect 391934 32824 391940 32836
rect 384448 32796 391940 32824
rect 384448 32784 384454 32796
rect 391934 32784 391940 32796
rect 391992 32784 391998 32836
rect 139670 32716 139676 32768
rect 139728 32756 139734 32768
rect 187694 32756 187700 32768
rect 139728 32728 187700 32756
rect 139728 32716 139734 32728
rect 187694 32716 187700 32728
rect 187752 32716 187758 32768
rect 370498 32716 370504 32768
rect 370556 32756 370562 32768
rect 378134 32756 378140 32768
rect 370556 32728 378140 32756
rect 370556 32716 370562 32728
rect 378134 32716 378140 32728
rect 378192 32716 378198 32768
rect 141142 32648 141148 32700
rect 141200 32688 141206 32700
rect 201494 32688 201500 32700
rect 141200 32660 201500 32688
rect 141200 32648 141206 32660
rect 201494 32648 201500 32660
rect 201552 32648 201558 32700
rect 266998 32648 267004 32700
rect 267056 32688 267062 32700
rect 275278 32688 275284 32700
rect 267056 32660 275284 32688
rect 267056 32648 267062 32660
rect 275278 32648 275284 32660
rect 275336 32648 275342 32700
rect 285674 32648 285680 32700
rect 285732 32688 285738 32700
rect 293954 32688 293960 32700
rect 285732 32660 293960 32688
rect 285732 32648 285738 32660
rect 293954 32648 293960 32660
rect 294012 32648 294018 32700
rect 362126 32648 362132 32700
rect 362184 32688 362190 32700
rect 374730 32688 374736 32700
rect 362184 32660 374736 32688
rect 362184 32648 362190 32660
rect 374730 32648 374736 32660
rect 374788 32648 374794 32700
rect 160830 32580 160836 32632
rect 160888 32620 160894 32632
rect 447134 32620 447140 32632
rect 160888 32592 447140 32620
rect 160888 32580 160894 32592
rect 447134 32580 447140 32592
rect 447192 32580 447198 32632
rect 3418 32512 3424 32564
rect 3476 32552 3482 32564
rect 7650 32552 7656 32564
rect 3476 32524 7656 32552
rect 3476 32512 3482 32524
rect 7650 32512 7656 32524
rect 7708 32512 7714 32564
rect 166166 32512 166172 32564
rect 166224 32552 166230 32564
rect 473998 32552 474004 32564
rect 166224 32524 474004 32552
rect 166224 32512 166230 32524
rect 473998 32512 474004 32524
rect 474056 32512 474062 32564
rect 163130 32444 163136 32496
rect 163188 32484 163194 32496
rect 485774 32484 485780 32496
rect 163188 32456 485780 32484
rect 163188 32444 163194 32456
rect 485774 32444 485780 32456
rect 485832 32444 485838 32496
rect 31754 32376 31760 32428
rect 31812 32416 31818 32428
rect 120718 32416 120724 32428
rect 31812 32388 120724 32416
rect 31812 32376 31818 32388
rect 120718 32376 120724 32388
rect 120776 32376 120782 32428
rect 164694 32376 164700 32428
rect 164752 32416 164758 32428
rect 503714 32416 503720 32428
rect 164752 32388 503720 32416
rect 164752 32376 164758 32388
rect 503714 32376 503720 32388
rect 503772 32376 503778 32428
rect 374638 31764 374644 31816
rect 374696 31804 374702 31816
rect 377398 31804 377404 31816
rect 374696 31776 377404 31804
rect 374696 31764 374702 31776
rect 377398 31764 377404 31776
rect 377456 31764 377462 31816
rect 349798 31696 349804 31748
rect 349856 31736 349862 31748
rect 353386 31736 353392 31748
rect 349856 31708 353392 31736
rect 349856 31696 349862 31708
rect 353386 31696 353392 31708
rect 353444 31696 353450 31748
rect 318058 31492 318064 31544
rect 318116 31532 318122 31544
rect 322934 31532 322940 31544
rect 318116 31504 322940 31532
rect 318116 31492 318122 31504
rect 322934 31492 322940 31504
rect 322992 31492 322998 31544
rect 326430 31220 326436 31272
rect 326488 31260 326494 31272
rect 331214 31260 331220 31272
rect 326488 31232 331220 31260
rect 326488 31220 326494 31232
rect 331214 31220 331220 31232
rect 331272 31220 331278 31272
rect 291838 31152 291844 31204
rect 291896 31192 291902 31204
rect 301590 31192 301596 31204
rect 291896 31164 301596 31192
rect 291896 31152 291902 31164
rect 301590 31152 301596 31164
rect 301648 31152 301654 31204
rect 337378 31152 337384 31204
rect 337436 31192 337442 31204
rect 347038 31192 347044 31204
rect 337436 31164 347044 31192
rect 337436 31152 337442 31164
rect 347038 31152 347044 31164
rect 347096 31152 347102 31204
rect 299198 31084 299204 31136
rect 299256 31124 299262 31136
rect 313274 31124 313280 31136
rect 299256 31096 313280 31124
rect 299256 31084 299262 31096
rect 313274 31084 313280 31096
rect 313332 31084 313338 31136
rect 342898 31084 342904 31136
rect 342956 31124 342962 31136
rect 353478 31124 353484 31136
rect 342956 31096 353484 31124
rect 342956 31084 342962 31096
rect 353478 31084 353484 31096
rect 353536 31084 353542 31136
rect 371878 31084 371884 31136
rect 371936 31124 371942 31136
rect 378778 31124 378784 31136
rect 371936 31096 378784 31124
rect 371936 31084 371942 31096
rect 378778 31084 378784 31096
rect 378836 31084 378842 31136
rect 164602 31016 164608 31068
rect 164660 31056 164666 31068
rect 499574 31056 499580 31068
rect 164660 31028 499580 31056
rect 164660 31016 164666 31028
rect 499574 31016 499580 31028
rect 499632 31016 499638 31068
rect 279418 30268 279424 30320
rect 279476 30308 279482 30320
rect 286318 30308 286324 30320
rect 279476 30280 286324 30308
rect 279476 30268 279482 30280
rect 286318 30268 286324 30280
rect 286376 30268 286382 30320
rect 387058 30268 387064 30320
rect 387116 30308 387122 30320
rect 392578 30308 392584 30320
rect 387116 30280 392584 30308
rect 387116 30268 387122 30280
rect 392578 30268 392584 30280
rect 392636 30268 392642 30320
rect 298278 29996 298284 30048
rect 298336 30036 298342 30048
rect 311158 30036 311164 30048
rect 298336 30008 311164 30036
rect 298336 29996 298342 30008
rect 311158 29996 311164 30008
rect 311216 29996 311222 30048
rect 293954 29928 293960 29980
rect 294012 29968 294018 29980
rect 320818 29968 320824 29980
rect 294012 29940 320824 29968
rect 294012 29928 294018 29940
rect 320818 29928 320824 29940
rect 320876 29928 320882 29980
rect 148042 29860 148048 29912
rect 148100 29900 148106 29912
rect 285674 29900 285680 29912
rect 148100 29872 285680 29900
rect 148100 29860 148106 29872
rect 285674 29860 285680 29872
rect 285732 29860 285738 29912
rect 298738 29860 298744 29912
rect 298796 29900 298802 29912
rect 326430 29900 326436 29912
rect 298796 29872 326436 29900
rect 298796 29860 298802 29872
rect 326430 29860 326436 29872
rect 326488 29860 326494 29912
rect 154114 29792 154120 29844
rect 154172 29832 154178 29844
rect 332594 29832 332600 29844
rect 154172 29804 332600 29832
rect 154172 29792 154178 29804
rect 332594 29792 332600 29804
rect 332652 29792 332658 29844
rect 152366 29724 152372 29776
rect 152424 29764 152430 29776
rect 339494 29764 339500 29776
rect 152424 29736 339500 29764
rect 152424 29724 152430 29736
rect 339494 29724 339500 29736
rect 339552 29724 339558 29776
rect 152274 29656 152280 29708
rect 152332 29696 152338 29708
rect 346394 29696 346400 29708
rect 152332 29668 346400 29696
rect 152332 29656 152338 29668
rect 346394 29656 346400 29668
rect 346452 29656 346458 29708
rect 391934 29656 391940 29708
rect 391992 29696 391998 29708
rect 397546 29696 397552 29708
rect 391992 29668 397552 29696
rect 391992 29656 391998 29668
rect 397546 29656 397552 29668
rect 397604 29656 397610 29708
rect 157794 29588 157800 29640
rect 157852 29628 157858 29640
rect 409874 29628 409880 29640
rect 157852 29600 409880 29628
rect 157852 29588 157858 29600
rect 409874 29588 409880 29600
rect 409932 29588 409938 29640
rect 287698 28908 287704 28960
rect 287756 28948 287762 28960
rect 291102 28948 291108 28960
rect 287756 28920 291108 28948
rect 287756 28908 287762 28920
rect 291102 28908 291108 28920
rect 291160 28908 291166 28960
rect 378134 28908 378140 28960
rect 378192 28948 378198 28960
rect 381538 28948 381544 28960
rect 378192 28920 381544 28948
rect 378192 28908 378198 28920
rect 381538 28908 381544 28920
rect 381596 28908 381602 28960
rect 360838 28772 360844 28824
rect 360896 28812 360902 28824
rect 365162 28812 365168 28824
rect 360896 28784 365168 28812
rect 360896 28772 360902 28784
rect 365162 28772 365168 28784
rect 365220 28772 365226 28824
rect 143994 28568 144000 28620
rect 144052 28608 144058 28620
rect 242894 28608 242900 28620
rect 144052 28580 242900 28608
rect 144052 28568 144058 28580
rect 242894 28568 242900 28580
rect 242952 28568 242958 28620
rect 145282 28500 145288 28552
rect 145340 28540 145346 28552
rect 251266 28540 251272 28552
rect 145340 28512 251272 28540
rect 145340 28500 145346 28512
rect 251266 28500 251272 28512
rect 251324 28500 251330 28552
rect 145190 28432 145196 28484
rect 145248 28472 145254 28484
rect 253934 28472 253940 28484
rect 145248 28444 253940 28472
rect 145248 28432 145254 28444
rect 253934 28432 253940 28444
rect 253992 28432 253998 28484
rect 344370 28432 344376 28484
rect 344428 28472 344434 28484
rect 348878 28472 348884 28484
rect 344428 28444 348884 28472
rect 344428 28432 344434 28444
rect 348878 28432 348884 28444
rect 348936 28432 348942 28484
rect 145374 28364 145380 28416
rect 145432 28404 145438 28416
rect 258074 28404 258080 28416
rect 145432 28376 258080 28404
rect 145432 28364 145438 28376
rect 258074 28364 258080 28376
rect 258132 28364 258138 28416
rect 304258 28364 304264 28416
rect 304316 28404 304322 28416
rect 323486 28404 323492 28416
rect 304316 28376 323492 28404
rect 304316 28364 304322 28376
rect 323486 28364 323492 28376
rect 323544 28364 323550 28416
rect 347590 28364 347596 28416
rect 347648 28404 347654 28416
rect 356698 28404 356704 28416
rect 347648 28376 356704 28404
rect 347648 28364 347654 28376
rect 356698 28364 356704 28376
rect 356756 28364 356762 28416
rect 171778 28296 171784 28348
rect 171836 28336 171842 28348
rect 397454 28336 397460 28348
rect 171836 28308 397460 28336
rect 171836 28296 171842 28308
rect 397454 28296 397460 28308
rect 397512 28296 397518 28348
rect 167638 28228 167644 28280
rect 167696 28268 167702 28280
rect 539686 28268 539692 28280
rect 167696 28240 539692 28268
rect 167696 28228 167702 28240
rect 539686 28228 539692 28240
rect 539744 28228 539750 28280
rect 353386 27684 353392 27736
rect 353444 27724 353450 27736
rect 356054 27724 356060 27736
rect 353444 27696 356060 27724
rect 353444 27684 353450 27696
rect 356054 27684 356060 27696
rect 356112 27684 356118 27736
rect 378778 27684 378784 27736
rect 378836 27724 378842 27736
rect 385034 27724 385040 27736
rect 378836 27696 385040 27724
rect 378836 27684 378842 27696
rect 385034 27684 385040 27696
rect 385092 27684 385098 27736
rect 330478 27548 330484 27600
rect 330536 27588 330542 27600
rect 334250 27588 334256 27600
rect 330536 27560 334256 27588
rect 330536 27548 330542 27560
rect 334250 27548 334256 27560
rect 334308 27548 334314 27600
rect 359550 27548 359556 27600
rect 359608 27588 359614 27600
rect 363322 27588 363328 27600
rect 359608 27560 363328 27588
rect 359608 27548 359614 27560
rect 363322 27548 363328 27560
rect 363380 27548 363386 27600
rect 397546 27548 397552 27600
rect 397604 27588 397610 27600
rect 400858 27588 400864 27600
rect 397604 27560 400864 27588
rect 397604 27548 397610 27560
rect 400858 27548 400864 27560
rect 400916 27548 400922 27600
rect 140958 27344 140964 27396
rect 141016 27384 141022 27396
rect 204254 27384 204260 27396
rect 141016 27356 204260 27384
rect 141016 27344 141022 27356
rect 204254 27344 204260 27356
rect 204312 27344 204318 27396
rect 141050 27276 141056 27328
rect 141108 27316 141114 27328
rect 208394 27316 208400 27328
rect 141108 27288 208400 27316
rect 141108 27276 141114 27288
rect 208394 27276 208400 27288
rect 208452 27276 208458 27328
rect 142430 27208 142436 27260
rect 142488 27248 142494 27260
rect 215294 27248 215300 27260
rect 142488 27220 215300 27248
rect 142488 27208 142494 27220
rect 215294 27208 215300 27220
rect 215352 27208 215358 27260
rect 142338 27140 142344 27192
rect 142396 27180 142402 27192
rect 218146 27180 218152 27192
rect 142396 27152 218152 27180
rect 142396 27140 142402 27152
rect 218146 27140 218152 27152
rect 218204 27140 218210 27192
rect 143902 27072 143908 27124
rect 143960 27112 143966 27124
rect 235994 27112 236000 27124
rect 143960 27084 236000 27112
rect 143960 27072 143966 27084
rect 235994 27072 236000 27084
rect 236052 27072 236058 27124
rect 295978 27072 295984 27124
rect 296036 27112 296042 27124
rect 302878 27112 302884 27124
rect 296036 27084 302884 27112
rect 296036 27072 296042 27084
rect 302878 27072 302884 27084
rect 302936 27072 302942 27124
rect 149514 27004 149520 27056
rect 149572 27044 149578 27056
rect 303614 27044 303620 27056
rect 149572 27016 303620 27044
rect 149572 27004 149578 27016
rect 303614 27004 303620 27016
rect 303672 27004 303678 27056
rect 313274 27004 313280 27056
rect 313332 27044 313338 27056
rect 321738 27044 321744 27056
rect 313332 27016 321744 27044
rect 313332 27004 313338 27016
rect 321738 27004 321744 27016
rect 321796 27004 321802 27056
rect 171686 26936 171692 26988
rect 171744 26976 171750 26988
rect 411254 26976 411260 26988
rect 171744 26948 411260 26976
rect 171744 26936 171750 26948
rect 411254 26936 411260 26948
rect 411312 26936 411318 26988
rect 168926 26868 168932 26920
rect 168984 26908 168990 26920
rect 560294 26908 560300 26920
rect 168984 26880 560300 26908
rect 168984 26868 168990 26880
rect 560294 26868 560300 26880
rect 560352 26868 560358 26920
rect 331214 26460 331220 26512
rect 331272 26500 331278 26512
rect 335354 26500 335360 26512
rect 331272 26472 335360 26500
rect 331272 26460 331278 26472
rect 335354 26460 335360 26472
rect 335412 26460 335418 26512
rect 353478 26256 353484 26308
rect 353536 26296 353542 26308
rect 356146 26296 356152 26308
rect 353536 26268 356152 26296
rect 353536 26256 353542 26268
rect 356146 26256 356152 26268
rect 356204 26256 356210 26308
rect 140406 25984 140412 26036
rect 140464 26024 140470 26036
rect 176746 26024 176752 26036
rect 140464 25996 176752 26024
rect 140464 25984 140470 25996
rect 176746 25984 176752 25996
rect 176804 25984 176810 26036
rect 139486 25916 139492 25968
rect 139544 25956 139550 25968
rect 179414 25956 179420 25968
rect 139544 25928 179420 25956
rect 139544 25916 139550 25928
rect 179414 25916 179420 25928
rect 179472 25916 179478 25968
rect 139578 25848 139584 25900
rect 139636 25888 139642 25900
rect 183554 25888 183560 25900
rect 139636 25860 183560 25888
rect 139636 25848 139642 25860
rect 183554 25848 183560 25860
rect 183612 25848 183618 25900
rect 139394 25780 139400 25832
rect 139452 25820 139458 25832
rect 186314 25820 186320 25832
rect 139452 25792 186320 25820
rect 139452 25780 139458 25792
rect 186314 25780 186320 25792
rect 186372 25780 186378 25832
rect 140866 25712 140872 25764
rect 140924 25752 140930 25764
rect 201586 25752 201592 25764
rect 140924 25724 201592 25752
rect 140924 25712 140930 25724
rect 201586 25712 201592 25724
rect 201644 25712 201650 25764
rect 291102 25712 291108 25764
rect 291160 25752 291166 25764
rect 302234 25752 302240 25764
rect 291160 25724 302240 25752
rect 291160 25712 291166 25724
rect 302234 25712 302240 25724
rect 302292 25712 302298 25764
rect 147950 25644 147956 25696
rect 148008 25684 148014 25696
rect 292666 25684 292672 25696
rect 148008 25656 292672 25684
rect 148008 25644 148014 25656
rect 292666 25644 292672 25656
rect 292724 25644 292730 25696
rect 374730 25644 374736 25696
rect 374788 25684 374794 25696
rect 381630 25684 381636 25696
rect 374788 25656 381636 25684
rect 374788 25644 374794 25656
rect 381630 25644 381636 25656
rect 381688 25644 381694 25696
rect 157702 25576 157708 25628
rect 157760 25616 157766 25628
rect 414014 25616 414020 25628
rect 157760 25588 414020 25616
rect 157760 25576 157766 25588
rect 414014 25576 414020 25588
rect 414072 25576 414078 25628
rect 167546 25508 167552 25560
rect 167604 25548 167610 25560
rect 535454 25548 535460 25560
rect 167604 25520 535460 25548
rect 167604 25508 167610 25520
rect 535454 25508 535460 25520
rect 535512 25508 535518 25560
rect 348878 25236 348884 25288
rect 348936 25276 348942 25288
rect 351822 25276 351828 25288
rect 348936 25248 351828 25276
rect 348936 25236 348942 25248
rect 351822 25236 351828 25248
rect 351880 25236 351886 25288
rect 301498 24828 301504 24880
rect 301556 24868 301562 24880
rect 305638 24868 305644 24880
rect 301556 24840 305644 24868
rect 301556 24828 301562 24840
rect 305638 24828 305644 24840
rect 305696 24828 305702 24880
rect 377398 24828 377404 24880
rect 377456 24868 377462 24880
rect 380158 24868 380164 24880
rect 377456 24840 380164 24868
rect 377456 24828 377462 24840
rect 380158 24828 380164 24840
rect 380216 24828 380222 24880
rect 286318 24692 286324 24744
rect 286376 24732 286382 24744
rect 292758 24732 292764 24744
rect 286376 24704 292764 24732
rect 286376 24692 286382 24704
rect 292758 24692 292764 24704
rect 292816 24692 292822 24744
rect 363322 24692 363328 24744
rect 363380 24732 363386 24744
rect 369118 24732 369124 24744
rect 363380 24704 369124 24732
rect 363380 24692 363386 24704
rect 369118 24692 369124 24704
rect 369176 24692 369182 24744
rect 147858 24624 147864 24676
rect 147916 24664 147922 24676
rect 289814 24664 289820 24676
rect 147916 24636 289820 24664
rect 147916 24624 147922 24636
rect 289814 24624 289820 24636
rect 289872 24624 289878 24676
rect 334250 24624 334256 24676
rect 334308 24664 334314 24676
rect 342254 24664 342260 24676
rect 334308 24636 342260 24664
rect 334308 24624 334314 24636
rect 342254 24624 342260 24636
rect 342312 24624 342318 24676
rect 356054 24624 356060 24676
rect 356112 24664 356118 24676
rect 369854 24664 369860 24676
rect 356112 24636 369860 24664
rect 356112 24624 356118 24636
rect 369854 24624 369860 24636
rect 369912 24624 369918 24676
rect 384482 24624 384488 24676
rect 384540 24664 384546 24676
rect 407206 24664 407212 24676
rect 384540 24636 407212 24664
rect 384540 24624 384546 24636
rect 407206 24624 407212 24636
rect 407264 24624 407270 24676
rect 157610 24556 157616 24608
rect 157668 24596 157674 24608
rect 416774 24596 416780 24608
rect 157668 24568 416780 24596
rect 157668 24556 157674 24568
rect 416774 24556 416780 24568
rect 416832 24556 416838 24608
rect 168742 24488 168748 24540
rect 168800 24528 168806 24540
rect 552014 24528 552020 24540
rect 168800 24500 552020 24528
rect 168800 24488 168806 24500
rect 552014 24488 552020 24500
rect 552072 24488 552078 24540
rect 169662 24420 169668 24472
rect 169720 24460 169726 24472
rect 556154 24460 556160 24472
rect 169720 24432 556160 24460
rect 169720 24420 169726 24432
rect 556154 24420 556160 24432
rect 556212 24420 556218 24472
rect 168834 24352 168840 24404
rect 168892 24392 168898 24404
rect 563054 24392 563060 24404
rect 168892 24364 563060 24392
rect 168892 24352 168898 24364
rect 563054 24352 563060 24364
rect 563112 24352 563118 24404
rect 3326 24284 3332 24336
rect 3384 24324 3390 24336
rect 179874 24324 179880 24336
rect 3384 24296 179880 24324
rect 3384 24284 3390 24296
rect 179874 24284 179880 24296
rect 179932 24284 179938 24336
rect 183002 24284 183008 24336
rect 183060 24324 183066 24336
rect 579614 24324 579620 24336
rect 183060 24296 579620 24324
rect 183060 24284 183066 24296
rect 579614 24284 579620 24296
rect 579672 24284 579678 24336
rect 169938 24216 169944 24268
rect 169996 24256 170002 24268
rect 569954 24256 569960 24268
rect 169996 24228 569960 24256
rect 169996 24216 170002 24228
rect 569954 24216 569960 24228
rect 570012 24216 570018 24268
rect 169846 24148 169852 24200
rect 169904 24188 169910 24200
rect 571334 24188 571340 24200
rect 169904 24160 571340 24188
rect 169904 24148 169910 24160
rect 571334 24148 571340 24160
rect 571392 24148 571398 24200
rect 170030 24080 170036 24132
rect 170088 24120 170094 24132
rect 572806 24120 572812 24132
rect 170088 24092 572812 24120
rect 170088 24080 170094 24092
rect 572806 24080 572812 24092
rect 572864 24080 572870 24132
rect 320818 24012 320824 24064
rect 320876 24052 320882 24064
rect 327718 24052 327724 24064
rect 320876 24024 327724 24052
rect 320876 24012 320882 24024
rect 327718 24012 327724 24024
rect 327776 24012 327782 24064
rect 135990 23400 135996 23452
rect 136048 23440 136054 23452
rect 142338 23440 142344 23452
rect 136048 23412 142344 23440
rect 136048 23400 136054 23412
rect 142338 23400 142344 23412
rect 142396 23400 142402 23452
rect 319438 23400 319444 23452
rect 319496 23440 319502 23452
rect 326338 23440 326344 23452
rect 319496 23412 326344 23440
rect 319496 23400 319502 23412
rect 326338 23400 326344 23412
rect 326396 23400 326402 23452
rect 391198 23400 391204 23452
rect 391256 23440 391262 23452
rect 393314 23440 393320 23452
rect 391256 23412 393320 23440
rect 391256 23400 391262 23412
rect 393314 23400 393320 23412
rect 393372 23400 393378 23452
rect 302234 23264 302240 23316
rect 302292 23304 302298 23316
rect 313274 23304 313280 23316
rect 302292 23276 313280 23304
rect 302292 23264 302298 23276
rect 313274 23264 313280 23276
rect 313332 23264 313338 23316
rect 3418 23196 3424 23248
rect 3476 23236 3482 23248
rect 173986 23236 173992 23248
rect 3476 23208 173992 23236
rect 3476 23196 3482 23208
rect 173986 23196 173992 23208
rect 174044 23196 174050 23248
rect 284938 23196 284944 23248
rect 284996 23236 285002 23248
rect 299290 23236 299296 23248
rect 284996 23208 299296 23236
rect 284996 23196 285002 23208
rect 299290 23196 299296 23208
rect 299348 23196 299354 23248
rect 311158 23196 311164 23248
rect 311216 23236 311222 23248
rect 323578 23236 323584 23248
rect 311216 23208 323584 23236
rect 311216 23196 311222 23208
rect 323578 23196 323584 23208
rect 323636 23196 323642 23248
rect 356146 23196 356152 23248
rect 356204 23236 356210 23248
rect 369946 23236 369952 23248
rect 356204 23208 369952 23236
rect 356204 23196 356210 23208
rect 369946 23196 369952 23208
rect 370004 23196 370010 23248
rect 172238 23128 172244 23180
rect 172296 23168 172302 23180
rect 404354 23168 404360 23180
rect 172296 23140 404360 23168
rect 172296 23128 172302 23140
rect 404354 23128 404360 23140
rect 404412 23128 404418 23180
rect 163038 23060 163044 23112
rect 163096 23100 163102 23112
rect 492674 23100 492680 23112
rect 163096 23072 492680 23100
rect 163096 23060 163102 23072
rect 492674 23060 492680 23072
rect 492732 23060 492738 23112
rect 167362 22992 167368 23044
rect 167420 23032 167426 23044
rect 534074 23032 534080 23044
rect 167420 23004 534080 23032
rect 167420 22992 167426 23004
rect 534074 22992 534080 23004
rect 534132 22992 534138 23044
rect 63494 22924 63500 22976
rect 63552 22964 63558 22976
rect 126330 22964 126336 22976
rect 63552 22936 126336 22964
rect 63552 22924 63558 22936
rect 126330 22924 126336 22936
rect 126388 22924 126394 22976
rect 167454 22924 167460 22976
rect 167512 22964 167518 22976
rect 538214 22964 538220 22976
rect 167512 22936 538220 22964
rect 167512 22924 167518 22936
rect 538214 22924 538220 22936
rect 538272 22924 538278 22976
rect 35894 22856 35900 22908
rect 35952 22896 35958 22908
rect 126974 22896 126980 22908
rect 35952 22868 126980 22896
rect 35952 22856 35958 22868
rect 126974 22856 126980 22868
rect 127032 22856 127038 22908
rect 167178 22856 167184 22908
rect 167236 22896 167242 22908
rect 540974 22896 540980 22908
rect 167236 22868 540980 22896
rect 167236 22856 167242 22868
rect 540974 22856 540980 22868
rect 541032 22856 541038 22908
rect 22094 22788 22100 22840
rect 22152 22828 22158 22840
rect 127526 22828 127532 22840
rect 22152 22800 127532 22828
rect 22152 22788 22158 22800
rect 127526 22788 127532 22800
rect 127584 22788 127590 22840
rect 167270 22788 167276 22840
rect 167328 22828 167334 22840
rect 545114 22828 545120 22840
rect 167328 22800 545120 22828
rect 167328 22788 167334 22800
rect 545114 22788 545120 22800
rect 545172 22788 545178 22840
rect 118326 22720 118332 22772
rect 118384 22760 118390 22772
rect 580258 22760 580264 22772
rect 118384 22732 580264 22760
rect 118384 22720 118390 22732
rect 580258 22720 580264 22732
rect 580316 22720 580322 22772
rect 321738 22108 321744 22160
rect 321796 22148 321802 22160
rect 324314 22148 324320 22160
rect 321796 22120 324320 22148
rect 321796 22108 321802 22120
rect 324314 22108 324320 22120
rect 324372 22108 324378 22160
rect 301590 21768 301596 21820
rect 301648 21808 301654 21820
rect 304258 21808 304264 21820
rect 301648 21780 304264 21808
rect 301648 21768 301654 21780
rect 304258 21768 304264 21780
rect 304316 21768 304322 21820
rect 329098 21768 329104 21820
rect 329156 21808 329162 21820
rect 344278 21808 344284 21820
rect 329156 21780 344284 21808
rect 329156 21768 329162 21780
rect 344278 21768 344284 21780
rect 344336 21768 344342 21820
rect 152182 21700 152188 21752
rect 152240 21740 152246 21752
rect 343634 21740 343640 21752
rect 152240 21712 343640 21740
rect 152240 21700 152246 21712
rect 343634 21700 343640 21712
rect 343692 21700 343698 21752
rect 160738 21632 160744 21684
rect 160796 21672 160802 21684
rect 454034 21672 454040 21684
rect 160796 21644 454040 21672
rect 160796 21632 160802 21644
rect 454034 21632 454040 21644
rect 454092 21632 454098 21684
rect 165982 21564 165988 21616
rect 166040 21604 166046 21616
rect 516134 21604 516140 21616
rect 166040 21576 516140 21604
rect 166040 21564 166046 21576
rect 516134 21564 516140 21576
rect 516192 21564 516198 21616
rect 165798 21496 165804 21548
rect 165856 21536 165862 21548
rect 520274 21536 520280 21548
rect 165856 21508 520280 21536
rect 165856 21496 165862 21508
rect 520274 21496 520280 21508
rect 520332 21496 520338 21548
rect 165890 21428 165896 21480
rect 165948 21468 165954 21480
rect 523126 21468 523132 21480
rect 165948 21440 523132 21468
rect 165948 21428 165954 21440
rect 523126 21428 523132 21440
rect 523184 21428 523190 21480
rect 85574 21360 85580 21412
rect 85632 21400 85638 21412
rect 131758 21400 131764 21412
rect 85632 21372 131764 21400
rect 85632 21360 85638 21372
rect 131758 21360 131764 21372
rect 131816 21360 131822 21412
rect 166074 21360 166080 21412
rect 166132 21400 166138 21412
rect 527174 21400 527180 21412
rect 166132 21372 527180 21400
rect 166132 21360 166138 21372
rect 527174 21360 527180 21372
rect 527232 21360 527238 21412
rect 362218 20612 362224 20664
rect 362276 20652 362282 20664
rect 365070 20652 365076 20664
rect 362276 20624 365076 20652
rect 362276 20612 362282 20624
rect 365070 20612 365076 20624
rect 365128 20612 365134 20664
rect 396718 20612 396724 20664
rect 396776 20652 396782 20664
rect 398926 20652 398932 20664
rect 396776 20624 398932 20652
rect 396776 20612 396782 20624
rect 398926 20612 398932 20624
rect 398984 20612 398990 20664
rect 299290 20340 299296 20392
rect 299348 20380 299354 20392
rect 326522 20380 326528 20392
rect 299348 20352 326528 20380
rect 299348 20340 299354 20352
rect 326522 20340 326528 20352
rect 326580 20340 326586 20392
rect 145098 20272 145104 20324
rect 145156 20312 145162 20324
rect 262214 20312 262220 20324
rect 145156 20284 262220 20312
rect 145156 20272 145162 20284
rect 262214 20272 262220 20284
rect 262272 20272 262278 20324
rect 313274 20272 313280 20324
rect 313332 20312 313338 20324
rect 322198 20312 322204 20324
rect 313332 20284 322204 20312
rect 313332 20272 313338 20284
rect 322198 20272 322204 20284
rect 322256 20272 322262 20324
rect 323486 20272 323492 20324
rect 323544 20312 323550 20324
rect 358078 20312 358084 20324
rect 323544 20284 358084 20312
rect 323544 20272 323550 20284
rect 358078 20272 358084 20284
rect 358136 20272 358142 20324
rect 369854 20272 369860 20324
rect 369912 20312 369918 20324
rect 379514 20312 379520 20324
rect 369912 20284 379520 20312
rect 369912 20272 369918 20284
rect 379514 20272 379520 20284
rect 379572 20272 379578 20324
rect 145006 20204 145012 20256
rect 145064 20244 145070 20256
rect 255314 20244 255320 20256
rect 145064 20216 255320 20244
rect 145064 20204 145070 20216
rect 255314 20204 255320 20216
rect 255372 20204 255378 20256
rect 255958 20204 255964 20256
rect 256016 20244 256022 20256
rect 456794 20244 456800 20256
rect 256016 20216 456800 20244
rect 256016 20204 256022 20216
rect 456794 20204 456800 20216
rect 456852 20204 456858 20256
rect 143810 20136 143816 20188
rect 143868 20176 143874 20188
rect 241514 20176 241520 20188
rect 143868 20148 241520 20176
rect 143868 20136 143874 20148
rect 241514 20136 241520 20148
rect 241572 20136 241578 20188
rect 242158 20136 242164 20188
rect 242216 20176 242222 20188
rect 449894 20176 449900 20188
rect 242216 20148 449900 20176
rect 242216 20136 242222 20148
rect 449894 20136 449900 20148
rect 449952 20136 449958 20188
rect 157518 20068 157524 20120
rect 157576 20108 157582 20120
rect 415394 20108 415400 20120
rect 157576 20080 415400 20108
rect 157576 20068 157582 20080
rect 415394 20068 415400 20080
rect 415452 20068 415458 20120
rect 164418 20000 164424 20052
rect 164476 20040 164482 20052
rect 506566 20040 506572 20052
rect 164476 20012 506572 20040
rect 164476 20000 164482 20012
rect 506566 20000 506572 20012
rect 506624 20000 506630 20052
rect 164510 19932 164516 19984
rect 164568 19972 164574 19984
rect 509234 19972 509240 19984
rect 164568 19944 509240 19972
rect 164568 19932 164574 19944
rect 509234 19932 509240 19944
rect 509292 19932 509298 19984
rect 356698 19252 356704 19304
rect 356756 19292 356762 19304
rect 359550 19292 359556 19304
rect 356756 19264 359556 19292
rect 356756 19252 356762 19264
rect 359550 19252 359556 19264
rect 359608 19252 359614 19304
rect 369118 18980 369124 19032
rect 369176 19020 369182 19032
rect 378686 19020 378692 19032
rect 369176 18992 378692 19020
rect 369176 18980 369182 18992
rect 378686 18980 378692 18992
rect 378744 18980 378750 19032
rect 359458 18912 359464 18964
rect 359516 18952 359522 18964
rect 377398 18952 377404 18964
rect 359516 18924 377404 18952
rect 359516 18912 359522 18924
rect 377398 18912 377404 18924
rect 377456 18912 377462 18964
rect 143718 18844 143724 18896
rect 143776 18884 143782 18896
rect 234614 18884 234620 18896
rect 143776 18856 234620 18884
rect 143776 18844 143782 18856
rect 234614 18844 234620 18856
rect 234672 18844 234678 18896
rect 275278 18844 275284 18896
rect 275336 18884 275342 18896
rect 288434 18884 288440 18896
rect 275336 18856 288440 18884
rect 275336 18844 275342 18856
rect 288434 18844 288440 18856
rect 288492 18844 288498 18896
rect 292758 18844 292764 18896
rect 292816 18884 292822 18896
rect 302050 18884 302056 18896
rect 292816 18856 302056 18884
rect 292816 18844 292822 18856
rect 302050 18844 302056 18856
rect 302108 18844 302114 18896
rect 347038 18844 347044 18896
rect 347096 18884 347102 18896
rect 388530 18884 388536 18896
rect 347096 18856 388536 18884
rect 347096 18844 347102 18856
rect 388530 18844 388536 18856
rect 388588 18844 388594 18896
rect 164234 18776 164240 18828
rect 164292 18816 164298 18828
rect 498286 18816 498292 18828
rect 164292 18788 498292 18816
rect 164292 18776 164298 18788
rect 498286 18776 498292 18788
rect 498344 18776 498350 18828
rect 164326 18708 164332 18760
rect 164384 18748 164390 18760
rect 502334 18748 502340 18760
rect 164384 18720 502340 18748
rect 164384 18708 164390 18720
rect 502334 18708 502340 18720
rect 502392 18708 502398 18760
rect 168466 18640 168472 18692
rect 168524 18680 168530 18692
rect 553394 18680 553400 18692
rect 168524 18652 553400 18680
rect 168524 18640 168530 18652
rect 553394 18640 553400 18652
rect 553452 18640 553458 18692
rect 81434 18572 81440 18624
rect 81492 18612 81498 18624
rect 131666 18612 131672 18624
rect 81492 18584 131672 18612
rect 81492 18572 81498 18584
rect 131666 18572 131672 18584
rect 131724 18572 131730 18624
rect 168558 18572 168564 18624
rect 168616 18612 168622 18624
rect 556246 18612 556252 18624
rect 168616 18584 556252 18612
rect 168616 18572 168622 18584
rect 556246 18572 556252 18584
rect 556304 18572 556310 18624
rect 351822 18028 351828 18080
rect 351880 18068 351886 18080
rect 354766 18068 354772 18080
rect 351880 18040 354772 18068
rect 351880 18028 351886 18040
rect 354766 18028 354772 18040
rect 354824 18028 354830 18080
rect 400858 17960 400864 18012
rect 400916 18000 400922 18012
rect 402974 18000 402980 18012
rect 400916 17972 402980 18000
rect 400916 17960 400922 17972
rect 402974 17960 402980 17972
rect 403032 17960 403038 18012
rect 365162 17892 365168 17944
rect 365220 17932 365226 17944
rect 373442 17932 373448 17944
rect 365220 17904 373448 17932
rect 365220 17892 365226 17904
rect 373442 17892 373448 17904
rect 373500 17892 373506 17944
rect 379514 17892 379520 17944
rect 379572 17932 379578 17944
rect 382274 17932 382280 17944
rect 379572 17904 382280 17932
rect 379572 17892 379578 17904
rect 382274 17892 382280 17904
rect 382332 17892 382338 17944
rect 369946 17348 369952 17400
rect 370004 17388 370010 17400
rect 375374 17388 375380 17400
rect 370004 17360 375380 17388
rect 370004 17348 370010 17360
rect 375374 17348 375380 17360
rect 375432 17348 375438 17400
rect 342254 17212 342260 17264
rect 342312 17252 342318 17264
rect 348694 17252 348700 17264
rect 342312 17224 348700 17252
rect 342312 17212 342318 17224
rect 348694 17212 348700 17224
rect 348752 17212 348758 17264
rect 392578 17212 392584 17264
rect 392636 17252 392642 17264
rect 397178 17252 397184 17264
rect 392636 17224 397184 17252
rect 392636 17212 392642 17224
rect 397178 17212 397184 17224
rect 397236 17212 397242 17264
rect 324314 17008 324320 17060
rect 324372 17048 324378 17060
rect 327074 17048 327080 17060
rect 324372 17020 327080 17048
rect 324372 17008 324378 17020
rect 327074 17008 327080 17020
rect 327132 17008 327138 17060
rect 143626 16124 143632 16176
rect 143684 16164 143690 16176
rect 237650 16164 237656 16176
rect 143684 16136 237656 16164
rect 143684 16124 143690 16136
rect 237650 16124 237656 16136
rect 237708 16124 237714 16176
rect 288434 16124 288440 16176
rect 288492 16164 288498 16176
rect 298738 16164 298744 16176
rect 288492 16136 298744 16164
rect 288492 16124 288498 16136
rect 298738 16124 298744 16136
rect 298796 16124 298802 16176
rect 302878 16124 302884 16176
rect 302936 16164 302942 16176
rect 313918 16164 313924 16176
rect 302936 16136 313924 16164
rect 302936 16124 302942 16136
rect 313918 16124 313924 16136
rect 313976 16124 313982 16176
rect 326522 16124 326528 16176
rect 326580 16164 326586 16176
rect 337010 16164 337016 16176
rect 326580 16136 337016 16164
rect 326580 16124 326586 16136
rect 337010 16124 337016 16136
rect 337068 16124 337074 16176
rect 152090 16056 152096 16108
rect 152148 16096 152154 16108
rect 342898 16096 342904 16108
rect 152148 16068 342904 16096
rect 152148 16056 152154 16068
rect 342898 16056 342904 16068
rect 342956 16056 342962 16108
rect 344278 16056 344284 16108
rect 344336 16096 344342 16108
rect 357342 16096 357348 16108
rect 344336 16068 357348 16096
rect 344336 16056 344342 16068
rect 357342 16056 357348 16068
rect 357400 16056 357406 16108
rect 358078 16056 358084 16108
rect 358136 16096 358142 16108
rect 385862 16096 385868 16108
rect 358136 16068 385868 16096
rect 358136 16056 358142 16068
rect 385862 16056 385868 16068
rect 385920 16056 385926 16108
rect 153470 15988 153476 16040
rect 153528 16028 153534 16040
rect 361114 16028 361120 16040
rect 153528 16000 361120 16028
rect 153528 15988 153534 16000
rect 361114 15988 361120 16000
rect 361172 15988 361178 16040
rect 385678 15988 385684 16040
rect 385736 16028 385742 16040
rect 390554 16028 390560 16040
rect 385736 16000 390560 16028
rect 385736 15988 385742 16000
rect 390554 15988 390560 16000
rect 390612 15988 390618 16040
rect 157426 15920 157432 15972
rect 157484 15960 157490 15972
rect 415486 15960 415492 15972
rect 157484 15932 415492 15960
rect 157484 15920 157490 15932
rect 415486 15920 415492 15932
rect 415544 15920 415550 15972
rect 157334 15852 157340 15904
rect 157392 15892 157398 15904
rect 420178 15892 420184 15904
rect 157392 15864 420184 15892
rect 157392 15852 157398 15864
rect 420178 15852 420184 15864
rect 420236 15852 420242 15904
rect 302050 15240 302056 15292
rect 302108 15280 302114 15292
rect 304258 15280 304264 15292
rect 302108 15252 304264 15280
rect 302108 15240 302114 15252
rect 304258 15240 304264 15252
rect 304316 15240 304322 15292
rect 380158 15172 380164 15224
rect 380216 15212 380222 15224
rect 382918 15212 382924 15224
rect 380216 15184 382924 15212
rect 380216 15172 380222 15184
rect 382918 15172 382924 15184
rect 382976 15172 382982 15224
rect 305638 14832 305644 14884
rect 305696 14872 305702 14884
rect 309594 14872 309600 14884
rect 305696 14844 309600 14872
rect 305696 14832 305702 14844
rect 309594 14832 309600 14844
rect 309652 14832 309658 14884
rect 149422 14764 149428 14816
rect 149480 14804 149486 14816
rect 311434 14804 311440 14816
rect 149480 14776 311440 14804
rect 149480 14764 149486 14776
rect 311434 14764 311440 14776
rect 311492 14764 311498 14816
rect 382366 14804 382372 14816
rect 373966 14776 382372 14804
rect 159634 14696 159640 14748
rect 159692 14736 159698 14748
rect 373966 14736 373994 14776
rect 382366 14764 382372 14776
rect 382424 14764 382430 14816
rect 159692 14708 373994 14736
rect 159692 14696 159698 14708
rect 382274 14696 382280 14748
rect 382332 14736 382338 14748
rect 402514 14736 402520 14748
rect 382332 14708 402520 14736
rect 382332 14696 382338 14708
rect 402514 14696 402520 14708
rect 402572 14696 402578 14748
rect 159266 14628 159272 14680
rect 159324 14668 159330 14680
rect 429194 14668 429200 14680
rect 159324 14640 429200 14668
rect 159324 14628 159330 14640
rect 429194 14628 429200 14640
rect 429252 14628 429258 14680
rect 159358 14560 159364 14612
rect 159416 14600 159422 14612
rect 436738 14600 436744 14612
rect 159416 14572 436744 14600
rect 159416 14560 159422 14572
rect 436738 14560 436744 14572
rect 436796 14560 436802 14612
rect 159174 14492 159180 14544
rect 159232 14532 159238 14544
rect 439130 14532 439136 14544
rect 159232 14504 439136 14532
rect 159232 14492 159238 14504
rect 439130 14492 439136 14504
rect 439188 14492 439194 14544
rect 162946 14424 162952 14476
rect 163004 14464 163010 14476
rect 492306 14464 492312 14476
rect 163004 14436 492312 14464
rect 163004 14424 163010 14436
rect 492306 14424 492312 14436
rect 492364 14424 492370 14476
rect 377398 13812 377404 13864
rect 377456 13852 377462 13864
rect 380894 13852 380900 13864
rect 377456 13824 380900 13852
rect 377456 13812 377462 13824
rect 380894 13812 380900 13824
rect 380952 13812 380958 13864
rect 304258 13744 304264 13796
rect 304316 13784 304322 13796
rect 307018 13784 307024 13796
rect 304316 13756 307024 13784
rect 304316 13744 304322 13756
rect 307018 13744 307024 13756
rect 307076 13744 307082 13796
rect 385862 13744 385868 13796
rect 385920 13784 385926 13796
rect 392578 13784 392584 13796
rect 385920 13756 392584 13784
rect 385920 13744 385926 13756
rect 392578 13744 392584 13756
rect 392636 13744 392642 13796
rect 153286 13132 153292 13184
rect 153344 13172 153350 13184
rect 357526 13172 357532 13184
rect 153344 13144 357532 13172
rect 153344 13132 153350 13144
rect 357526 13132 357532 13144
rect 357584 13132 357590 13184
rect 153378 13064 153384 13116
rect 153436 13104 153442 13116
rect 365806 13104 365812 13116
rect 153436 13076 365812 13104
rect 153436 13064 153442 13076
rect 365806 13064 365812 13076
rect 365864 13064 365870 13116
rect 375374 13064 375380 13116
rect 375432 13104 375438 13116
rect 381722 13104 381728 13116
rect 375432 13076 381728 13104
rect 375432 13064 375438 13076
rect 381722 13064 381728 13076
rect 381780 13064 381786 13116
rect 323578 12384 323584 12436
rect 323636 12424 323642 12436
rect 326246 12424 326252 12436
rect 323636 12396 326252 12424
rect 323636 12384 323642 12396
rect 326246 12384 326252 12396
rect 326304 12384 326310 12436
rect 348694 12384 348700 12436
rect 348752 12424 348758 12436
rect 357066 12424 357072 12436
rect 348752 12396 357072 12424
rect 348752 12384 348758 12396
rect 357066 12384 357072 12396
rect 357124 12384 357130 12436
rect 381630 12384 381636 12436
rect 381688 12424 381694 12436
rect 384390 12424 384396 12436
rect 381688 12396 384396 12424
rect 381688 12384 381694 12396
rect 384390 12384 384396 12396
rect 384448 12384 384454 12436
rect 390554 12384 390560 12436
rect 390612 12424 390618 12436
rect 395338 12424 395344 12436
rect 390612 12396 395344 12424
rect 390612 12384 390618 12396
rect 395338 12384 395344 12396
rect 395396 12384 395402 12436
rect 397178 12384 397184 12436
rect 397236 12424 397242 12436
rect 403710 12424 403716 12436
rect 397236 12396 403716 12424
rect 397236 12384 397242 12396
rect 403710 12384 403716 12396
rect 403768 12384 403774 12436
rect 304350 12316 304356 12368
rect 304408 12356 304414 12368
rect 312538 12356 312544 12368
rect 304408 12328 312544 12356
rect 304408 12316 304414 12328
rect 312538 12316 312544 12328
rect 312596 12316 312602 12368
rect 326430 12316 326436 12368
rect 326488 12356 326494 12368
rect 332686 12356 332692 12368
rect 326488 12328 332692 12356
rect 326488 12316 326494 12328
rect 332686 12316 332692 12328
rect 332744 12316 332750 12368
rect 151998 12248 152004 12300
rect 152056 12288 152062 12300
rect 345290 12288 345296 12300
rect 152056 12260 345296 12288
rect 152056 12248 152062 12260
rect 345290 12248 345296 12260
rect 345348 12248 345354 12300
rect 357342 12248 357348 12300
rect 357400 12288 357406 12300
rect 373350 12288 373356 12300
rect 357400 12260 373356 12288
rect 357400 12248 357406 12260
rect 373350 12248 373356 12260
rect 373408 12248 373414 12300
rect 373442 12248 373448 12300
rect 373500 12288 373506 12300
rect 379514 12288 379520 12300
rect 373500 12260 379520 12288
rect 373500 12248 373506 12260
rect 379514 12248 379520 12260
rect 379572 12248 379578 12300
rect 151906 12180 151912 12232
rect 151964 12220 151970 12232
rect 349246 12220 349252 12232
rect 151964 12192 349252 12220
rect 151964 12180 151970 12192
rect 349246 12180 349252 12192
rect 349304 12180 349310 12232
rect 354766 12180 354772 12232
rect 354824 12220 354830 12232
rect 376018 12220 376024 12232
rect 354824 12192 376024 12220
rect 354824 12180 354830 12192
rect 376018 12180 376024 12192
rect 376076 12180 376082 12232
rect 162210 12112 162216 12164
rect 162268 12152 162274 12164
rect 390646 12152 390652 12164
rect 162268 12124 390652 12152
rect 162268 12112 162274 12124
rect 390646 12112 390652 12124
rect 390704 12112 390710 12164
rect 159082 12044 159088 12096
rect 159140 12084 159146 12096
rect 428458 12084 428464 12096
rect 159140 12056 428464 12084
rect 159140 12044 159146 12056
rect 428458 12044 428464 12056
rect 428516 12044 428522 12096
rect 158898 11976 158904 12028
rect 158956 12016 158962 12028
rect 432046 12016 432052 12028
rect 158956 11988 432052 12016
rect 158956 11976 158962 11988
rect 432046 11976 432052 11988
rect 432104 11976 432110 12028
rect 158806 11908 158812 11960
rect 158864 11948 158870 11960
rect 435082 11948 435088 11960
rect 158864 11920 435088 11948
rect 158864 11908 158870 11920
rect 435082 11908 435088 11920
rect 435140 11908 435146 11960
rect 160002 11840 160008 11892
rect 160060 11880 160066 11892
rect 440326 11880 440332 11892
rect 160060 11852 440332 11880
rect 160060 11840 160066 11852
rect 440326 11840 440332 11852
rect 440384 11840 440390 11892
rect 162026 11772 162032 11824
rect 162084 11812 162090 11824
rect 468202 11812 468208 11824
rect 162084 11784 468208 11812
rect 162084 11772 162090 11784
rect 468202 11772 468208 11784
rect 468260 11772 468266 11824
rect 169754 11704 169760 11756
rect 169812 11744 169818 11756
rect 574646 11744 574652 11756
rect 169812 11716 574652 11744
rect 169812 11704 169818 11716
rect 574646 11704 574652 11716
rect 574704 11704 574710 11756
rect 364978 11636 364984 11688
rect 365036 11676 365042 11688
rect 367738 11676 367744 11688
rect 365036 11648 367744 11676
rect 365036 11636 365042 11648
rect 367738 11636 367744 11648
rect 367796 11636 367802 11688
rect 378686 11636 378692 11688
rect 378744 11676 378750 11688
rect 381262 11676 381268 11688
rect 378744 11648 381268 11676
rect 378744 11636 378750 11648
rect 381262 11636 381268 11648
rect 381320 11636 381326 11688
rect 117314 10548 117320 10600
rect 117372 10588 117378 10600
rect 134242 10588 134248 10600
rect 117372 10560 134248 10588
rect 117372 10548 117378 10560
rect 134242 10548 134248 10560
rect 134300 10548 134306 10600
rect 106458 10480 106464 10532
rect 106516 10520 106522 10532
rect 133046 10520 133052 10532
rect 106516 10492 133052 10520
rect 106516 10480 106522 10492
rect 133046 10480 133052 10492
rect 133104 10480 133110 10532
rect 78122 10412 78128 10464
rect 78180 10452 78186 10464
rect 129090 10452 129096 10464
rect 78180 10424 129096 10452
rect 78180 10412 78186 10424
rect 129090 10412 129096 10424
rect 129148 10412 129154 10464
rect 149330 10412 149336 10464
rect 149388 10452 149394 10464
rect 309778 10452 309784 10464
rect 149388 10424 309784 10452
rect 149388 10412 149394 10424
rect 309778 10412 309784 10424
rect 309836 10412 309842 10464
rect 25314 10344 25320 10396
rect 25372 10384 25378 10396
rect 93118 10384 93124 10396
rect 25372 10356 93124 10384
rect 25372 10344 25378 10356
rect 93118 10344 93124 10356
rect 93176 10344 93182 10396
rect 99834 10344 99840 10396
rect 99892 10384 99898 10396
rect 132954 10384 132960 10396
rect 99892 10356 132960 10384
rect 99892 10344 99898 10356
rect 132954 10344 132960 10356
rect 133012 10344 133018 10396
rect 149238 10344 149244 10396
rect 149296 10384 149302 10396
rect 313826 10384 313832 10396
rect 149296 10356 313832 10384
rect 149296 10344 149302 10356
rect 313826 10344 313832 10356
rect 313884 10344 313890 10396
rect 35986 10276 35992 10328
rect 36044 10316 36050 10328
rect 127434 10316 127440 10328
rect 36044 10288 127440 10316
rect 36044 10276 36050 10288
rect 127434 10276 127440 10288
rect 127492 10276 127498 10328
rect 166994 10276 167000 10328
rect 167052 10316 167058 10328
rect 542722 10316 542728 10328
rect 167052 10288 542728 10316
rect 167052 10276 167058 10288
rect 542722 10276 542728 10288
rect 542780 10276 542786 10328
rect 147766 9596 147772 9648
rect 147824 9636 147830 9648
rect 296070 9636 296076 9648
rect 147824 9608 296076 9636
rect 147824 9596 147830 9608
rect 296070 9596 296076 9608
rect 296128 9596 296134 9648
rect 309594 9596 309600 9648
rect 309652 9636 309658 9648
rect 313090 9636 313096 9648
rect 309652 9608 313096 9636
rect 309652 9596 309658 9608
rect 313090 9596 313096 9608
rect 313148 9596 313154 9648
rect 315298 9596 315304 9648
rect 315356 9636 315362 9648
rect 465166 9636 465172 9648
rect 315356 9608 465172 9636
rect 315356 9596 315362 9608
rect 465166 9596 465172 9608
rect 465224 9596 465230 9648
rect 160186 9528 160192 9580
rect 160244 9568 160250 9580
rect 445018 9568 445024 9580
rect 160244 9540 445024 9568
rect 160244 9528 160250 9540
rect 445018 9528 445024 9540
rect 445076 9528 445082 9580
rect 165706 9460 165712 9512
rect 165764 9500 165770 9512
rect 449894 9500 449900 9512
rect 165764 9472 449900 9500
rect 165764 9460 165770 9472
rect 449894 9460 449900 9472
rect 449952 9460 449958 9512
rect 160278 9392 160284 9444
rect 160336 9432 160342 9444
rect 446214 9432 446220 9444
rect 160336 9404 446220 9432
rect 160336 9392 160342 9404
rect 446214 9392 446220 9404
rect 446272 9392 446278 9444
rect 160462 9324 160468 9376
rect 160520 9364 160526 9376
rect 448606 9364 448612 9376
rect 160520 9336 448612 9364
rect 160520 9324 160526 9336
rect 448606 9324 448612 9336
rect 448664 9324 448670 9376
rect 60826 9256 60832 9308
rect 60884 9296 60890 9308
rect 128354 9296 128360 9308
rect 60884 9268 128360 9296
rect 60884 9256 60890 9268
rect 128354 9256 128360 9268
rect 128412 9256 128418 9308
rect 161198 9256 161204 9308
rect 161256 9296 161262 9308
rect 449802 9296 449808 9308
rect 161256 9268 449808 9296
rect 161256 9256 161262 9268
rect 449802 9256 449808 9268
rect 449860 9256 449866 9308
rect 59630 9188 59636 9240
rect 59688 9228 59694 9240
rect 130102 9228 130108 9240
rect 59688 9200 130108 9228
rect 59688 9188 59694 9200
rect 130102 9188 130108 9200
rect 130160 9188 130166 9240
rect 160554 9188 160560 9240
rect 160612 9228 160618 9240
rect 452102 9228 452108 9240
rect 160612 9200 452108 9228
rect 160612 9188 160618 9200
rect 452102 9188 452108 9200
rect 452160 9188 452166 9240
rect 53742 9120 53748 9172
rect 53800 9160 53806 9172
rect 128722 9160 128728 9172
rect 53800 9132 128728 9160
rect 53800 9120 53806 9132
rect 128722 9120 128728 9132
rect 128780 9120 128786 9172
rect 160370 9120 160376 9172
rect 160428 9160 160434 9172
rect 453298 9160 453304 9172
rect 160428 9132 453304 9160
rect 160428 9120 160434 9132
rect 453298 9120 453304 9132
rect 453356 9120 453362 9172
rect 52546 9052 52552 9104
rect 52604 9092 52610 9104
rect 128630 9092 128636 9104
rect 52604 9064 128636 9092
rect 52604 9052 52610 9064
rect 128630 9052 128636 9064
rect 128688 9052 128694 9104
rect 160646 9052 160652 9104
rect 160704 9092 160710 9104
rect 455690 9092 455696 9104
rect 160704 9064 455696 9092
rect 160704 9052 160710 9064
rect 455690 9052 455696 9064
rect 455748 9052 455754 9104
rect 45462 8984 45468 9036
rect 45520 9024 45526 9036
rect 128538 9024 128544 9036
rect 45520 8996 128544 9024
rect 45520 8984 45526 8996
rect 128538 8984 128544 8996
rect 128596 8984 128602 9036
rect 161842 8984 161848 9036
rect 161900 9024 161906 9036
rect 463970 9024 463976 9036
rect 161900 8996 463976 9024
rect 161900 8984 161906 8996
rect 463970 8984 463976 8996
rect 464028 8984 464034 9036
rect 9950 8916 9956 8968
rect 10008 8956 10014 8968
rect 126146 8956 126152 8968
rect 10008 8928 126152 8956
rect 10008 8916 10014 8928
rect 126146 8916 126152 8928
rect 126204 8916 126210 8968
rect 161934 8916 161940 8968
rect 161992 8956 161998 8968
rect 467466 8956 467472 8968
rect 161992 8928 467472 8956
rect 161992 8916 161998 8928
rect 467466 8916 467472 8928
rect 467524 8916 467530 8968
rect 327718 8848 327724 8900
rect 327776 8888 327782 8900
rect 330386 8888 330392 8900
rect 327776 8860 330392 8888
rect 327776 8848 327782 8860
rect 330386 8848 330392 8860
rect 330444 8848 330450 8900
rect 357066 8848 357072 8900
rect 357124 8888 357130 8900
rect 362310 8888 362316 8900
rect 357124 8860 362316 8888
rect 357124 8848 357130 8860
rect 362310 8848 362316 8860
rect 362368 8848 362374 8900
rect 322198 8304 322204 8356
rect 322256 8344 322262 8356
rect 327074 8344 327080 8356
rect 322256 8316 327080 8344
rect 322256 8304 322262 8316
rect 327074 8304 327080 8316
rect 327132 8304 327138 8356
rect 116394 8032 116400 8084
rect 116452 8072 116458 8084
rect 134150 8072 134156 8084
rect 116452 8044 134156 8072
rect 116452 8032 116458 8044
rect 134150 8032 134156 8044
rect 134208 8032 134214 8084
rect 105722 7964 105728 8016
rect 105780 8004 105786 8016
rect 132862 8004 132868 8016
rect 105780 7976 132868 8004
rect 105780 7964 105786 7976
rect 132862 7964 132868 7976
rect 132920 7964 132926 8016
rect 98638 7896 98644 7948
rect 98696 7936 98702 7948
rect 132770 7936 132776 7948
rect 98696 7908 132776 7936
rect 98696 7896 98702 7908
rect 132770 7896 132776 7908
rect 132828 7896 132834 7948
rect 142246 7896 142252 7948
rect 142304 7936 142310 7948
rect 222746 7936 222752 7948
rect 142304 7908 222752 7936
rect 142304 7896 142310 7908
rect 222746 7896 222752 7908
rect 222804 7896 222810 7948
rect 84470 7828 84476 7880
rect 84528 7868 84534 7880
rect 131574 7868 131580 7880
rect 84528 7840 131580 7868
rect 84528 7828 84534 7840
rect 131574 7828 131580 7840
rect 131632 7828 131638 7880
rect 143534 7828 143540 7880
rect 143592 7868 143598 7880
rect 242986 7868 242992 7880
rect 143592 7840 242992 7868
rect 143592 7828 143598 7840
rect 242986 7828 242992 7840
rect 243044 7828 243050 7880
rect 48958 7760 48964 7812
rect 49016 7800 49022 7812
rect 129182 7800 129188 7812
rect 49016 7772 129188 7800
rect 49016 7760 49022 7772
rect 129182 7760 129188 7772
rect 129240 7760 129246 7812
rect 144914 7760 144920 7812
rect 144972 7800 144978 7812
rect 260650 7800 260656 7812
rect 144972 7772 260656 7800
rect 144972 7760 144978 7772
rect 260650 7760 260656 7772
rect 260708 7760 260714 7812
rect 34790 7692 34796 7744
rect 34848 7732 34854 7744
rect 127342 7732 127348 7744
rect 34848 7704 127348 7732
rect 34848 7692 34854 7704
rect 127342 7692 127348 7704
rect 127400 7692 127406 7744
rect 147030 7692 147036 7744
rect 147088 7732 147094 7744
rect 278314 7732 278320 7744
rect 147088 7704 278320 7732
rect 147088 7692 147094 7704
rect 278314 7692 278320 7704
rect 278372 7692 278378 7744
rect 373258 7692 373264 7744
rect 373316 7732 373322 7744
rect 381170 7732 381176 7744
rect 373316 7704 381176 7732
rect 373316 7692 373322 7704
rect 381170 7692 381176 7704
rect 381228 7692 381234 7744
rect 381538 7692 381544 7744
rect 381596 7732 381602 7744
rect 391842 7732 391848 7744
rect 381596 7704 391848 7732
rect 381596 7692 381602 7704
rect 391842 7692 391848 7704
rect 391900 7692 391906 7744
rect 24210 7624 24216 7676
rect 24268 7664 24274 7676
rect 122098 7664 122104 7676
rect 24268 7636 122104 7664
rect 24268 7624 24274 7636
rect 122098 7624 122104 7636
rect 122156 7624 122162 7676
rect 149054 7624 149060 7676
rect 149112 7664 149118 7676
rect 307938 7664 307944 7676
rect 149112 7636 307944 7664
rect 149112 7624 149118 7636
rect 307938 7624 307944 7636
rect 307996 7624 308002 7676
rect 365070 7624 365076 7676
rect 365128 7664 365134 7676
rect 376478 7664 376484 7676
rect 365128 7636 376484 7664
rect 365128 7624 365134 7636
rect 376478 7624 376484 7636
rect 376536 7624 376542 7676
rect 380894 7624 380900 7676
rect 380952 7664 380958 7676
rect 393038 7664 393044 7676
rect 380952 7636 393044 7664
rect 380952 7624 380958 7636
rect 393038 7624 393044 7636
rect 393096 7624 393102 7676
rect 27706 7556 27712 7608
rect 27764 7596 27770 7608
rect 127250 7596 127256 7608
rect 27764 7568 127256 7596
rect 27764 7556 27770 7568
rect 127250 7556 127256 7568
rect 127308 7556 127314 7608
rect 165614 7556 165620 7608
rect 165672 7596 165678 7608
rect 449158 7596 449164 7608
rect 165672 7568 449164 7596
rect 165672 7556 165678 7568
rect 449158 7556 449164 7568
rect 449216 7556 449222 7608
rect 381262 6876 381268 6928
rect 381320 6916 381326 6928
rect 384758 6916 384764 6928
rect 381320 6888 384764 6916
rect 381320 6876 381326 6888
rect 384758 6876 384764 6888
rect 384816 6876 384822 6928
rect 140774 6808 140780 6860
rect 140832 6848 140838 6860
rect 203886 6848 203892 6860
rect 140832 6820 203892 6848
rect 140832 6808 140838 6820
rect 203886 6808 203892 6820
rect 203944 6808 203950 6860
rect 162302 6740 162308 6792
rect 162360 6780 162366 6792
rect 235810 6780 235816 6792
rect 162360 6752 235816 6780
rect 162360 6740 162366 6752
rect 235810 6740 235816 6752
rect 235868 6740 235874 6792
rect 160922 6672 160928 6724
rect 160980 6712 160986 6724
rect 271230 6712 271236 6724
rect 160980 6684 271236 6712
rect 160980 6672 160986 6684
rect 271230 6672 271236 6684
rect 271288 6672 271294 6724
rect 104526 6604 104532 6656
rect 104584 6644 104590 6656
rect 132678 6644 132684 6656
rect 104584 6616 132684 6644
rect 104584 6604 104590 6616
rect 132678 6604 132684 6616
rect 132736 6604 132742 6656
rect 146938 6604 146944 6656
rect 146996 6644 147002 6656
rect 270034 6644 270040 6656
rect 146996 6616 270040 6644
rect 146996 6604 147002 6616
rect 270034 6604 270040 6616
rect 270092 6604 270098 6656
rect 80882 6536 80888 6588
rect 80940 6576 80946 6588
rect 131482 6576 131488 6588
rect 80940 6548 131488 6576
rect 80940 6536 80946 6548
rect 131482 6536 131488 6548
rect 131540 6536 131546 6588
rect 146846 6536 146852 6588
rect 146904 6576 146910 6588
rect 273622 6576 273628 6588
rect 146904 6548 273628 6576
rect 146904 6536 146910 6548
rect 273622 6536 273628 6548
rect 273680 6536 273686 6588
rect 77386 6468 77392 6520
rect 77444 6508 77450 6520
rect 131390 6508 131396 6520
rect 77444 6480 131396 6508
rect 77444 6468 77450 6480
rect 131390 6468 131396 6480
rect 131448 6468 131454 6520
rect 146754 6468 146760 6520
rect 146812 6508 146818 6520
rect 276014 6508 276020 6520
rect 146812 6480 276020 6508
rect 146812 6468 146818 6480
rect 276014 6468 276020 6480
rect 276072 6468 276078 6520
rect 313918 6468 313924 6520
rect 313976 6508 313982 6520
rect 322750 6508 322756 6520
rect 313976 6480 322756 6508
rect 313976 6468 313982 6480
rect 322750 6468 322756 6480
rect 322808 6468 322814 6520
rect 66714 6400 66720 6452
rect 66772 6440 66778 6452
rect 130010 6440 130016 6452
rect 66772 6412 130016 6440
rect 66772 6400 66778 6412
rect 130010 6400 130016 6412
rect 130068 6400 130074 6452
rect 146570 6400 146576 6452
rect 146628 6440 146634 6452
rect 277118 6440 277124 6452
rect 146628 6412 277124 6440
rect 146628 6400 146634 6412
rect 277118 6400 277124 6412
rect 277176 6400 277182 6452
rect 307018 6400 307024 6452
rect 307076 6440 307082 6452
rect 329190 6440 329196 6452
rect 307076 6412 329196 6440
rect 307076 6400 307082 6412
rect 329190 6400 329196 6412
rect 329248 6400 329254 6452
rect 44266 6332 44272 6384
rect 44324 6372 44330 6384
rect 128814 6372 128820 6384
rect 44324 6344 128820 6372
rect 44324 6332 44330 6344
rect 128814 6332 128820 6344
rect 128872 6332 128878 6384
rect 146662 6332 146668 6384
rect 146720 6372 146726 6384
rect 279510 6372 279516 6384
rect 146720 6344 279516 6372
rect 146720 6332 146726 6344
rect 279510 6332 279516 6344
rect 279568 6332 279574 6384
rect 298738 6332 298744 6384
rect 298796 6372 298802 6384
rect 320910 6372 320916 6384
rect 298796 6344 320916 6372
rect 298796 6332 298802 6344
rect 320910 6332 320916 6344
rect 320968 6332 320974 6384
rect 392578 6332 392584 6384
rect 392636 6372 392642 6384
rect 398098 6372 398104 6384
rect 392636 6344 398104 6372
rect 392636 6332 392642 6344
rect 398098 6332 398104 6344
rect 398156 6332 398162 6384
rect 33594 6264 33600 6316
rect 33652 6304 33658 6316
rect 127158 6304 127164 6316
rect 33652 6276 127164 6304
rect 33652 6264 33658 6276
rect 127158 6264 127164 6276
rect 127216 6264 127222 6316
rect 151814 6264 151820 6316
rect 151872 6304 151878 6316
rect 348050 6304 348056 6316
rect 151872 6276 348056 6304
rect 151872 6264 151878 6276
rect 348050 6264 348056 6276
rect 348108 6264 348114 6316
rect 373350 6264 373356 6316
rect 373408 6304 373414 6316
rect 378042 6304 378048 6316
rect 373408 6276 378048 6304
rect 373408 6264 373414 6276
rect 378042 6264 378048 6276
rect 378100 6264 378106 6316
rect 381722 6264 381728 6316
rect 381780 6304 381786 6316
rect 395246 6304 395252 6316
rect 381780 6276 395252 6304
rect 381780 6264 381786 6276
rect 395246 6264 395252 6276
rect 395304 6264 395310 6316
rect 19426 6196 19432 6248
rect 19484 6236 19490 6248
rect 124950 6236 124956 6248
rect 19484 6208 124956 6236
rect 19484 6196 19490 6208
rect 124950 6196 124956 6208
rect 125008 6196 125014 6248
rect 161750 6196 161756 6248
rect 161808 6236 161814 6248
rect 471054 6236 471060 6248
rect 161808 6208 471060 6236
rect 161808 6196 161814 6208
rect 471054 6196 471060 6208
rect 471112 6196 471118 6248
rect 18230 6128 18236 6180
rect 18288 6168 18294 6180
rect 126054 6168 126060 6180
rect 18288 6140 126060 6168
rect 18288 6128 18294 6140
rect 126054 6128 126060 6140
rect 126112 6128 126118 6180
rect 137094 6128 137100 6180
rect 137152 6168 137158 6180
rect 145926 6168 145932 6180
rect 137152 6140 145932 6168
rect 137152 6128 137158 6140
rect 145926 6128 145932 6140
rect 145984 6128 145990 6180
rect 171042 6128 171048 6180
rect 171100 6168 171106 6180
rect 576302 6168 576308 6180
rect 171100 6140 576308 6168
rect 171100 6128 171106 6140
rect 576302 6128 576308 6140
rect 576360 6128 576366 6180
rect 313090 5516 313096 5568
rect 313148 5556 313154 5568
rect 314654 5556 314660 5568
rect 313148 5528 314660 5556
rect 313148 5516 313154 5528
rect 314654 5516 314660 5528
rect 314712 5516 314718 5568
rect 376018 5516 376024 5568
rect 376076 5556 376082 5568
rect 378870 5556 378876 5568
rect 376076 5528 378876 5556
rect 376076 5516 376082 5528
rect 378870 5516 378876 5528
rect 378928 5516 378934 5568
rect 384298 5516 384304 5568
rect 384356 5556 384362 5568
rect 387150 5556 387156 5568
rect 384356 5528 387156 5556
rect 384356 5516 384362 5528
rect 387150 5516 387156 5528
rect 387208 5516 387214 5568
rect 114002 5312 114008 5364
rect 114060 5352 114066 5364
rect 134058 5352 134064 5364
rect 114060 5324 134064 5352
rect 114060 5312 114066 5324
rect 134058 5312 134064 5324
rect 134116 5312 134122 5364
rect 101030 5244 101036 5296
rect 101088 5284 101094 5296
rect 133230 5284 133236 5296
rect 101088 5256 133236 5284
rect 101088 5244 101094 5256
rect 133230 5244 133236 5256
rect 133288 5244 133294 5296
rect 136910 5244 136916 5296
rect 136968 5284 136974 5296
rect 154206 5284 154212 5296
rect 136968 5256 154212 5284
rect 136968 5244 136974 5256
rect 154206 5244 154212 5256
rect 154264 5244 154270 5296
rect 93946 5176 93952 5228
rect 94004 5216 94010 5228
rect 133138 5216 133144 5228
rect 94004 5188 133144 5216
rect 94004 5176 94010 5188
rect 133138 5176 133144 5188
rect 133196 5176 133202 5228
rect 137002 5176 137008 5228
rect 137060 5216 137066 5228
rect 157794 5216 157800 5228
rect 137060 5188 157800 5216
rect 137060 5176 137066 5188
rect 157794 5176 157800 5188
rect 157852 5176 157858 5228
rect 63218 5108 63224 5160
rect 63276 5148 63282 5160
rect 129918 5148 129924 5160
rect 63276 5120 129924 5148
rect 63276 5108 63282 5120
rect 129918 5108 129924 5120
rect 129976 5108 129982 5160
rect 138290 5108 138296 5160
rect 138348 5148 138354 5160
rect 169570 5148 169576 5160
rect 138348 5120 169576 5148
rect 138348 5108 138354 5120
rect 169570 5108 169576 5120
rect 169628 5108 169634 5160
rect 30098 5040 30104 5092
rect 30156 5080 30162 5092
rect 127802 5080 127808 5092
rect 30156 5052 127808 5080
rect 30156 5040 30162 5052
rect 127802 5040 127808 5052
rect 127860 5040 127866 5092
rect 136818 5040 136824 5092
rect 136876 5080 136882 5092
rect 148318 5080 148324 5092
rect 136876 5052 148324 5080
rect 136876 5040 136882 5052
rect 148318 5040 148324 5052
rect 148376 5040 148382 5092
rect 154390 5040 154396 5092
rect 154448 5080 154454 5092
rect 213086 5080 213092 5092
rect 154448 5052 213092 5080
rect 154448 5040 154454 5052
rect 213086 5040 213092 5052
rect 213144 5040 213150 5092
rect 15930 4972 15936 5024
rect 15988 5012 15994 5024
rect 113818 5012 113824 5024
rect 15988 4984 113824 5012
rect 15988 4972 15994 4984
rect 113818 4972 113824 4984
rect 113876 4972 113882 5024
rect 142154 4972 142160 5024
rect 142212 5012 142218 5024
rect 216858 5012 216864 5024
rect 142212 4984 216864 5012
rect 142212 4972 142218 4984
rect 216858 4972 216864 4984
rect 216916 4972 216922 5024
rect 436830 4972 436836 5024
rect 436888 5012 436894 5024
rect 436888 4984 451274 5012
rect 436888 4972 436894 4984
rect 28902 4904 28908 4956
rect 28960 4944 28966 4956
rect 127894 4944 127900 4956
rect 28960 4916 127900 4944
rect 28960 4904 28966 4916
rect 127894 4904 127900 4916
rect 127952 4904 127958 4956
rect 148686 4904 148692 4956
rect 148744 4944 148750 4956
rect 294874 4944 294880 4956
rect 148744 4916 294880 4944
rect 148744 4904 148750 4916
rect 294874 4904 294880 4916
rect 294932 4904 294938 4956
rect 451246 4944 451274 4984
rect 479334 4944 479340 4956
rect 451246 4916 479340 4944
rect 479334 4904 479340 4916
rect 479392 4904 479398 4956
rect 6454 4836 6460 4888
rect 6512 4876 6518 4888
rect 10318 4876 10324 4888
rect 6512 4848 10324 4876
rect 6512 4836 6518 4848
rect 10318 4836 10324 4848
rect 10376 4836 10382 4888
rect 13538 4836 13544 4888
rect 13596 4876 13602 4888
rect 125962 4876 125968 4888
rect 13596 4848 125968 4876
rect 13596 4836 13602 4848
rect 125962 4836 125968 4848
rect 126020 4836 126026 4888
rect 138198 4836 138204 4888
rect 138256 4876 138262 4888
rect 162486 4876 162492 4888
rect 138256 4848 162492 4876
rect 138256 4836 138262 4848
rect 162486 4836 162492 4848
rect 162544 4836 162550 4888
rect 162854 4836 162860 4888
rect 162912 4876 162918 4888
rect 487614 4876 487620 4888
rect 162912 4848 487620 4876
rect 162912 4836 162918 4848
rect 487614 4836 487620 4848
rect 487672 4836 487678 4888
rect 8754 4768 8760 4820
rect 8812 4808 8818 4820
rect 125870 4808 125876 4820
rect 8812 4780 125876 4808
rect 8812 4768 8818 4780
rect 125870 4768 125876 4780
rect 125928 4768 125934 4820
rect 138106 4768 138112 4820
rect 138164 4808 138170 4820
rect 166074 4808 166080 4820
rect 138164 4780 166080 4808
rect 138164 4768 138170 4780
rect 166074 4768 166080 4780
rect 166132 4768 166138 4820
rect 169478 4768 169484 4820
rect 169536 4808 169542 4820
rect 562042 4808 562048 4820
rect 169536 4780 562048 4808
rect 169536 4768 169542 4780
rect 562042 4768 562048 4780
rect 562100 4768 562106 4820
rect 136726 4428 136732 4480
rect 136784 4468 136790 4480
rect 144730 4468 144736 4480
rect 136784 4440 144736 4468
rect 136784 4428 136790 4440
rect 144730 4428 144736 4440
rect 144788 4428 144794 4480
rect 184934 4156 184940 4208
rect 184992 4196 184998 4208
rect 186130 4196 186136 4208
rect 184992 4168 186136 4196
rect 184992 4156 184998 4168
rect 186130 4156 186136 4168
rect 186188 4156 186194 4208
rect 201494 4156 201500 4208
rect 201552 4196 201558 4208
rect 202690 4196 202696 4208
rect 201552 4168 202696 4196
rect 201552 4156 201558 4168
rect 202690 4156 202696 4168
rect 202748 4156 202754 4208
rect 242894 4156 242900 4208
rect 242952 4196 242958 4208
rect 244090 4196 244096 4208
rect 242952 4168 244096 4196
rect 242952 4156 242958 4168
rect 244090 4156 244096 4168
rect 244148 4156 244154 4208
rect 251174 4156 251180 4208
rect 251232 4196 251238 4208
rect 252370 4196 252376 4208
rect 251232 4168 252376 4196
rect 251232 4156 251238 4168
rect 252370 4156 252376 4168
rect 252428 4156 252434 4208
rect 566 4088 572 4140
rect 624 4128 630 4140
rect 7558 4128 7564 4140
rect 624 4100 7564 4128
rect 624 4088 630 4100
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 11146 4088 11152 4140
rect 11204 4128 11210 4140
rect 126422 4128 126428 4140
rect 11204 4100 126428 4128
rect 11204 4088 11210 4100
rect 126422 4088 126428 4100
rect 126480 4088 126486 4140
rect 144362 4088 144368 4140
rect 144420 4128 144426 4140
rect 153010 4128 153016 4140
rect 144420 4100 153016 4128
rect 144420 4088 144426 4100
rect 153010 4088 153016 4100
rect 153068 4088 153074 4140
rect 172330 4088 172336 4140
rect 172388 4128 172394 4140
rect 288986 4128 288992 4140
rect 172388 4100 288992 4128
rect 172388 4088 172394 4100
rect 288986 4088 288992 4100
rect 289044 4088 289050 4140
rect 124858 4060 124864 4072
rect 122806 4032 124864 4060
rect 87966 3952 87972 4004
rect 88024 3992 88030 4004
rect 122806 3992 122834 4032
rect 124858 4020 124864 4032
rect 124916 4020 124922 4072
rect 125870 4020 125876 4072
rect 125928 4060 125934 4072
rect 134518 4060 134524 4072
rect 125928 4032 134524 4060
rect 125928 4020 125934 4032
rect 134518 4020 134524 4032
rect 134576 4020 134582 4072
rect 146478 4020 146484 4072
rect 146536 4060 146542 4072
rect 268838 4060 268844 4072
rect 146536 4032 268844 4060
rect 146536 4020 146542 4032
rect 268838 4020 268844 4032
rect 268896 4020 268902 4072
rect 88024 3964 122834 3992
rect 88024 3952 88030 3964
rect 124674 3952 124680 4004
rect 124732 3992 124738 4004
rect 134610 3992 134616 4004
rect 124732 3964 134616 3992
rect 124732 3952 124738 3964
rect 134610 3952 134616 3964
rect 134668 3952 134674 4004
rect 138934 3952 138940 4004
rect 138992 3992 138998 4004
rect 143534 3992 143540 4004
rect 138992 3964 143540 3992
rect 138992 3952 138998 3964
rect 143534 3952 143540 3964
rect 143592 3952 143598 4004
rect 146386 3952 146392 4004
rect 146444 3992 146450 4004
rect 272426 3992 272432 4004
rect 146444 3964 272432 3992
rect 146444 3952 146450 3964
rect 272426 3952 272432 3964
rect 272484 3952 272490 4004
rect 314654 3952 314660 4004
rect 314712 3992 314718 4004
rect 324406 3992 324412 4004
rect 314712 3964 324412 3992
rect 314712 3952 314718 3964
rect 324406 3952 324412 3964
rect 324464 3952 324470 4004
rect 86862 3884 86868 3936
rect 86920 3924 86926 3936
rect 131206 3924 131212 3936
rect 86920 3896 131212 3924
rect 86920 3884 86926 3896
rect 131206 3884 131212 3896
rect 131264 3884 131270 3936
rect 144454 3884 144460 3936
rect 144512 3924 144518 3936
rect 156598 3924 156604 3936
rect 144512 3896 156604 3924
rect 144512 3884 144518 3896
rect 156598 3884 156604 3896
rect 156656 3884 156662 3936
rect 163774 3884 163780 3936
rect 163832 3924 163838 3936
rect 303154 3924 303160 3936
rect 163832 3896 303160 3924
rect 163832 3884 163838 3896
rect 303154 3884 303160 3896
rect 303212 3884 303218 3936
rect 312538 3884 312544 3936
rect 312596 3924 312602 3936
rect 322106 3924 322112 3936
rect 312596 3896 322112 3924
rect 312596 3884 312602 3896
rect 322106 3884 322112 3896
rect 322164 3884 322170 3936
rect 83274 3816 83280 3868
rect 83332 3856 83338 3868
rect 131942 3856 131948 3868
rect 83332 3828 131948 3856
rect 83332 3816 83338 3828
rect 131942 3816 131948 3828
rect 132000 3816 132006 3868
rect 142798 3816 142804 3868
rect 142856 3856 142862 3868
rect 163682 3856 163688 3868
rect 142856 3828 163688 3856
rect 142856 3816 142862 3828
rect 163682 3816 163688 3828
rect 163740 3816 163746 3868
rect 173618 3816 173624 3868
rect 173676 3856 173682 3868
rect 212166 3856 212172 3868
rect 173676 3828 212172 3856
rect 173676 3816 173682 3828
rect 212166 3816 212172 3828
rect 212224 3816 212230 3868
rect 213086 3816 213092 3868
rect 213144 3856 213150 3868
rect 364610 3856 364616 3868
rect 213144 3828 364616 3856
rect 213144 3816 213150 3828
rect 364610 3816 364616 3828
rect 364668 3816 364674 3868
rect 367738 3816 367744 3868
rect 367796 3856 367802 3868
rect 377674 3856 377680 3868
rect 367796 3828 377680 3856
rect 367796 3816 367802 3828
rect 377674 3816 377680 3828
rect 377732 3816 377738 3868
rect 388438 3816 388444 3868
rect 388496 3856 388502 3868
rect 396534 3856 396540 3868
rect 388496 3828 396540 3856
rect 388496 3816 388502 3828
rect 396534 3816 396540 3828
rect 396592 3816 396598 3868
rect 398098 3816 398104 3868
rect 398156 3856 398162 3868
rect 408402 3856 408408 3868
rect 398156 3828 408408 3856
rect 398156 3816 398162 3828
rect 408402 3816 408408 3828
rect 408460 3816 408466 3868
rect 79686 3748 79692 3800
rect 79744 3788 79750 3800
rect 131298 3788 131304 3800
rect 79744 3760 131304 3788
rect 79744 3748 79750 3760
rect 131298 3748 131304 3760
rect 131356 3748 131362 3800
rect 140222 3748 140228 3800
rect 140280 3788 140286 3800
rect 164878 3788 164884 3800
rect 140280 3760 164884 3788
rect 140280 3748 140286 3760
rect 164878 3748 164884 3760
rect 164936 3748 164942 3800
rect 172422 3748 172428 3800
rect 172480 3788 172486 3800
rect 356330 3788 356336 3800
rect 172480 3760 356336 3788
rect 172480 3748 172486 3760
rect 356330 3748 356336 3760
rect 356388 3748 356394 3800
rect 359550 3748 359556 3800
rect 359608 3788 359614 3800
rect 368198 3788 368204 3800
rect 359608 3760 368204 3788
rect 359608 3748 359614 3760
rect 368198 3748 368204 3760
rect 368256 3748 368262 3800
rect 382918 3748 382924 3800
rect 382976 3788 382982 3800
rect 388254 3788 388260 3800
rect 382976 3760 388260 3788
rect 382976 3748 382982 3760
rect 388254 3748 388260 3760
rect 388312 3748 388318 3800
rect 388530 3748 388536 3800
rect 388588 3788 388594 3800
rect 398834 3788 398840 3800
rect 388588 3760 398840 3788
rect 388588 3748 388594 3760
rect 398834 3748 398840 3760
rect 398892 3748 398898 3800
rect 449158 3748 449164 3800
rect 449216 3788 449222 3800
rect 521838 3788 521844 3800
rect 449216 3760 521844 3788
rect 449216 3748 449222 3760
rect 521838 3748 521844 3760
rect 521896 3748 521902 3800
rect 69106 3680 69112 3732
rect 69164 3720 69170 3732
rect 126238 3720 126244 3732
rect 69164 3692 126244 3720
rect 69164 3680 69170 3692
rect 126238 3680 126244 3692
rect 126296 3680 126302 3732
rect 130654 3720 130660 3732
rect 126716 3692 130660 3720
rect 65518 3612 65524 3664
rect 65576 3652 65582 3664
rect 126716 3652 126744 3692
rect 130654 3680 130660 3692
rect 130712 3680 130718 3732
rect 142982 3680 142988 3732
rect 143040 3720 143046 3732
rect 155402 3720 155408 3732
rect 143040 3692 155408 3720
rect 143040 3680 143046 3692
rect 155402 3680 155408 3692
rect 155460 3680 155466 3732
rect 159818 3680 159824 3732
rect 159876 3720 159882 3732
rect 437934 3720 437940 3732
rect 159876 3692 437940 3720
rect 159876 3680 159882 3692
rect 437934 3680 437940 3692
rect 437992 3680 437998 3732
rect 449894 3680 449900 3732
rect 449952 3720 449958 3732
rect 525426 3720 525432 3732
rect 449952 3692 525432 3720
rect 449952 3680 449958 3692
rect 525426 3680 525432 3692
rect 525484 3680 525490 3732
rect 65576 3624 126744 3652
rect 65576 3612 65582 3624
rect 126974 3612 126980 3664
rect 127032 3652 127038 3664
rect 130286 3652 130292 3664
rect 127032 3624 130292 3652
rect 127032 3612 127038 3624
rect 130286 3612 130292 3624
rect 130344 3612 130350 3664
rect 140130 3612 140136 3664
rect 140188 3652 140194 3664
rect 170766 3652 170772 3664
rect 140188 3624 170772 3652
rect 140188 3612 140194 3624
rect 170766 3612 170772 3624
rect 170824 3612 170830 3664
rect 176654 3612 176660 3664
rect 176712 3652 176718 3664
rect 177850 3652 177856 3664
rect 176712 3624 177856 3652
rect 176712 3612 176718 3624
rect 177850 3612 177856 3624
rect 177908 3612 177914 3664
rect 177942 3612 177948 3664
rect 178000 3652 178006 3664
rect 461578 3652 461584 3664
rect 178000 3624 461584 3652
rect 178000 3612 178006 3624
rect 461578 3612 461584 3624
rect 461636 3612 461642 3664
rect 17034 3544 17040 3596
rect 17092 3584 17098 3596
rect 125778 3584 125784 3596
rect 17092 3556 125784 3584
rect 17092 3544 17098 3556
rect 125778 3544 125784 3556
rect 125836 3544 125842 3596
rect 129366 3544 129372 3596
rect 129424 3584 129430 3596
rect 130470 3584 130476 3596
rect 129424 3556 130476 3584
rect 129424 3544 129430 3556
rect 130470 3544 130476 3556
rect 130528 3544 130534 3596
rect 131758 3544 131764 3596
rect 131816 3584 131822 3596
rect 135806 3584 135812 3596
rect 131816 3556 135812 3584
rect 131816 3544 131822 3556
rect 135806 3544 135812 3556
rect 135864 3544 135870 3596
rect 138658 3544 138664 3596
rect 138716 3584 138722 3596
rect 151814 3584 151820 3596
rect 138716 3556 151820 3584
rect 138716 3544 138722 3556
rect 151814 3544 151820 3556
rect 151872 3544 151878 3596
rect 161658 3544 161664 3596
rect 161716 3584 161722 3596
rect 462774 3584 462780 3596
rect 161716 3556 462780 3584
rect 161716 3544 161722 3556
rect 462774 3544 462780 3556
rect 462832 3544 462838 3596
rect 481634 3544 481640 3596
rect 481692 3584 481698 3596
rect 482462 3584 482468 3596
rect 481692 3556 482468 3584
rect 481692 3544 481698 3556
rect 482462 3544 482468 3556
rect 482520 3544 482526 3596
rect 506474 3544 506480 3596
rect 506532 3584 506538 3596
rect 507302 3584 507308 3596
rect 506532 3556 507308 3584
rect 506532 3544 506538 3556
rect 507302 3544 507308 3556
rect 507360 3544 507366 3596
rect 518342 3584 518348 3596
rect 509206 3556 518348 3584
rect 12342 3476 12348 3528
rect 12400 3516 12406 3528
rect 126606 3516 126612 3528
rect 12400 3488 126612 3516
rect 12400 3476 12406 3488
rect 126606 3476 126612 3488
rect 126664 3476 126670 3528
rect 135254 3476 135260 3528
rect 135312 3516 135318 3528
rect 136542 3516 136548 3528
rect 135312 3488 136548 3516
rect 135312 3476 135318 3488
rect 136542 3476 136548 3488
rect 136600 3476 136606 3528
rect 162762 3476 162768 3528
rect 162820 3516 162826 3528
rect 466270 3516 466276 3528
rect 162820 3488 466276 3516
rect 162820 3476 162826 3488
rect 466270 3476 466276 3488
rect 466328 3476 466334 3528
rect 473998 3476 474004 3528
rect 474056 3516 474062 3528
rect 509206 3516 509234 3556
rect 518342 3544 518348 3556
rect 518400 3544 518406 3596
rect 574738 3544 574744 3596
rect 574796 3584 574802 3596
rect 574796 3556 576854 3584
rect 574796 3544 574802 3556
rect 474056 3488 509234 3516
rect 474056 3476 474062 3488
rect 514754 3476 514760 3528
rect 514812 3516 514818 3528
rect 515582 3516 515588 3528
rect 514812 3488 515588 3516
rect 514812 3476 514818 3488
rect 515582 3476 515588 3488
rect 515640 3476 515646 3528
rect 539594 3476 539600 3528
rect 539652 3516 539658 3528
rect 540422 3516 540428 3528
rect 539652 3488 540428 3516
rect 539652 3476 539658 3488
rect 540422 3476 540428 3488
rect 540480 3476 540486 3528
rect 564434 3476 564440 3528
rect 564492 3516 564498 3528
rect 565262 3516 565268 3528
rect 564492 3488 565268 3516
rect 564492 3476 564498 3488
rect 565262 3476 565268 3488
rect 565320 3476 565326 3528
rect 35894 3408 35900 3460
rect 35952 3448 35958 3460
rect 36814 3448 36820 3460
rect 35952 3420 36820 3448
rect 35952 3408 35958 3420
rect 36814 3408 36820 3420
rect 36872 3408 36878 3460
rect 118694 3408 118700 3460
rect 118752 3448 118758 3460
rect 119890 3448 119896 3460
rect 118752 3420 119896 3448
rect 118752 3408 118758 3420
rect 119890 3408 119896 3420
rect 119948 3408 119954 3460
rect 135898 3408 135904 3460
rect 135956 3448 135962 3460
rect 138842 3448 138848 3460
rect 135956 3420 138848 3448
rect 135956 3408 135962 3420
rect 138842 3408 138848 3420
rect 138900 3408 138906 3460
rect 139026 3408 139032 3460
rect 139084 3448 139090 3460
rect 168374 3448 168380 3460
rect 139084 3420 168380 3448
rect 139084 3408 139090 3420
rect 168374 3408 168380 3420
rect 168432 3408 168438 3460
rect 172054 3408 172060 3460
rect 172112 3448 172118 3460
rect 179046 3448 179052 3460
rect 172112 3420 179052 3448
rect 172112 3408 172118 3420
rect 179046 3408 179052 3420
rect 179104 3408 179110 3460
rect 181438 3448 181444 3460
rect 179156 3420 181444 3448
rect 135714 3340 135720 3392
rect 135772 3380 135778 3392
rect 141234 3380 141240 3392
rect 135772 3352 141240 3380
rect 135772 3340 135778 3352
rect 141234 3340 141240 3352
rect 141292 3340 141298 3392
rect 173250 3340 173256 3392
rect 173308 3380 173314 3392
rect 177942 3380 177948 3392
rect 173308 3352 177948 3380
rect 173308 3340 173314 3352
rect 177942 3340 177948 3352
rect 178000 3340 178006 3392
rect 137830 3272 137836 3324
rect 137888 3312 137894 3324
rect 150618 3312 150624 3324
rect 137888 3284 150624 3312
rect 137888 3272 137894 3284
rect 150618 3272 150624 3284
rect 150676 3272 150682 3324
rect 154482 3272 154488 3324
rect 154540 3312 154546 3324
rect 173158 3312 173164 3324
rect 154540 3284 173164 3312
rect 154540 3272 154546 3284
rect 173158 3272 173164 3284
rect 173216 3272 173222 3324
rect 173434 3272 173440 3324
rect 173492 3312 173498 3324
rect 179156 3312 179184 3420
rect 181438 3408 181444 3420
rect 181496 3408 181502 3460
rect 181530 3408 181536 3460
rect 181588 3448 181594 3460
rect 519538 3448 519544 3460
rect 181588 3420 519544 3448
rect 181588 3408 181594 3420
rect 519538 3408 519544 3420
rect 519596 3408 519602 3460
rect 576826 3448 576854 3556
rect 580994 3448 581000 3460
rect 576826 3420 581000 3448
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 285398 3380 285404 3392
rect 173492 3284 179184 3312
rect 179248 3352 285404 3380
rect 173492 3272 173498 3284
rect 132954 3136 132960 3188
rect 133012 3176 133018 3188
rect 135438 3176 135444 3188
rect 133012 3148 135444 3176
rect 133012 3136 133018 3148
rect 135438 3136 135444 3148
rect 135496 3136 135502 3188
rect 135530 3136 135536 3188
rect 135588 3176 135594 3188
rect 140038 3176 140044 3188
rect 135588 3148 140044 3176
rect 135588 3136 135594 3148
rect 140038 3136 140044 3148
rect 140096 3136 140102 3188
rect 171870 3136 171876 3188
rect 171928 3176 171934 3188
rect 179248 3176 179276 3352
rect 285398 3340 285404 3352
rect 285456 3340 285462 3392
rect 307754 3340 307760 3392
rect 307812 3380 307818 3392
rect 309042 3380 309048 3392
rect 307812 3352 309048 3380
rect 307812 3340 307818 3352
rect 309042 3340 309048 3352
rect 309100 3340 309106 3392
rect 316034 3340 316040 3392
rect 316092 3380 316098 3392
rect 317322 3380 317328 3392
rect 316092 3352 317328 3380
rect 316092 3340 316098 3352
rect 317322 3340 317328 3352
rect 317380 3340 317386 3392
rect 332686 3340 332692 3392
rect 332744 3380 332750 3392
rect 333882 3380 333888 3392
rect 332744 3352 333888 3380
rect 332744 3340 332750 3352
rect 333882 3340 333888 3352
rect 333940 3340 333946 3392
rect 340966 3340 340972 3392
rect 341024 3380 341030 3392
rect 342162 3380 342168 3392
rect 341024 3352 342168 3380
rect 341024 3340 341030 3352
rect 342162 3340 342168 3352
rect 342220 3340 342226 3392
rect 365806 3340 365812 3392
rect 365864 3380 365870 3392
rect 367002 3380 367008 3392
rect 365864 3352 367008 3380
rect 365864 3340 365870 3352
rect 367002 3340 367008 3352
rect 367060 3340 367066 3392
rect 374086 3340 374092 3392
rect 374144 3380 374150 3392
rect 375282 3380 375288 3392
rect 374144 3352 375288 3380
rect 374144 3340 374150 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 382366 3340 382372 3392
rect 382424 3380 382430 3392
rect 383562 3380 383568 3392
rect 382424 3352 383568 3380
rect 382424 3340 382430 3352
rect 383562 3340 383568 3352
rect 383620 3340 383626 3392
rect 398926 3340 398932 3392
rect 398984 3380 398990 3392
rect 400122 3380 400128 3392
rect 398984 3352 400128 3380
rect 398984 3340 398990 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 415486 3340 415492 3392
rect 415544 3380 415550 3392
rect 416682 3380 416688 3392
rect 415544 3352 416688 3380
rect 415544 3340 415550 3352
rect 416682 3340 416688 3352
rect 416740 3340 416746 3392
rect 423766 3340 423772 3392
rect 423824 3380 423830 3392
rect 424962 3380 424968 3392
rect 423824 3352 424968 3380
rect 423824 3340 423830 3352
rect 424962 3340 424968 3352
rect 425020 3340 425026 3392
rect 431954 3340 431960 3392
rect 432012 3380 432018 3392
rect 433242 3380 433248 3392
rect 432012 3352 433248 3380
rect 432012 3340 432018 3352
rect 433242 3340 433248 3352
rect 433300 3340 433306 3392
rect 440326 3340 440332 3392
rect 440384 3380 440390 3392
rect 441522 3380 441528 3392
rect 440384 3352 441528 3380
rect 440384 3340 440390 3352
rect 441522 3340 441528 3352
rect 441580 3340 441586 3392
rect 456794 3340 456800 3392
rect 456852 3380 456858 3392
rect 458082 3380 458088 3392
rect 456852 3352 458088 3380
rect 456852 3340 456858 3352
rect 458082 3340 458088 3352
rect 458140 3340 458146 3392
rect 322750 3272 322756 3324
rect 322808 3312 322814 3324
rect 325602 3312 325608 3324
rect 322808 3284 325608 3312
rect 322808 3272 322814 3284
rect 325602 3272 325608 3284
rect 325660 3272 325666 3324
rect 403710 3272 403716 3324
rect 403768 3312 403774 3324
rect 406010 3312 406016 3324
rect 403768 3284 406016 3312
rect 403768 3272 403774 3284
rect 406010 3272 406016 3284
rect 406068 3272 406074 3324
rect 395338 3204 395344 3256
rect 395396 3244 395402 3256
rect 401318 3244 401324 3256
rect 395396 3216 401324 3244
rect 395396 3204 395402 3216
rect 401318 3204 401324 3216
rect 401376 3204 401382 3256
rect 171928 3148 179276 3176
rect 171928 3136 171934 3148
rect 384390 3136 384396 3188
rect 384448 3176 384454 3188
rect 389450 3176 389456 3188
rect 384448 3148 389456 3176
rect 384448 3136 384454 3148
rect 389450 3136 389456 3148
rect 389508 3136 389514 3188
rect 173710 3068 173716 3120
rect 173768 3108 173774 3120
rect 182542 3108 182548 3120
rect 173768 3080 182548 3108
rect 173768 3068 173774 3080
rect 182542 3068 182548 3080
rect 182600 3068 182606 3120
rect 326430 3068 326436 3120
rect 326488 3108 326494 3120
rect 331582 3108 331588 3120
rect 326488 3080 331588 3108
rect 326488 3068 326494 3080
rect 331582 3068 331588 3080
rect 331640 3068 331646 3120
rect 135622 3000 135628 3052
rect 135680 3040 135686 3052
rect 137646 3040 137652 3052
rect 135680 3012 137652 3040
rect 135680 3000 135686 3012
rect 137646 3000 137652 3012
rect 137704 3000 137710 3052
rect 378042 3000 378048 3052
rect 378100 3040 378106 3052
rect 382366 3040 382372 3052
rect 378100 3012 382372 3040
rect 378100 3000 378106 3012
rect 382366 3000 382372 3012
rect 382424 3000 382430 3052
rect 165062 2932 165068 2984
rect 165120 2972 165126 2984
rect 171962 2972 171968 2984
rect 165120 2944 171968 2972
rect 165120 2932 165126 2944
rect 171962 2932 171968 2944
rect 172020 2932 172026 2984
rect 327074 2932 327080 2984
rect 327132 2972 327138 2984
rect 335078 2972 335084 2984
rect 327132 2944 335084 2972
rect 327132 2932 327138 2944
rect 335078 2932 335084 2944
rect 335136 2932 335142 2984
rect 357434 2456 357440 2508
rect 357492 2496 357498 2508
rect 358722 2496 358728 2508
rect 357492 2468 358728 2496
rect 357492 2456 357498 2468
rect 358722 2456 358728 2468
rect 358780 2456 358786 2508
rect 349154 1232 349160 1284
rect 349212 1272 349218 1284
rect 350442 1272 350448 1284
rect 349212 1244 350448 1272
rect 349212 1232 349218 1244
rect 350442 1232 350448 1244
rect 350500 1232 350506 1284
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 196624 700612 196676 700664
rect 218980 700612 219032 700664
rect 193864 700544 193916 700596
rect 283840 700544 283892 700596
rect 192484 700476 192536 700528
rect 348792 700476 348844 700528
rect 189724 700408 189776 700460
rect 413652 700408 413704 700460
rect 188344 700340 188396 700392
rect 478512 700340 478564 700392
rect 89168 700272 89220 700324
rect 180800 700272 180852 700324
rect 185584 700272 185636 700324
rect 543464 700272 543516 700324
rect 105452 699660 105504 699712
rect 106924 699660 106976 699712
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 2780 683680 2832 683732
rect 4804 683680 4856 683732
rect 184204 683136 184256 683188
rect 579620 683136 579672 683188
rect 3516 670692 3568 670744
rect 180892 670692 180944 670744
rect 182824 643084 182876 643136
rect 580172 643084 580224 643136
rect 3516 632068 3568 632120
rect 7564 632068 7616 632120
rect 184296 630640 184348 630692
rect 579712 630640 579764 630692
rect 3516 618264 3568 618316
rect 180984 618264 181036 618316
rect 120724 616836 120776 616888
rect 580172 616836 580224 616888
rect 3516 579640 3568 579692
rect 17224 579640 17276 579692
rect 184388 576852 184440 576904
rect 580172 576852 580224 576904
rect 3056 565836 3108 565888
rect 179420 565836 179472 565888
rect 120816 563048 120868 563100
rect 580172 563048 580224 563100
rect 180064 536800 180116 536852
rect 580172 536800 580224 536852
rect 3516 527824 3568 527876
rect 8944 527824 8996 527876
rect 214564 524424 214616 524476
rect 579804 524424 579856 524476
rect 3516 514768 3568 514820
rect 181076 514768 181128 514820
rect 120908 510620 120960 510672
rect 579988 510620 580040 510672
rect 182916 484372 182968 484424
rect 580172 484372 580224 484424
rect 3516 474716 3568 474768
rect 10324 474716 10376 474768
rect 211804 470568 211856 470620
rect 579620 470568 579672 470620
rect 121000 456764 121052 456816
rect 579620 456764 579672 456816
rect 118700 431196 118752 431248
rect 580540 431196 580592 431248
rect 2964 422288 3016 422340
rect 13084 422288 13136 422340
rect 183008 418140 183060 418192
rect 580172 418140 580224 418192
rect 3056 409844 3108 409896
rect 179512 409844 179564 409896
rect 118608 404336 118660 404388
rect 580172 404336 580224 404388
rect 3332 371220 3384 371272
rect 84844 371220 84896 371272
rect 224224 364352 224276 364404
rect 580172 364352 580224 364404
rect 3332 357416 3384 357468
rect 181168 357416 181220 357468
rect 118516 351908 118568 351960
rect 580172 351908 580224 351960
rect 3332 318792 3384 318844
rect 14464 318792 14516 318844
rect 221464 311856 221516 311908
rect 580172 311856 580224 311908
rect 3332 304988 3384 305040
rect 182180 304988 182232 305040
rect 146944 298120 146996 298172
rect 580172 298120 580224 298172
rect 183100 271872 183152 271924
rect 580172 271872 580224 271924
rect 3332 266364 3384 266416
rect 18604 266364 18656 266416
rect 220084 258068 220136 258120
rect 579620 258068 579672 258120
rect 3332 253920 3384 253972
rect 178684 253920 178736 253972
rect 126244 244264 126296 244316
rect 580172 244264 580224 244316
rect 3332 240116 3384 240168
rect 82084 240116 82136 240168
rect 217324 218016 217376 218068
rect 580172 218016 580224 218068
rect 3332 213936 3384 213988
rect 31024 213936 31076 213988
rect 122104 205640 122156 205692
rect 580172 205640 580224 205692
rect 3332 201492 3384 201544
rect 178776 201492 178828 201544
rect 3332 187688 3384 187740
rect 119344 187688 119396 187740
rect 215944 178032 215996 178084
rect 580172 178032 580224 178084
rect 3516 166268 3568 166320
rect 179696 166268 179748 166320
rect 122196 165588 122248 165640
rect 580172 165588 580224 165640
rect 3516 162868 3568 162920
rect 21364 162868 21416 162920
rect 183192 151784 183244 151836
rect 579988 151784 580040 151836
rect 3516 149064 3568 149116
rect 179604 149064 179656 149116
rect 119068 145596 119120 145648
rect 234620 145596 234672 145648
rect 23480 145528 23532 145580
rect 179788 145528 179840 145580
rect 119160 144168 119212 144220
rect 299480 144168 299532 144220
rect 118240 142876 118292 142928
rect 146944 142876 146996 142928
rect 153200 142876 153252 142928
rect 181444 142876 181496 142928
rect 118976 142808 119028 142860
rect 429200 142808 429252 142860
rect 118148 141516 118200 141568
rect 126244 141516 126296 141568
rect 136640 141516 136692 141568
rect 181352 141516 181404 141568
rect 118056 141448 118108 141500
rect 169760 141448 169812 141500
rect 118884 141380 118936 141432
rect 494060 141380 494112 141432
rect 119252 140088 119304 140140
rect 364340 140088 364392 140140
rect 118792 140020 118844 140072
rect 558920 140020 558972 140072
rect 118332 139544 118384 139596
rect 122104 139544 122156 139596
rect 118424 139476 118476 139528
rect 122196 139476 122248 139528
rect 3332 139408 3384 139460
rect 181536 139408 181588 139460
rect 178684 139340 178736 139392
rect 182272 139340 182324 139392
rect 178776 139272 178828 139324
rect 182364 139272 182416 139324
rect 196716 137980 196768 138032
rect 580172 137980 580224 138032
rect 3516 137776 3568 137828
rect 121092 137776 121144 137828
rect 7656 136688 7708 136740
rect 117320 136688 117372 136740
rect 9036 135260 9088 135312
rect 117320 135260 117372 135312
rect 3424 135056 3476 135108
rect 3424 134852 3476 134904
rect 22744 133900 22796 133952
rect 117320 133900 117372 133952
rect 21364 133832 21416 133884
rect 117412 133832 117464 133884
rect 31024 132404 31076 132456
rect 117320 132404 117372 132456
rect 18604 131044 18656 131096
rect 117320 131044 117372 131096
rect 14464 129684 14516 129736
rect 117320 129684 117372 129736
rect 84844 128256 84896 128308
rect 117320 128256 117372 128308
rect 13084 126896 13136 126948
rect 117320 126896 117372 126948
rect 10324 124108 10376 124160
rect 117320 124108 117372 124160
rect 8944 122748 8996 122800
rect 117320 122748 117372 122800
rect 17224 121388 17276 121440
rect 117320 121388 117372 121440
rect 7564 120028 7616 120080
rect 117320 120028 117372 120080
rect 4804 118600 4856 118652
rect 117320 118600 117372 118652
rect 40040 117240 40092 117292
rect 117320 117240 117372 117292
rect 106924 115880 106976 115932
rect 117320 115880 117372 115932
rect 180156 111800 180208 111852
rect 579988 111800 580040 111852
rect 3332 111732 3384 111784
rect 22744 111732 22796 111784
rect 183468 108944 183520 108996
rect 196624 108944 196676 108996
rect 183468 107584 183520 107636
rect 193864 107584 193916 107636
rect 183468 106224 183520 106276
rect 192484 106224 192536 106276
rect 182732 104796 182784 104848
rect 189724 104796 189776 104848
rect 183468 102620 183520 102672
rect 188344 102620 188396 102672
rect 182272 101464 182324 101516
rect 185584 101464 185636 101516
rect 182456 99968 182508 100020
rect 184204 99968 184256 100020
rect 193864 99356 193916 99408
rect 580172 99356 580224 99408
rect 182180 98472 182232 98524
rect 184296 98472 184348 98524
rect 182548 97384 182600 97436
rect 184388 97384 184440 97436
rect 183468 96568 183520 96620
rect 214564 96568 214616 96620
rect 183468 95140 183520 95192
rect 211804 95140 211856 95192
rect 182548 93100 182600 93152
rect 224224 93100 224276 93152
rect 183468 91740 183520 91792
rect 221464 91740 221516 91792
rect 183376 90312 183428 90364
rect 220084 90312 220136 90364
rect 580172 89088 580224 89140
rect 580632 89088 580684 89140
rect 183468 88952 183520 89004
rect 217324 88952 217376 89004
rect 580632 88952 580684 89004
rect 580908 88952 580960 89004
rect 183376 87592 183428 87644
rect 215944 87592 215996 87644
rect 183468 85484 183520 85536
rect 196716 85484 196768 85536
rect 3516 84192 3568 84244
rect 120724 84192 120776 84244
rect 183468 84124 183520 84176
rect 193864 84124 193916 84176
rect 120908 80792 120960 80844
rect 122104 80588 122156 80640
rect 6920 79976 6972 80028
rect 122104 79976 122156 80028
rect 125232 79908 125284 79960
rect 125830 79908 125882 79960
rect 126566 79908 126618 79960
rect 126658 79908 126710 79960
rect 126934 79908 126986 79960
rect 127026 79908 127078 79960
rect 127394 79908 127446 79960
rect 127486 79908 127538 79960
rect 126014 79840 126066 79892
rect 125876 79772 125928 79824
rect 126106 79772 126158 79824
rect 82084 79704 82136 79756
rect 120908 79704 120960 79756
rect 125968 79704 126020 79756
rect 3700 79568 3752 79620
rect 125140 79636 125192 79688
rect 125784 79568 125836 79620
rect 126750 79772 126802 79824
rect 126888 79772 126940 79824
rect 126980 79772 127032 79824
rect 126796 79636 126848 79688
rect 126704 79568 126756 79620
rect 127348 79568 127400 79620
rect 127670 79908 127722 79960
rect 127762 79908 127814 79960
rect 127854 79908 127906 79960
rect 127808 79772 127860 79824
rect 127900 79704 127952 79756
rect 126612 79500 126664 79552
rect 127440 79500 127492 79552
rect 127624 79500 127676 79552
rect 128314 79908 128366 79960
rect 128406 79908 128458 79960
rect 129050 79908 129102 79960
rect 129142 79908 129194 79960
rect 129418 79908 129470 79960
rect 128222 79840 128274 79892
rect 128590 79772 128642 79824
rect 128360 79704 128412 79756
rect 129004 79704 129056 79756
rect 128636 79636 128688 79688
rect 128820 79636 128872 79688
rect 129234 79840 129286 79892
rect 129464 79636 129516 79688
rect 129372 79568 129424 79620
rect 129786 79908 129838 79960
rect 129740 79636 129792 79688
rect 130246 79908 130298 79960
rect 129970 79840 130022 79892
rect 130062 79840 130114 79892
rect 130154 79840 130206 79892
rect 130016 79636 130068 79688
rect 130108 79568 130160 79620
rect 130200 79568 130252 79620
rect 128084 79432 128136 79484
rect 128176 79432 128228 79484
rect 128912 79432 128964 79484
rect 130522 79908 130574 79960
rect 130798 79908 130850 79960
rect 130890 79908 130942 79960
rect 131166 79908 131218 79960
rect 131258 79908 131310 79960
rect 131442 79908 131494 79960
rect 131534 79908 131586 79960
rect 131994 79908 132046 79960
rect 130614 79840 130666 79892
rect 130476 79636 130528 79688
rect 130982 79840 131034 79892
rect 130936 79704 130988 79756
rect 130568 79500 130620 79552
rect 130752 79500 130804 79552
rect 131120 79636 131172 79688
rect 3884 79296 3936 79348
rect 124404 79296 124456 79348
rect 127716 79296 127768 79348
rect 128544 79364 128596 79416
rect 130936 79432 130988 79484
rect 131442 79772 131494 79824
rect 131810 79772 131862 79824
rect 131902 79772 131954 79824
rect 131396 79568 131448 79620
rect 131672 79568 131724 79620
rect 131764 79568 131816 79620
rect 131580 79500 131632 79552
rect 131672 79432 131724 79484
rect 132178 79908 132230 79960
rect 132270 79840 132322 79892
rect 132040 79636 132092 79688
rect 132316 79704 132368 79756
rect 132914 79908 132966 79960
rect 133006 79908 133058 79960
rect 132638 79840 132690 79892
rect 133374 79908 133426 79960
rect 133466 79908 133518 79960
rect 133558 79908 133610 79960
rect 133834 79908 133886 79960
rect 134110 79908 134162 79960
rect 134202 79908 134254 79960
rect 132500 79636 132552 79688
rect 132224 79500 132276 79552
rect 133282 79840 133334 79892
rect 132730 79772 132782 79824
rect 132960 79772 133012 79824
rect 133512 79772 133564 79824
rect 133420 79704 133472 79756
rect 132684 79636 132736 79688
rect 133328 79636 133380 79688
rect 132776 79568 132828 79620
rect 133926 79840 133978 79892
rect 133788 79568 133840 79620
rect 134064 79568 134116 79620
rect 135122 79908 135174 79960
rect 135214 79908 135266 79960
rect 135306 79908 135358 79960
rect 135398 79908 135450 79960
rect 136042 79908 136094 79960
rect 136134 79908 136186 79960
rect 134846 79840 134898 79892
rect 134892 79704 134944 79756
rect 135582 79840 135634 79892
rect 135766 79840 135818 79892
rect 135352 79772 135404 79824
rect 134984 79636 135036 79688
rect 135168 79636 135220 79688
rect 135674 79772 135726 79824
rect 135812 79704 135864 79756
rect 134524 79568 134576 79620
rect 135260 79568 135312 79620
rect 135720 79636 135772 79688
rect 135536 79568 135588 79620
rect 135904 79636 135956 79688
rect 135996 79636 136048 79688
rect 136088 79568 136140 79620
rect 136318 79908 136370 79960
rect 136686 79908 136738 79960
rect 136778 79908 136830 79960
rect 137054 79908 137106 79960
rect 137146 79908 137198 79960
rect 137238 79908 137290 79960
rect 137330 79908 137382 79960
rect 137422 79908 137474 79960
rect 137606 79908 137658 79960
rect 133144 79500 133196 79552
rect 134156 79500 134208 79552
rect 135904 79500 135956 79552
rect 136870 79840 136922 79892
rect 136732 79772 136784 79824
rect 136916 79636 136968 79688
rect 136824 79568 136876 79620
rect 137376 79704 137428 79756
rect 137100 79568 137152 79620
rect 137192 79568 137244 79620
rect 137008 79500 137060 79552
rect 137468 79500 137520 79552
rect 137882 79908 137934 79960
rect 137698 79840 137750 79892
rect 137790 79840 137842 79892
rect 137928 79772 137980 79824
rect 137744 79636 137796 79688
rect 135628 79432 135680 79484
rect 136180 79432 136232 79484
rect 129924 79364 129976 79416
rect 135536 79364 135588 79416
rect 136180 79296 136232 79348
rect 138342 79908 138394 79960
rect 138802 79908 138854 79960
rect 138894 79908 138946 79960
rect 138986 79908 139038 79960
rect 139354 79908 139406 79960
rect 139538 79908 139590 79960
rect 138250 79840 138302 79892
rect 138112 79636 138164 79688
rect 138710 79840 138762 79892
rect 138526 79772 138578 79824
rect 138664 79704 138716 79756
rect 138480 79568 138532 79620
rect 138572 79500 138624 79552
rect 139262 79840 139314 79892
rect 139124 79636 139176 79688
rect 139492 79772 139544 79824
rect 139722 79908 139774 79960
rect 139814 79908 139866 79960
rect 140182 79908 140234 79960
rect 139400 79636 139452 79688
rect 139584 79636 139636 79688
rect 139308 79568 139360 79620
rect 140274 79840 140326 79892
rect 140366 79840 140418 79892
rect 140228 79636 140280 79688
rect 140044 79568 140096 79620
rect 139124 79500 139176 79552
rect 138388 79432 138440 79484
rect 140320 79500 140372 79552
rect 140642 79908 140694 79960
rect 141010 79908 141062 79960
rect 141746 79908 141798 79960
rect 141838 79908 141890 79960
rect 141930 79908 141982 79960
rect 142390 79908 142442 79960
rect 140826 79840 140878 79892
rect 141194 79840 141246 79892
rect 141562 79840 141614 79892
rect 140964 79772 141016 79824
rect 140780 79704 140832 79756
rect 140872 79704 140924 79756
rect 140596 79636 140648 79688
rect 141332 79500 141384 79552
rect 141792 79772 141844 79824
rect 141700 79568 141752 79620
rect 141976 79568 142028 79620
rect 142160 79568 142212 79620
rect 142482 79840 142534 79892
rect 143126 79908 143178 79960
rect 142942 79840 142994 79892
rect 142436 79500 142488 79552
rect 142620 79500 142672 79552
rect 143310 79908 143362 79960
rect 143494 79908 143546 79960
rect 143862 79908 143914 79960
rect 143172 79772 143224 79824
rect 143586 79840 143638 79892
rect 144046 79908 144098 79960
rect 144230 79908 144282 79960
rect 144322 79908 144374 79960
rect 144506 79908 144558 79960
rect 144690 79908 144742 79960
rect 144782 79908 144834 79960
rect 143356 79772 143408 79824
rect 143678 79772 143730 79824
rect 143080 79636 143132 79688
rect 143264 79500 143316 79552
rect 143540 79568 143592 79620
rect 144000 79500 144052 79552
rect 144276 79772 144328 79824
rect 144506 79772 144558 79824
rect 144460 79568 144512 79620
rect 145426 79908 145478 79960
rect 145518 79908 145570 79960
rect 145702 79908 145754 79960
rect 145794 79908 145846 79960
rect 146530 79908 146582 79960
rect 146622 79908 146674 79960
rect 144966 79840 145018 79892
rect 145150 79840 145202 79892
rect 144920 79704 144972 79756
rect 145334 79840 145386 79892
rect 145564 79704 145616 79756
rect 145656 79704 145708 79756
rect 145012 79636 145064 79688
rect 145196 79636 145248 79688
rect 145380 79636 145432 79688
rect 145978 79840 146030 79892
rect 146438 79772 146490 79824
rect 145840 79636 145892 79688
rect 145932 79636 145984 79688
rect 146714 79840 146766 79892
rect 146484 79636 146536 79688
rect 146898 79908 146950 79960
rect 147358 79908 147410 79960
rect 146760 79636 146812 79688
rect 146392 79568 146444 79620
rect 146576 79568 146628 79620
rect 146668 79568 146720 79620
rect 147174 79840 147226 79892
rect 147266 79840 147318 79892
rect 147726 79840 147778 79892
rect 147128 79568 147180 79620
rect 146208 79500 146260 79552
rect 147036 79500 147088 79552
rect 147910 79772 147962 79824
rect 148002 79772 148054 79824
rect 148094 79772 148146 79824
rect 147496 79568 147548 79620
rect 147588 79568 147640 79620
rect 147772 79500 147824 79552
rect 148048 79568 148100 79620
rect 143172 79432 143224 79484
rect 147864 79432 147916 79484
rect 148370 79840 148422 79892
rect 148554 79840 148606 79892
rect 148692 79636 148744 79688
rect 149014 79908 149066 79960
rect 150302 79908 150354 79960
rect 150578 79908 150630 79960
rect 150762 79908 150814 79960
rect 150854 79908 150906 79960
rect 150946 79908 150998 79960
rect 151222 79908 151274 79960
rect 151498 79908 151550 79960
rect 149382 79840 149434 79892
rect 149474 79840 149526 79892
rect 149842 79840 149894 79892
rect 149934 79840 149986 79892
rect 149106 79772 149158 79824
rect 148600 79568 148652 79620
rect 148968 79568 149020 79620
rect 149060 79568 149112 79620
rect 149152 79568 149204 79620
rect 148416 79500 148468 79552
rect 149520 79636 149572 79688
rect 149336 79568 149388 79620
rect 150026 79772 150078 79824
rect 150164 79636 150216 79688
rect 150394 79840 150446 79892
rect 150440 79704 150492 79756
rect 150670 79840 150722 79892
rect 150532 79636 150584 79688
rect 150256 79568 150308 79620
rect 149612 79500 149664 79552
rect 149980 79500 150032 79552
rect 150348 79500 150400 79552
rect 150854 79772 150906 79824
rect 150992 79568 151044 79620
rect 150808 79500 150860 79552
rect 151314 79840 151366 79892
rect 151406 79840 151458 79892
rect 151866 79908 151918 79960
rect 151958 79908 152010 79960
rect 152510 79908 152562 79960
rect 152694 79908 152746 79960
rect 151452 79636 151504 79688
rect 151544 79636 151596 79688
rect 151728 79636 151780 79688
rect 151268 79568 151320 79620
rect 151360 79568 151412 79620
rect 152234 79840 152286 79892
rect 152142 79772 152194 79824
rect 152004 79636 152056 79688
rect 152096 79636 152148 79688
rect 152602 79840 152654 79892
rect 152556 79704 152608 79756
rect 151912 79568 151964 79620
rect 152970 79908 153022 79960
rect 153154 79908 153206 79960
rect 153246 79908 153298 79960
rect 153338 79908 153390 79960
rect 153430 79908 153482 79960
rect 153016 79704 153068 79756
rect 153108 79704 153160 79756
rect 153200 79704 153252 79756
rect 153292 79636 153344 79688
rect 152556 79500 152608 79552
rect 152832 79500 152884 79552
rect 152924 79500 152976 79552
rect 153568 79500 153620 79552
rect 580356 80792 580408 80844
rect 178592 80724 178644 80776
rect 580724 80724 580776 80776
rect 174728 80588 174780 80640
rect 174820 80588 174872 80640
rect 175004 80588 175056 80640
rect 580816 80656 580868 80708
rect 176108 80452 176160 80504
rect 181352 80452 181404 80504
rect 174452 80384 174504 80436
rect 174912 80316 174964 80368
rect 154074 79908 154126 79960
rect 154626 79908 154678 79960
rect 156006 79908 156058 79960
rect 156190 79908 156242 79960
rect 154902 79840 154954 79892
rect 154442 79772 154494 79824
rect 155086 79772 155138 79824
rect 155270 79772 155322 79824
rect 155362 79772 155414 79824
rect 155454 79772 155506 79824
rect 154120 79704 154172 79756
rect 154212 79636 154264 79688
rect 155040 79636 155092 79688
rect 155408 79636 155460 79688
rect 154212 79500 154264 79552
rect 154856 79568 154908 79620
rect 155316 79568 155368 79620
rect 155500 79568 155552 79620
rect 155822 79840 155874 79892
rect 156052 79772 156104 79824
rect 156374 79772 156426 79824
rect 156144 79704 156196 79756
rect 155868 79636 155920 79688
rect 155684 79500 155736 79552
rect 156328 79500 156380 79552
rect 156742 79908 156794 79960
rect 156834 79908 156886 79960
rect 157202 79908 157254 79960
rect 157294 79908 157346 79960
rect 157386 79908 157438 79960
rect 157156 79772 157208 79824
rect 156880 79704 156932 79756
rect 157478 79840 157530 79892
rect 156788 79636 156840 79688
rect 157248 79636 157300 79688
rect 156696 79568 156748 79620
rect 157570 79772 157622 79824
rect 157524 79636 157576 79688
rect 158030 79908 158082 79960
rect 158122 79908 158174 79960
rect 158076 79704 158128 79756
rect 157616 79568 157668 79620
rect 157984 79568 158036 79620
rect 156788 79500 156840 79552
rect 157800 79500 157852 79552
rect 158260 79568 158312 79620
rect 174544 80248 174596 80300
rect 176384 80248 176436 80300
rect 200120 80248 200172 80300
rect 174636 80180 174688 80232
rect 231860 80180 231912 80232
rect 158858 79908 158910 79960
rect 159042 79908 159094 79960
rect 159318 79908 159370 79960
rect 160054 79908 160106 79960
rect 160146 79908 160198 79960
rect 160422 79908 160474 79960
rect 160606 79908 160658 79960
rect 160790 79908 160842 79960
rect 160882 79908 160934 79960
rect 161526 79908 161578 79960
rect 161894 79908 161946 79960
rect 162446 79908 162498 79960
rect 158582 79840 158634 79892
rect 158536 79636 158588 79688
rect 158766 79840 158818 79892
rect 159226 79840 159278 79892
rect 158904 79772 158956 79824
rect 158628 79568 158680 79620
rect 139952 79364 140004 79416
rect 152648 79364 152700 79416
rect 153476 79364 153528 79416
rect 153660 79364 153712 79416
rect 144552 79296 144604 79348
rect 155132 79364 155184 79416
rect 158168 79364 158220 79416
rect 158352 79364 158404 79416
rect 159502 79840 159554 79892
rect 159594 79840 159646 79892
rect 159456 79636 159508 79688
rect 159916 79636 159968 79688
rect 160330 79840 160382 79892
rect 160146 79772 160198 79824
rect 159456 79500 159508 79552
rect 160008 79500 160060 79552
rect 159732 79364 159784 79416
rect 160008 79364 160060 79416
rect 160468 79636 160520 79688
rect 160882 79772 160934 79824
rect 160744 79636 160796 79688
rect 161158 79840 161210 79892
rect 161250 79840 161302 79892
rect 161342 79840 161394 79892
rect 161112 79704 161164 79756
rect 161204 79636 161256 79688
rect 161710 79840 161762 79892
rect 161526 79772 161578 79824
rect 161572 79636 161624 79688
rect 161986 79840 162038 79892
rect 161940 79704 161992 79756
rect 162032 79636 162084 79688
rect 162354 79840 162406 79892
rect 162308 79704 162360 79756
rect 162400 79636 162452 79688
rect 162492 79636 162544 79688
rect 161756 79568 161808 79620
rect 162308 79568 162360 79620
rect 160928 79500 160980 79552
rect 162584 79500 162636 79552
rect 163090 79908 163142 79960
rect 164194 79908 164246 79960
rect 164286 79908 164338 79960
rect 164838 79908 164890 79960
rect 164930 79908 164982 79960
rect 162998 79840 163050 79892
rect 163458 79840 163510 79892
rect 163550 79840 163602 79892
rect 163734 79840 163786 79892
rect 162860 79568 162912 79620
rect 163688 79704 163740 79756
rect 162952 79500 163004 79552
rect 163044 79500 163096 79552
rect 163228 79500 163280 79552
rect 160836 79432 160888 79484
rect 160560 79364 160612 79416
rect 161388 79364 161440 79416
rect 161572 79364 161624 79416
rect 162308 79364 162360 79416
rect 120724 79228 120776 79280
rect 162676 79296 162728 79348
rect 163044 79364 163096 79416
rect 163504 79364 163556 79416
rect 164010 79840 164062 79892
rect 164148 79636 164200 79688
rect 164470 79840 164522 79892
rect 164608 79568 164660 79620
rect 164976 79636 165028 79688
rect 164516 79500 164568 79552
rect 164792 79500 164844 79552
rect 165666 79908 165718 79960
rect 165758 79908 165810 79960
rect 166494 79908 166546 79960
rect 166862 79908 166914 79960
rect 168426 79908 168478 79960
rect 168610 79908 168662 79960
rect 168794 79908 168846 79960
rect 165390 79840 165442 79892
rect 165482 79840 165534 79892
rect 165574 79840 165626 79892
rect 165436 79704 165488 79756
rect 165528 79636 165580 79688
rect 165252 79568 165304 79620
rect 165620 79568 165672 79620
rect 165436 79500 165488 79552
rect 166126 79772 166178 79824
rect 166218 79772 166270 79824
rect 166448 79704 166500 79756
rect 167690 79840 167742 79892
rect 167966 79840 168018 79892
rect 167874 79772 167926 79824
rect 168058 79772 168110 79824
rect 167920 79636 167972 79688
rect 168518 79840 168570 79892
rect 168380 79704 168432 79756
rect 168104 79636 168156 79688
rect 168472 79636 168524 79688
rect 169254 79840 169306 79892
rect 169162 79772 169214 79824
rect 166264 79568 166316 79620
rect 166356 79568 166408 79620
rect 166540 79568 166592 79620
rect 166816 79568 166868 79620
rect 167092 79568 167144 79620
rect 167644 79568 167696 79620
rect 167736 79568 167788 79620
rect 167828 79568 167880 79620
rect 168564 79568 168616 79620
rect 169300 79636 169352 79688
rect 169898 79908 169950 79960
rect 169990 79908 170042 79960
rect 170266 79908 170318 79960
rect 169806 79840 169858 79892
rect 169760 79704 169812 79756
rect 170174 79840 170226 79892
rect 169944 79636 169996 79688
rect 169208 79568 169260 79620
rect 169576 79568 169628 79620
rect 169852 79568 169904 79620
rect 170128 79704 170180 79756
rect 172014 79908 172066 79960
rect 174820 80112 174872 80164
rect 174912 80112 174964 80164
rect 252560 80112 252612 80164
rect 175464 80044 175516 80096
rect 175556 80044 175608 80096
rect 430580 80044 430632 80096
rect 172382 79908 172434 79960
rect 170542 79840 170594 79892
rect 178592 79976 178644 80028
rect 172658 79908 172710 79960
rect 172750 79908 172802 79960
rect 172934 79908 172986 79960
rect 173118 79908 173170 79960
rect 170220 79636 170272 79688
rect 170404 79636 170456 79688
rect 170312 79568 170364 79620
rect 170726 79772 170778 79824
rect 171094 79772 171146 79824
rect 171462 79772 171514 79824
rect 171324 79704 171376 79756
rect 171140 79636 171192 79688
rect 171232 79636 171284 79688
rect 172152 79636 172204 79688
rect 172612 79636 172664 79688
rect 171324 79568 171376 79620
rect 172336 79568 172388 79620
rect 173302 79840 173354 79892
rect 172888 79704 172940 79756
rect 173256 79704 173308 79756
rect 173578 79908 173630 79960
rect 173670 79908 173722 79960
rect 173762 79908 173814 79960
rect 173854 79908 173906 79960
rect 174728 79908 174780 79960
rect 174544 79840 174596 79892
rect 175556 79840 175608 79892
rect 173808 79772 173860 79824
rect 173624 79704 173676 79756
rect 173716 79704 173768 79756
rect 173440 79636 173492 79688
rect 201500 79568 201552 79620
rect 165988 79500 166040 79552
rect 166172 79500 166224 79552
rect 164424 79432 164476 79484
rect 171876 79500 171928 79552
rect 172428 79500 172480 79552
rect 180064 79500 180116 79552
rect 164056 79364 164108 79416
rect 167368 79432 167420 79484
rect 171784 79432 171836 79484
rect 172244 79432 172296 79484
rect 527180 79432 527232 79484
rect 121092 79160 121144 79212
rect 125324 79024 125376 79076
rect 125416 78956 125468 79008
rect 157340 79228 157392 79280
rect 157432 79228 157484 79280
rect 157892 79228 157944 79280
rect 157984 79228 158036 79280
rect 171232 79364 171284 79416
rect 166632 79296 166684 79348
rect 171048 79296 171100 79348
rect 173532 79364 173584 79416
rect 176292 79364 176344 79416
rect 580540 79364 580592 79416
rect 171876 79296 171928 79348
rect 173992 79296 174044 79348
rect 176200 79296 176252 79348
rect 580172 79296 580224 79348
rect 136180 79092 136232 79144
rect 161572 79160 161624 79212
rect 165804 79160 165856 79212
rect 172336 79228 172388 79280
rect 183100 79228 183152 79280
rect 167092 79160 167144 79212
rect 167276 79160 167328 79212
rect 168012 79160 168064 79212
rect 152648 79092 152700 79144
rect 154212 79092 154264 79144
rect 155132 79092 155184 79144
rect 167368 79092 167420 79144
rect 168380 79092 168432 79144
rect 168656 79092 168708 79144
rect 171048 79160 171100 79212
rect 174636 79160 174688 79212
rect 174728 79160 174780 79212
rect 183192 79160 183244 79212
rect 249800 79092 249852 79144
rect 135536 79024 135588 79076
rect 139952 79024 140004 79076
rect 145288 79024 145340 79076
rect 152372 79024 152424 79076
rect 153200 79024 153252 79076
rect 160100 79024 160152 79076
rect 161480 79024 161532 79076
rect 165804 79024 165856 79076
rect 167184 79024 167236 79076
rect 167552 79024 167604 79076
rect 168288 79024 168340 79076
rect 195980 79024 196032 79076
rect 151728 78956 151780 79008
rect 152648 78956 152700 79008
rect 153384 78956 153436 79008
rect 153844 78956 153896 79008
rect 154856 78956 154908 79008
rect 132776 78888 132828 78940
rect 148416 78888 148468 78940
rect 157432 78888 157484 78940
rect 157800 78888 157852 78940
rect 159180 78888 159232 78940
rect 160652 78956 160704 79008
rect 161020 78956 161072 79008
rect 162216 78956 162268 79008
rect 267832 78956 267884 79008
rect 167184 78888 167236 78940
rect 167276 78888 167328 78940
rect 213920 78888 213972 78940
rect 131028 78820 131080 78872
rect 137376 78820 137428 78872
rect 137836 78820 137888 78872
rect 150992 78820 151044 78872
rect 151728 78820 151780 78872
rect 157340 78820 157392 78872
rect 160836 78820 160888 78872
rect 161020 78820 161072 78872
rect 172152 78820 172204 78872
rect 172244 78820 172296 78872
rect 174728 78820 174780 78872
rect 176752 78820 176804 78872
rect 266360 78820 266412 78872
rect 129648 78752 129700 78804
rect 130108 78752 130160 78804
rect 132592 78752 132644 78804
rect 133052 78752 133104 78804
rect 140964 78752 141016 78804
rect 141424 78752 141476 78804
rect 148048 78752 148100 78804
rect 127164 78684 127216 78736
rect 127992 78684 128044 78736
rect 129004 78684 129056 78736
rect 129188 78684 129240 78736
rect 132776 78684 132828 78736
rect 133236 78684 133288 78736
rect 152280 78684 152332 78736
rect 152464 78684 152516 78736
rect 158628 78752 158680 78804
rect 159088 78752 159140 78804
rect 159640 78752 159692 78804
rect 160100 78752 160152 78804
rect 171508 78752 171560 78804
rect 171968 78752 172020 78804
rect 172428 78752 172480 78804
rect 172520 78752 172572 78804
rect 397460 78752 397512 78804
rect 125784 78616 125836 78668
rect 129924 78616 129976 78668
rect 132868 78616 132920 78668
rect 133052 78616 133104 78668
rect 144460 78616 144512 78668
rect 144828 78616 144880 78668
rect 147772 78616 147824 78668
rect 148140 78616 148192 78668
rect 150440 78616 150492 78668
rect 154304 78616 154356 78668
rect 426440 78684 426492 78736
rect 162584 78616 162636 78668
rect 162952 78616 163004 78668
rect 163320 78616 163372 78668
rect 166264 78616 166316 78668
rect 168012 78616 168064 78668
rect 168380 78616 168432 78668
rect 173808 78616 173860 78668
rect 122196 78548 122248 78600
rect 128636 78548 128688 78600
rect 141148 78548 141200 78600
rect 141976 78548 142028 78600
rect 146300 78548 146352 78600
rect 162216 78548 162268 78600
rect 166908 78548 166960 78600
rect 171968 78548 172020 78600
rect 172612 78548 172664 78600
rect 176752 78548 176804 78600
rect 125784 78480 125836 78532
rect 127072 78480 127124 78532
rect 146760 78480 146812 78532
rect 155868 78480 155920 78532
rect 156696 78480 156748 78532
rect 157432 78480 157484 78532
rect 161020 78480 161072 78532
rect 167184 78480 167236 78532
rect 170864 78480 170916 78532
rect 171876 78480 171928 78532
rect 255964 78480 256016 78532
rect 160100 78412 160152 78464
rect 160376 78412 160428 78464
rect 160744 78412 160796 78464
rect 162308 78412 162360 78464
rect 315304 78412 315356 78464
rect 126980 78344 127032 78396
rect 128360 78344 128412 78396
rect 150348 78344 150400 78396
rect 150716 78344 150768 78396
rect 162768 78344 162820 78396
rect 436744 78344 436796 78396
rect 120724 78276 120776 78328
rect 128268 78276 128320 78328
rect 148968 78276 149020 78328
rect 166264 78276 166316 78328
rect 116584 78208 116636 78260
rect 128820 78208 128872 78260
rect 142436 78208 142488 78260
rect 142712 78208 142764 78260
rect 145012 78208 145064 78260
rect 145748 78208 145800 78260
rect 155408 78208 155460 78260
rect 159640 78208 159692 78260
rect 161756 78208 161808 78260
rect 171876 78276 171928 78328
rect 172060 78276 172112 78328
rect 178776 78276 178828 78328
rect 167368 78208 167420 78260
rect 167552 78208 167604 78260
rect 169024 78208 169076 78260
rect 169208 78208 169260 78260
rect 113824 78140 113876 78192
rect 126796 78140 126848 78192
rect 139400 78140 139452 78192
rect 140136 78140 140188 78192
rect 142068 78140 142120 78192
rect 128268 78072 128320 78124
rect 150624 78072 150676 78124
rect 152372 78140 152424 78192
rect 158260 78140 158312 78192
rect 158720 78140 158772 78192
rect 162308 78140 162360 78192
rect 163136 78140 163188 78192
rect 483020 78208 483072 78260
rect 153384 78072 153436 78124
rect 154120 78072 154172 78124
rect 155500 78072 155552 78124
rect 155868 78072 155920 78124
rect 156144 78072 156196 78124
rect 156420 78072 156472 78124
rect 160100 78072 160152 78124
rect 161296 78072 161348 78124
rect 163228 78072 163280 78124
rect 171784 78072 171836 78124
rect 93124 78004 93176 78056
rect 127440 78004 127492 78056
rect 140504 78004 140556 78056
rect 146300 78004 146352 78056
rect 150992 78004 151044 78056
rect 151176 78004 151228 78056
rect 151636 78004 151688 78056
rect 154488 78004 154540 78056
rect 158628 78004 158680 78056
rect 159180 78004 159232 78056
rect 10324 77936 10376 77988
rect 125968 77936 126020 77988
rect 126796 77936 126848 77988
rect 128544 77936 128596 77988
rect 131764 77936 131816 77988
rect 132224 77936 132276 77988
rect 133236 77936 133288 77988
rect 133420 77936 133472 77988
rect 141608 77936 141660 77988
rect 141792 77936 141844 77988
rect 142252 77936 142304 77988
rect 152372 77936 152424 77988
rect 152648 77936 152700 77988
rect 154120 77868 154172 77920
rect 155500 77868 155552 77920
rect 157616 77868 157668 77920
rect 161572 77936 161624 77988
rect 162124 77936 162176 77988
rect 145012 77800 145064 77852
rect 145380 77800 145432 77852
rect 154672 77800 154724 77852
rect 158260 77800 158312 77852
rect 162216 77868 162268 77920
rect 164516 78004 164568 78056
rect 498200 78140 498252 78192
rect 171968 78072 172020 78124
rect 532700 78072 532752 78124
rect 165620 77936 165672 77988
rect 170588 77936 170640 77988
rect 170680 77936 170732 77988
rect 574744 78004 574796 78056
rect 143172 77732 143224 77784
rect 148416 77732 148468 77784
rect 151452 77732 151504 77784
rect 153844 77732 153896 77784
rect 159180 77732 159232 77784
rect 168288 77732 168340 77784
rect 123484 77664 123536 77716
rect 134800 77664 134852 77716
rect 155960 77664 156012 77716
rect 162124 77664 162176 77716
rect 162308 77664 162360 77716
rect 167184 77664 167236 77716
rect 168472 77664 168524 77716
rect 168748 77664 168800 77716
rect 171324 77868 171376 77920
rect 581092 77936 581144 77988
rect 172704 77868 172756 77920
rect 331220 77868 331272 77920
rect 171600 77800 171652 77852
rect 176292 77800 176344 77852
rect 172152 77732 172204 77784
rect 171600 77664 171652 77716
rect 176200 77664 176252 77716
rect 182916 77664 182968 77716
rect 144920 77596 144972 77648
rect 145840 77596 145892 77648
rect 160928 77596 160980 77648
rect 242164 77596 242216 77648
rect 139676 77528 139728 77580
rect 122104 77460 122156 77512
rect 127348 77460 127400 77512
rect 128820 77460 128872 77512
rect 129832 77460 129884 77512
rect 140780 77460 140832 77512
rect 159180 77460 159232 77512
rect 172060 77528 172112 77580
rect 165620 77460 165672 77512
rect 166172 77460 166224 77512
rect 166264 77460 166316 77512
rect 166448 77460 166500 77512
rect 167184 77460 167236 77512
rect 167736 77460 167788 77512
rect 169668 77460 169720 77512
rect 170220 77460 170272 77512
rect 170404 77460 170456 77512
rect 172336 77460 172388 77512
rect 132868 77392 132920 77444
rect 133696 77392 133748 77444
rect 141976 77392 142028 77444
rect 176384 77392 176436 77444
rect 152372 77324 152424 77376
rect 167276 77324 167328 77376
rect 168564 77324 168616 77376
rect 168840 77324 168892 77376
rect 168932 77324 168984 77376
rect 169116 77324 169168 77376
rect 125048 77256 125100 77308
rect 126704 77256 126756 77308
rect 144828 77256 144880 77308
rect 166632 77256 166684 77308
rect 171784 77256 171836 77308
rect 480260 77256 480312 77308
rect 124864 77188 124916 77240
rect 131212 77188 131264 77240
rect 137008 77188 137060 77240
rect 138940 77188 138992 77240
rect 149336 77188 149388 77240
rect 150072 77188 150124 77240
rect 152372 77188 152424 77240
rect 226340 77188 226392 77240
rect 130292 77120 130344 77172
rect 130568 77120 130620 77172
rect 146208 77120 146260 77172
rect 240140 77120 240192 77172
rect 139308 77052 139360 77104
rect 140504 77052 140556 77104
rect 147312 77052 147364 77104
rect 260840 77052 260892 77104
rect 122840 76984 122892 77036
rect 134892 76984 134944 77036
rect 147956 76984 148008 77036
rect 296720 76984 296772 77036
rect 156052 76916 156104 76968
rect 331128 76916 331180 76968
rect 118700 76848 118752 76900
rect 134984 76848 135036 76900
rect 143080 76848 143132 76900
rect 152372 76848 152424 76900
rect 157432 76848 157484 76900
rect 158352 76848 158404 76900
rect 102140 76780 102192 76832
rect 133512 76780 133564 76832
rect 70400 76712 70452 76764
rect 125416 76712 125468 76764
rect 155040 76712 155092 76764
rect 346400 76848 346452 76900
rect 167276 76780 167328 76832
rect 167920 76780 167972 76832
rect 168840 76780 168892 76832
rect 169392 76780 169444 76832
rect 173992 76780 174044 76832
rect 174360 76780 174412 76832
rect 174452 76780 174504 76832
rect 374000 76780 374052 76832
rect 171232 76712 171284 76764
rect 408500 76712 408552 76764
rect 93860 76644 93912 76696
rect 132500 76644 132552 76696
rect 142620 76644 142672 76696
rect 144552 76644 144604 76696
rect 159456 76644 159508 76696
rect 433340 76644 433392 76696
rect 69020 76576 69072 76628
rect 130752 76576 130804 76628
rect 165804 76576 165856 76628
rect 166080 76576 166132 76628
rect 169116 76576 169168 76628
rect 169484 76576 169536 76628
rect 171784 76576 171836 76628
rect 471980 76576 472032 76628
rect 6920 76508 6972 76560
rect 125140 76508 125192 76560
rect 169208 76508 169260 76560
rect 558920 76508 558972 76560
rect 155224 76440 155276 76492
rect 208400 76440 208452 76492
rect 149060 76372 149112 76424
rect 149520 76372 149572 76424
rect 151636 76372 151688 76424
rect 197360 76372 197412 76424
rect 127440 76304 127492 76356
rect 128084 76304 128136 76356
rect 149428 76304 149480 76356
rect 149980 76304 150032 76356
rect 155684 76304 155736 76356
rect 172520 76304 172572 76356
rect 162492 76236 162544 76288
rect 171784 76236 171836 76288
rect 165896 76168 165948 76220
rect 166172 76168 166224 76220
rect 125140 76032 125192 76084
rect 132408 76032 132460 76084
rect 136088 76032 136140 76084
rect 136456 76032 136508 76084
rect 165896 76032 165948 76084
rect 166540 76032 166592 76084
rect 128544 75964 128596 76016
rect 129096 75964 129148 76016
rect 133880 75964 133932 76016
rect 135536 75964 135588 76016
rect 151728 75896 151780 75948
rect 154856 75896 154908 75948
rect 139952 75828 140004 75880
rect 173256 75896 173308 75948
rect 172520 75828 172572 75880
rect 243728 75828 243780 75880
rect 156788 75760 156840 75812
rect 229192 75760 229244 75812
rect 130476 75692 130528 75744
rect 135260 75692 135312 75744
rect 150624 75692 150676 75744
rect 258080 75692 258132 75744
rect 128636 75624 128688 75676
rect 129556 75624 129608 75676
rect 151084 75624 151136 75676
rect 259460 75624 259512 75676
rect 154580 75556 154632 75608
rect 288532 75556 288584 75608
rect 121460 75488 121512 75540
rect 135076 75488 135128 75540
rect 151360 75488 151412 75540
rect 288440 75488 288492 75540
rect 51080 75420 51132 75472
rect 129372 75420 129424 75472
rect 129740 75420 129792 75472
rect 135720 75420 135772 75472
rect 156144 75420 156196 75472
rect 340144 75420 340196 75472
rect 107660 75352 107712 75404
rect 133788 75352 133840 75404
rect 134156 75352 134208 75404
rect 134616 75352 134668 75404
rect 155684 75352 155736 75404
rect 359372 75352 359424 75404
rect 49700 75284 49752 75336
rect 129464 75284 129516 75336
rect 131212 75284 131264 75336
rect 132316 75284 132368 75336
rect 135536 75284 135588 75336
rect 136272 75284 136324 75336
rect 143816 75284 143868 75336
rect 144276 75284 144328 75336
rect 149244 75284 149296 75336
rect 150164 75284 150216 75336
rect 157432 75284 157484 75336
rect 158168 75284 158220 75336
rect 163596 75284 163648 75336
rect 46940 75216 46992 75268
rect 124680 75216 124732 75268
rect 129924 75216 129976 75268
rect 130384 75216 130436 75268
rect 131488 75216 131540 75268
rect 131856 75216 131908 75268
rect 132684 75216 132736 75268
rect 133604 75216 133656 75268
rect 134616 75216 134668 75268
rect 135168 75216 135220 75268
rect 135996 75216 136048 75268
rect 136548 75216 136600 75268
rect 137100 75216 137152 75268
rect 137284 75216 137336 75268
rect 138112 75216 138164 75268
rect 138296 75216 138348 75268
rect 138848 75216 138900 75268
rect 139032 75216 139084 75268
rect 139952 75216 140004 75268
rect 140228 75216 140280 75268
rect 141056 75216 141108 75268
rect 141332 75216 141384 75268
rect 142620 75216 142672 75268
rect 142988 75216 143040 75268
rect 145104 75216 145156 75268
rect 145288 75216 145340 75268
rect 145472 75216 145524 75268
rect 145656 75216 145708 75268
rect 146392 75216 146444 75268
rect 146668 75216 146720 75268
rect 146760 75216 146812 75268
rect 146944 75216 146996 75268
rect 147956 75216 148008 75268
rect 148600 75216 148652 75268
rect 149336 75216 149388 75268
rect 149796 75216 149848 75268
rect 152004 75216 152056 75268
rect 152464 75216 152516 75268
rect 157524 75216 157576 75268
rect 157800 75216 157852 75268
rect 158904 75216 158956 75268
rect 159088 75216 159140 75268
rect 160008 75216 160060 75268
rect 160836 75216 160888 75268
rect 163228 75216 163280 75268
rect 163688 75216 163740 75268
rect 164424 75216 164476 75268
rect 164976 75216 165028 75268
rect 165436 75284 165488 75336
rect 481640 75284 481692 75336
rect 489920 75216 489972 75268
rect 26240 75148 26292 75200
rect 125968 75148 126020 75200
rect 126612 75148 126664 75200
rect 130016 75148 130068 75200
rect 130660 75148 130712 75200
rect 131304 75148 131356 75200
rect 131580 75148 131632 75200
rect 135720 75148 135772 75200
rect 136364 75148 136416 75200
rect 139676 75148 139728 75200
rect 140320 75148 140372 75200
rect 142252 75148 142304 75200
rect 142896 75148 142948 75200
rect 144000 75148 144052 75200
rect 144460 75148 144512 75200
rect 147772 75148 147824 75200
rect 148692 75148 148744 75200
rect 149428 75148 149480 75200
rect 149888 75148 149940 75200
rect 151912 75148 151964 75200
rect 152372 75148 152424 75200
rect 126060 75080 126112 75132
rect 126888 75080 126940 75132
rect 132960 75080 133012 75132
rect 133328 75080 133380 75132
rect 138296 75080 138348 75132
rect 138756 75080 138808 75132
rect 141056 75080 141108 75132
rect 141792 75080 141844 75132
rect 145104 75080 145156 75132
rect 145932 75080 145984 75132
rect 146576 75080 146628 75132
rect 146944 75080 146996 75132
rect 149152 75080 149204 75132
rect 156696 75080 156748 75132
rect 131580 75012 131632 75064
rect 132132 75012 132184 75064
rect 136916 75012 136968 75064
rect 137560 75012 137612 75064
rect 143540 75012 143592 75064
rect 144368 75012 144420 75064
rect 146668 75012 146720 75064
rect 147496 75012 147548 75064
rect 124404 74944 124456 74996
rect 127256 74944 127308 74996
rect 127624 74944 127676 74996
rect 128452 74944 128504 74996
rect 128912 74944 128964 74996
rect 137008 74944 137060 74996
rect 137744 74944 137796 74996
rect 146576 74944 146628 74996
rect 147220 74944 147272 74996
rect 151912 74876 151964 74928
rect 153108 74876 153160 74928
rect 157616 75148 157668 75200
rect 158076 75148 158128 75200
rect 162952 75148 163004 75200
rect 163780 75148 163832 75200
rect 164516 75148 164568 75200
rect 165160 75148 165212 75200
rect 157524 75080 157576 75132
rect 157984 75080 158036 75132
rect 163044 75080 163096 75132
rect 163872 75080 163924 75132
rect 163688 74944 163740 74996
rect 164884 74944 164936 74996
rect 506480 75148 506532 75200
rect 169760 75080 169812 75132
rect 170128 75080 170180 75132
rect 171508 75012 171560 75064
rect 172428 75012 172480 75064
rect 173532 74876 173584 74928
rect 151820 74808 151872 74860
rect 152648 74808 152700 74860
rect 127348 74672 127400 74724
rect 128176 74672 128228 74724
rect 139124 74468 139176 74520
rect 140136 74468 140188 74520
rect 143080 74468 143132 74520
rect 223580 74468 223632 74520
rect 243728 74468 243780 74520
rect 347504 74468 347556 74520
rect 145748 74400 145800 74452
rect 251180 74400 251232 74452
rect 156236 74332 156288 74384
rect 270040 74332 270092 74384
rect 151544 74264 151596 74316
rect 189080 74264 189132 74316
rect 208400 74264 208452 74316
rect 322940 74264 322992 74316
rect 156604 74196 156656 74248
rect 301136 74196 301188 74248
rect 128268 74128 128320 74180
rect 229100 74128 229152 74180
rect 229192 74128 229244 74180
rect 382924 74128 382976 74180
rect 4160 74060 4212 74112
rect 125600 74060 125652 74112
rect 154304 74060 154356 74112
rect 318800 74060 318852 74112
rect 118792 73992 118844 74044
rect 134708 73992 134760 74044
rect 157248 73992 157300 74044
rect 324320 73992 324372 74044
rect 60740 73924 60792 73976
rect 130200 73924 130252 73976
rect 156972 73924 157024 73976
rect 331864 73924 331916 73976
rect 30380 73856 30432 73908
rect 126336 73856 126388 73908
rect 126796 73856 126848 73908
rect 156420 73856 156472 73908
rect 362960 73856 363012 73908
rect 127992 73788 128044 73840
rect 158628 73788 158680 73840
rect 368480 73788 368532 73840
rect 141700 73720 141752 73772
rect 209780 73720 209832 73772
rect 193864 73652 193916 73704
rect 214104 73652 214156 73704
rect 369124 73652 369176 73704
rect 374736 73652 374788 73704
rect 137376 73380 137428 73432
rect 142988 73380 143040 73432
rect 339132 73244 339184 73296
rect 341064 73244 341116 73296
rect 126244 73176 126296 73228
rect 130844 73176 130896 73228
rect 151268 73108 151320 73160
rect 155316 73108 155368 73160
rect 170864 73108 170916 73160
rect 580172 73108 580224 73160
rect 150716 73040 150768 73092
rect 155776 73040 155828 73092
rect 258080 72836 258132 72888
rect 268200 72836 268252 72888
rect 166724 72768 166776 72820
rect 181444 72768 181496 72820
rect 259460 72768 259512 72820
rect 275376 72768 275428 72820
rect 150900 72700 150952 72752
rect 280068 72700 280120 72752
rect 149980 72632 150032 72684
rect 307760 72632 307812 72684
rect 150072 72564 150124 72616
rect 311900 72564 311952 72616
rect 114560 72496 114612 72548
rect 134432 72496 134484 72548
rect 153200 72496 153252 72548
rect 340880 72496 340932 72548
rect 96620 72428 96672 72480
rect 132592 72428 132644 72480
rect 158352 72428 158404 72480
rect 354680 72428 354732 72480
rect 288440 72156 288492 72208
rect 296168 72156 296220 72208
rect 378416 71748 378468 71800
rect 384764 71748 384816 71800
rect 150992 71680 151044 71732
rect 215300 71680 215352 71732
rect 229100 71680 229152 71732
rect 258724 71680 258776 71732
rect 349804 71680 349856 71732
rect 355508 71680 355560 71732
rect 359372 71680 359424 71732
rect 365076 71680 365128 71732
rect 3424 71612 3476 71664
rect 9036 71612 9088 71664
rect 189080 71612 189132 71664
rect 286324 71612 286376 71664
rect 154672 71544 154724 71596
rect 255320 71544 255372 71596
rect 150808 71476 150860 71528
rect 264244 71476 264296 71528
rect 154856 71408 154908 71460
rect 271880 71408 271932 71460
rect 155500 71340 155552 71392
rect 287612 71340 287664 71392
rect 301136 71340 301188 71392
rect 311164 71340 311216 71392
rect 324320 71340 324372 71392
rect 330484 71340 330536 71392
rect 155408 71272 155460 71324
rect 316684 71272 316736 71324
rect 322940 71272 322992 71324
rect 332600 71272 332652 71324
rect 154764 71204 154816 71256
rect 339408 71204 339460 71256
rect 362960 71204 363012 71256
rect 370504 71204 370556 71256
rect 165068 71136 165120 71188
rect 500960 71136 501012 71188
rect 165528 71068 165580 71120
rect 507860 71068 507912 71120
rect 138020 71000 138072 71052
rect 165068 71000 165120 71052
rect 168012 71000 168064 71052
rect 539600 71000 539652 71052
rect 148416 70932 148468 70984
rect 190460 70932 190512 70984
rect 214104 70932 214156 70984
rect 257344 70932 257396 70984
rect 164056 70524 164108 70576
rect 170404 70524 170456 70576
rect 155316 70320 155368 70372
rect 250444 70320 250496 70372
rect 155776 70252 155828 70304
rect 271788 70252 271840 70304
rect 140044 70184 140096 70236
rect 173440 70184 173492 70236
rect 173532 70184 173584 70236
rect 327724 70184 327776 70236
rect 155960 70116 156012 70168
rect 326988 70116 327040 70168
rect 154672 70048 154724 70100
rect 327816 70048 327868 70100
rect 155868 69980 155920 70032
rect 338764 69980 338816 70032
rect 156880 69912 156932 69964
rect 361580 69912 361632 69964
rect 164792 69844 164844 69896
rect 505100 69844 505152 69896
rect 166356 69776 166408 69828
rect 523040 69776 523092 69828
rect 137284 69708 137336 69760
rect 149152 69708 149204 69760
rect 167092 69708 167144 69760
rect 536840 69708 536892 69760
rect 138572 69640 138624 69692
rect 140228 69640 140280 69692
rect 169116 69640 169168 69692
rect 564440 69640 564492 69692
rect 141516 69572 141568 69624
rect 209872 69572 209924 69624
rect 215300 68960 215352 69012
rect 218152 68960 218204 69012
rect 255320 68960 255372 69012
rect 258816 68960 258868 69012
rect 288532 68960 288584 69012
rect 295340 68960 295392 69012
rect 331128 68960 331180 69012
rect 336004 68960 336056 69012
rect 346400 68960 346452 69012
rect 349804 68960 349856 69012
rect 341064 68620 341116 68672
rect 352564 68620 352616 68672
rect 355508 68620 355560 68672
rect 359280 68620 359332 68672
rect 332600 68552 332652 68604
rect 347228 68552 347280 68604
rect 153752 68484 153804 68536
rect 358820 68484 358872 68536
rect 166264 68416 166316 68468
rect 525800 68416 525852 68468
rect 169024 68348 169076 68400
rect 557540 68348 557592 68400
rect 170772 68280 170824 68332
rect 564532 68280 564584 68332
rect 365076 68212 365128 68264
rect 369124 68212 369176 68264
rect 271880 68144 271932 68196
rect 275284 68144 275336 68196
rect 137192 67532 137244 67584
rect 138664 67532 138716 67584
rect 270040 67532 270092 67584
rect 275192 67532 275244 67584
rect 306932 67532 306984 67584
rect 309784 67532 309836 67584
rect 384764 67532 384816 67584
rect 387064 67532 387116 67584
rect 326988 67464 327040 67516
rect 329104 67464 329156 67516
rect 138480 67056 138532 67108
rect 167092 67056 167144 67108
rect 139952 66988 140004 67040
rect 189080 66988 189132 67040
rect 142804 66920 142856 66972
rect 220820 66920 220872 66972
rect 145564 66852 145616 66904
rect 256700 66852 256752 66904
rect 339408 66716 339460 66768
rect 345664 66716 345716 66768
rect 271788 66444 271840 66496
rect 278780 66444 278832 66496
rect 268200 66172 268252 66224
rect 271144 66172 271196 66224
rect 287612 66172 287664 66224
rect 291108 66172 291160 66224
rect 347504 66172 347556 66224
rect 349988 66172 350040 66224
rect 142712 65764 142764 65816
rect 218060 65764 218112 65816
rect 218152 65764 218204 65816
rect 226248 65764 226300 65816
rect 144184 65696 144236 65748
rect 238760 65696 238812 65748
rect 280068 65696 280120 65748
rect 292856 65696 292908 65748
rect 295340 65696 295392 65748
rect 303620 65696 303672 65748
rect 311164 65696 311216 65748
rect 316040 65696 316092 65748
rect 330484 65696 330536 65748
rect 340788 65696 340840 65748
rect 359280 65696 359332 65748
rect 370964 65696 371016 65748
rect 163412 65628 163464 65680
rect 484400 65628 484452 65680
rect 167736 65560 167788 65612
rect 543740 65560 543792 65612
rect 170220 65492 170272 65544
rect 572720 65492 572772 65544
rect 361580 64880 361632 64932
rect 364984 64880 365036 64932
rect 264244 64404 264296 64456
rect 269764 64404 269816 64456
rect 152556 64268 152608 64320
rect 338120 64268 338172 64320
rect 157984 64200 158036 64252
rect 374092 64200 374144 64252
rect 170128 64132 170180 64184
rect 568580 64132 568632 64184
rect 352564 63996 352616 64048
rect 357348 63996 357400 64048
rect 275376 63724 275428 63776
rect 278412 63724 278464 63776
rect 278780 63588 278832 63640
rect 283012 63588 283064 63640
rect 139860 63112 139912 63164
rect 184940 63112 184992 63164
rect 142620 63044 142672 63096
rect 224960 63044 225012 63096
rect 147128 62976 147180 63028
rect 274640 62976 274692 63028
rect 152464 62908 152516 62960
rect 340972 62908 341024 62960
rect 163320 62840 163372 62892
rect 481732 62840 481784 62892
rect 170680 62772 170732 62824
rect 514760 62772 514812 62824
rect 316040 62568 316092 62620
rect 318984 62568 319036 62620
rect 138388 62024 138440 62076
rect 142804 62024 142856 62076
rect 349988 61956 350040 62008
rect 353944 61956 353996 62008
rect 370964 61752 371016 61804
rect 376668 61752 376720 61804
rect 257344 61616 257396 61668
rect 262864 61616 262916 61668
rect 275192 61616 275244 61668
rect 297364 61616 297416 61668
rect 148324 61548 148376 61600
rect 292580 61548 292632 61600
rect 340788 61548 340840 61600
rect 354036 61548 354088 61600
rect 149704 61480 149756 61532
rect 306380 61480 306432 61532
rect 347228 61480 347280 61532
rect 363604 61480 363656 61532
rect 153660 61412 153712 61464
rect 362960 61412 363012 61464
rect 102232 61344 102284 61396
rect 125324 61344 125376 61396
rect 157892 61344 157944 61396
rect 412640 61344 412692 61396
rect 292856 60936 292908 60988
rect 295984 60936 296036 60988
rect 338764 60732 338816 60784
rect 344284 60732 344336 60784
rect 183284 60664 183336 60716
rect 580172 60664 580224 60716
rect 327816 60596 327868 60648
rect 332600 60596 332652 60648
rect 318984 60392 319036 60444
rect 327908 60392 327960 60444
rect 141424 60120 141476 60172
rect 207020 60120 207072 60172
rect 226248 60120 226300 60172
rect 247684 60120 247736 60172
rect 144092 60052 144144 60104
rect 233240 60052 233292 60104
rect 149612 59984 149664 60036
rect 305000 59984 305052 60036
rect 258816 59916 258868 59968
rect 264336 59916 264388 59968
rect 120080 59576 120132 59628
rect 123484 59576 123536 59628
rect 3056 59304 3108 59356
rect 181260 59304 181312 59356
rect 258724 59304 258776 59356
rect 261484 59304 261536 59356
rect 303620 59304 303672 59356
rect 307024 59304 307076 59356
rect 357348 59304 357400 59356
rect 363696 59304 363748 59356
rect 286324 58760 286376 58812
rect 298744 58760 298796 58812
rect 283012 58692 283064 58744
rect 291844 58692 291896 58744
rect 296168 58692 296220 58744
rect 313924 58692 313976 58744
rect 275284 58624 275336 58676
rect 283656 58624 283708 58676
rect 291108 58624 291160 58676
rect 311164 58624 311216 58676
rect 336004 58624 336056 58676
rect 362224 58624 362276 58676
rect 95240 57196 95292 57248
rect 125232 57196 125284 57248
rect 296076 57196 296128 57248
rect 301596 57196 301648 57248
rect 309784 57196 309836 57248
rect 323584 57196 323636 57248
rect 376668 57196 376720 57248
rect 384396 57196 384448 57248
rect 332600 56584 332652 56636
rect 336004 56584 336056 56636
rect 261484 56516 261536 56568
rect 264244 56516 264296 56568
rect 278412 56516 278464 56568
rect 280804 56516 280856 56568
rect 329104 56516 329156 56568
rect 333980 56516 334032 56568
rect 369124 56516 369176 56568
rect 371884 56516 371936 56568
rect 88340 55836 88392 55888
rect 125140 55836 125192 55888
rect 370504 55836 370556 55888
rect 387708 55836 387760 55888
rect 291844 54612 291896 54664
rect 295340 54612 295392 54664
rect 283656 54476 283708 54528
rect 292672 54476 292724 54528
rect 297364 54476 297416 54528
rect 326344 54476 326396 54528
rect 340144 54476 340196 54528
rect 343640 54476 343692 54528
rect 364984 54476 365036 54528
rect 374644 54476 374696 54528
rect 262864 54408 262916 54460
rect 269856 54408 269908 54460
rect 250444 54340 250496 54392
rect 253020 54340 253072 54392
rect 374736 54340 374788 54392
rect 380164 54340 380216 54392
rect 363604 53728 363656 53780
rect 366548 53728 366600 53780
rect 313924 53456 313976 53508
rect 316776 53456 316828 53508
rect 363696 53252 363748 53304
rect 367008 53252 367060 53304
rect 354036 53116 354088 53168
rect 356244 53116 356296 53168
rect 264336 53048 264388 53100
rect 281356 53048 281408 53100
rect 311164 53048 311216 53100
rect 318156 53048 318208 53100
rect 333980 53048 334032 53100
rect 340144 53048 340196 53100
rect 327908 52368 327960 52420
rect 332600 52368 332652 52420
rect 362224 52368 362276 52420
rect 365628 52368 365680 52420
rect 13820 51688 13872 51740
rect 125048 51688 125100 51740
rect 295340 51688 295392 51740
rect 318064 51688 318116 51740
rect 387708 51212 387760 51264
rect 391204 51212 391256 51264
rect 253020 51008 253072 51060
rect 258724 51008 258776 51060
rect 353944 51008 353996 51060
rect 356704 51008 356756 51060
rect 269764 50940 269816 50992
rect 273168 50940 273220 50992
rect 247684 50328 247736 50380
rect 274732 50328 274784 50380
rect 331864 50328 331916 50380
rect 339960 50328 340012 50380
rect 343640 50328 343692 50380
rect 359464 50328 359516 50380
rect 366548 49784 366600 49836
rect 373264 49784 373316 49836
rect 271144 49648 271196 49700
rect 277492 49648 277544 49700
rect 307024 49648 307076 49700
rect 311992 49648 312044 49700
rect 332600 49648 332652 49700
rect 337384 49648 337436 49700
rect 349804 48220 349856 48272
rect 352012 48220 352064 48272
rect 365628 48220 365680 48272
rect 370504 48220 370556 48272
rect 367008 48152 367060 48204
rect 371240 48152 371292 48204
rect 356244 47608 356296 47660
rect 374184 47608 374236 47660
rect 163228 47540 163280 47592
rect 488540 47540 488592 47592
rect 344284 47268 344336 47320
rect 346400 47268 346452 47320
rect 118516 46860 118568 46912
rect 580172 46860 580224 46912
rect 264244 46792 264296 46844
rect 267004 46792 267056 46844
rect 301596 46792 301648 46844
rect 304264 46792 304316 46844
rect 274732 46520 274784 46572
rect 279424 46520 279476 46572
rect 273168 46248 273220 46300
rect 282184 46248 282236 46300
rect 277492 46180 277544 46232
rect 288440 46180 288492 46232
rect 292672 46180 292724 46232
rect 301504 46180 301556 46232
rect 339960 46180 340012 46232
rect 349804 46180 349856 46232
rect 311992 46044 312044 46096
rect 317420 46044 317472 46096
rect 281356 45568 281408 45620
rect 287704 45568 287756 45620
rect 3424 45500 3476 45552
rect 174084 45500 174136 45552
rect 327724 45092 327776 45144
rect 332600 45092 332652 45144
rect 346400 44888 346452 44940
rect 359556 44888 359608 44940
rect 67640 44820 67692 44872
rect 130200 44820 130252 44872
rect 139768 44820 139820 44872
rect 185032 44820 185084 44872
rect 340144 44820 340196 44872
rect 352104 44820 352156 44872
rect 318156 44684 318208 44736
rect 324320 44684 324372 44736
rect 374184 44616 374236 44668
rect 383016 44616 383068 44668
rect 336004 44140 336056 44192
rect 339408 44140 339460 44192
rect 317420 43392 317472 43444
rect 344284 43392 344336 43444
rect 371240 43120 371292 43172
rect 376024 43120 376076 43172
rect 269856 42916 269908 42968
rect 276020 42916 276072 42968
rect 316776 42780 316828 42832
rect 319444 42780 319496 42832
rect 352012 42712 352064 42764
rect 355324 42712 355376 42764
rect 280804 42236 280856 42288
rect 284300 42236 284352 42288
rect 316684 41828 316736 41880
rect 319812 41828 319864 41880
rect 324320 40672 324372 40724
rect 330484 40672 330536 40724
rect 339408 40672 339460 40724
rect 341064 40672 341116 40724
rect 352104 40672 352156 40724
rect 375288 40672 375340 40724
rect 288440 39992 288492 40044
rect 291844 39992 291896 40044
rect 323584 39992 323636 40044
rect 326436 39992 326488 40044
rect 276020 39380 276072 39432
rect 284944 39380 284996 39432
rect 332600 39380 332652 39432
rect 340144 39380 340196 39432
rect 258724 39312 258776 39364
rect 278044 39312 278096 39364
rect 326344 39312 326396 39364
rect 337936 39312 337988 39364
rect 345664 39312 345716 39364
rect 362224 39312 362276 39364
rect 45560 37884 45612 37936
rect 116584 37884 116636 37936
rect 282184 37884 282236 37936
rect 298284 37884 298336 37936
rect 375288 37884 375340 37936
rect 388444 37884 388496 37936
rect 284300 37476 284352 37528
rect 287428 37476 287480 37528
rect 380164 37272 380216 37324
rect 384304 37272 384356 37324
rect 319812 37204 319864 37256
rect 322848 37204 322900 37256
rect 337936 37204 337988 37256
rect 342904 37204 342956 37256
rect 355324 37204 355376 37256
rect 360844 37204 360896 37256
rect 341064 37136 341116 37188
rect 344376 37136 344428 37188
rect 340144 36592 340196 36644
rect 362132 36592 362184 36644
rect 7564 36524 7616 36576
rect 124220 36524 124272 36576
rect 172152 36524 172204 36576
rect 418160 36524 418212 36576
rect 382924 35912 382976 35964
rect 385684 35912 385736 35964
rect 148140 35300 148192 35352
rect 287060 35300 287112 35352
rect 287428 35300 287480 35352
rect 299204 35300 299256 35352
rect 356704 35300 356756 35352
rect 361580 35300 361632 35352
rect 148232 35232 148284 35284
rect 291200 35232 291252 35284
rect 38660 35164 38712 35216
rect 122196 35164 122248 35216
rect 153568 35164 153620 35216
rect 357440 35164 357492 35216
rect 278044 34552 278096 34604
rect 285680 34552 285732 34604
rect 141332 33940 141384 33992
rect 198740 33940 198792 33992
rect 344284 33940 344336 33992
rect 347596 33940 347648 33992
rect 141240 33872 141292 33924
rect 205640 33872 205692 33924
rect 142528 33804 142580 33856
rect 219440 33804 219492 33856
rect 376024 33804 376076 33856
rect 384488 33804 384540 33856
rect 145472 33736 145524 33788
rect 259460 33736 259512 33788
rect 322848 33736 322900 33788
rect 329104 33736 329156 33788
rect 383016 33736 383068 33788
rect 396724 33736 396776 33788
rect 171968 33056 172020 33108
rect 580172 33056 580224 33108
rect 361580 32988 361632 33040
rect 364984 32988 365036 33040
rect 384396 32784 384448 32836
rect 391940 32784 391992 32836
rect 139676 32716 139728 32768
rect 187700 32716 187752 32768
rect 370504 32716 370556 32768
rect 378140 32716 378192 32768
rect 141148 32648 141200 32700
rect 201500 32648 201552 32700
rect 267004 32648 267056 32700
rect 275284 32648 275336 32700
rect 285680 32648 285732 32700
rect 293960 32648 294012 32700
rect 362132 32648 362184 32700
rect 374736 32648 374788 32700
rect 160836 32580 160888 32632
rect 447140 32580 447192 32632
rect 3424 32512 3476 32564
rect 7656 32512 7708 32564
rect 166172 32512 166224 32564
rect 474004 32512 474056 32564
rect 163136 32444 163188 32496
rect 485780 32444 485832 32496
rect 31760 32376 31812 32428
rect 120724 32376 120776 32428
rect 164700 32376 164752 32428
rect 503720 32376 503772 32428
rect 374644 31764 374696 31816
rect 377404 31764 377456 31816
rect 349804 31696 349856 31748
rect 353392 31696 353444 31748
rect 318064 31492 318116 31544
rect 322940 31492 322992 31544
rect 326436 31220 326488 31272
rect 331220 31220 331272 31272
rect 291844 31152 291896 31204
rect 301596 31152 301648 31204
rect 337384 31152 337436 31204
rect 347044 31152 347096 31204
rect 299204 31084 299256 31136
rect 313280 31084 313332 31136
rect 342904 31084 342956 31136
rect 353484 31084 353536 31136
rect 371884 31084 371936 31136
rect 378784 31084 378836 31136
rect 164608 31016 164660 31068
rect 499580 31016 499632 31068
rect 279424 30268 279476 30320
rect 286324 30268 286376 30320
rect 387064 30268 387116 30320
rect 392584 30268 392636 30320
rect 298284 29996 298336 30048
rect 311164 29996 311216 30048
rect 293960 29928 294012 29980
rect 320824 29928 320876 29980
rect 148048 29860 148100 29912
rect 285680 29860 285732 29912
rect 298744 29860 298796 29912
rect 326436 29860 326488 29912
rect 154120 29792 154172 29844
rect 332600 29792 332652 29844
rect 152372 29724 152424 29776
rect 339500 29724 339552 29776
rect 152280 29656 152332 29708
rect 346400 29656 346452 29708
rect 391940 29656 391992 29708
rect 397552 29656 397604 29708
rect 157800 29588 157852 29640
rect 409880 29588 409932 29640
rect 287704 28908 287756 28960
rect 291108 28908 291160 28960
rect 378140 28908 378192 28960
rect 381544 28908 381596 28960
rect 360844 28772 360896 28824
rect 365168 28772 365220 28824
rect 144000 28568 144052 28620
rect 242900 28568 242952 28620
rect 145288 28500 145340 28552
rect 251272 28500 251324 28552
rect 145196 28432 145248 28484
rect 253940 28432 253992 28484
rect 344376 28432 344428 28484
rect 348884 28432 348936 28484
rect 145380 28364 145432 28416
rect 258080 28364 258132 28416
rect 304264 28364 304316 28416
rect 323492 28364 323544 28416
rect 347596 28364 347648 28416
rect 356704 28364 356756 28416
rect 171784 28296 171836 28348
rect 397460 28296 397512 28348
rect 167644 28228 167696 28280
rect 539692 28228 539744 28280
rect 353392 27684 353444 27736
rect 356060 27684 356112 27736
rect 378784 27684 378836 27736
rect 385040 27684 385092 27736
rect 330484 27548 330536 27600
rect 334256 27548 334308 27600
rect 359556 27548 359608 27600
rect 363328 27548 363380 27600
rect 397552 27548 397604 27600
rect 400864 27548 400916 27600
rect 140964 27344 141016 27396
rect 204260 27344 204312 27396
rect 141056 27276 141108 27328
rect 208400 27276 208452 27328
rect 142436 27208 142488 27260
rect 215300 27208 215352 27260
rect 142344 27140 142396 27192
rect 218152 27140 218204 27192
rect 143908 27072 143960 27124
rect 236000 27072 236052 27124
rect 295984 27072 296036 27124
rect 302884 27072 302936 27124
rect 149520 27004 149572 27056
rect 303620 27004 303672 27056
rect 313280 27004 313332 27056
rect 321744 27004 321796 27056
rect 171692 26936 171744 26988
rect 411260 26936 411312 26988
rect 168932 26868 168984 26920
rect 560300 26868 560352 26920
rect 331220 26460 331272 26512
rect 335360 26460 335412 26512
rect 353484 26256 353536 26308
rect 356152 26256 356204 26308
rect 140412 25984 140464 26036
rect 176752 25984 176804 26036
rect 139492 25916 139544 25968
rect 179420 25916 179472 25968
rect 139584 25848 139636 25900
rect 183560 25848 183612 25900
rect 139400 25780 139452 25832
rect 186320 25780 186372 25832
rect 140872 25712 140924 25764
rect 201592 25712 201644 25764
rect 291108 25712 291160 25764
rect 302240 25712 302292 25764
rect 147956 25644 148008 25696
rect 292672 25644 292724 25696
rect 374736 25644 374788 25696
rect 381636 25644 381688 25696
rect 157708 25576 157760 25628
rect 414020 25576 414072 25628
rect 167552 25508 167604 25560
rect 535460 25508 535512 25560
rect 348884 25236 348936 25288
rect 351828 25236 351880 25288
rect 301504 24828 301556 24880
rect 305644 24828 305696 24880
rect 377404 24828 377456 24880
rect 380164 24828 380216 24880
rect 286324 24692 286376 24744
rect 292764 24692 292816 24744
rect 363328 24692 363380 24744
rect 369124 24692 369176 24744
rect 147864 24624 147916 24676
rect 289820 24624 289872 24676
rect 334256 24624 334308 24676
rect 342260 24624 342312 24676
rect 356060 24624 356112 24676
rect 369860 24624 369912 24676
rect 384488 24624 384540 24676
rect 407212 24624 407264 24676
rect 157616 24556 157668 24608
rect 416780 24556 416832 24608
rect 168748 24488 168800 24540
rect 552020 24488 552072 24540
rect 169668 24420 169720 24472
rect 556160 24420 556212 24472
rect 168840 24352 168892 24404
rect 563060 24352 563112 24404
rect 3332 24284 3384 24336
rect 179880 24284 179932 24336
rect 183008 24284 183060 24336
rect 579620 24284 579672 24336
rect 169944 24216 169996 24268
rect 569960 24216 570012 24268
rect 169852 24148 169904 24200
rect 571340 24148 571392 24200
rect 170036 24080 170088 24132
rect 572812 24080 572864 24132
rect 320824 24012 320876 24064
rect 327724 24012 327776 24064
rect 135996 23400 136048 23452
rect 142344 23400 142396 23452
rect 319444 23400 319496 23452
rect 326344 23400 326396 23452
rect 391204 23400 391256 23452
rect 393320 23400 393372 23452
rect 302240 23264 302292 23316
rect 313280 23264 313332 23316
rect 3424 23196 3476 23248
rect 173992 23196 174044 23248
rect 284944 23196 284996 23248
rect 299296 23196 299348 23248
rect 311164 23196 311216 23248
rect 323584 23196 323636 23248
rect 356152 23196 356204 23248
rect 369952 23196 370004 23248
rect 172244 23128 172296 23180
rect 404360 23128 404412 23180
rect 163044 23060 163096 23112
rect 492680 23060 492732 23112
rect 167368 22992 167420 23044
rect 534080 22992 534132 23044
rect 63500 22924 63552 22976
rect 126336 22924 126388 22976
rect 167460 22924 167512 22976
rect 538220 22924 538272 22976
rect 35900 22856 35952 22908
rect 126980 22856 127032 22908
rect 167184 22856 167236 22908
rect 540980 22856 541032 22908
rect 22100 22788 22152 22840
rect 127532 22788 127584 22840
rect 167276 22788 167328 22840
rect 545120 22788 545172 22840
rect 118332 22720 118384 22772
rect 580264 22720 580316 22772
rect 321744 22108 321796 22160
rect 324320 22108 324372 22160
rect 301596 21768 301648 21820
rect 304264 21768 304316 21820
rect 329104 21768 329156 21820
rect 344284 21768 344336 21820
rect 152188 21700 152240 21752
rect 343640 21700 343692 21752
rect 160744 21632 160796 21684
rect 454040 21632 454092 21684
rect 165988 21564 166040 21616
rect 516140 21564 516192 21616
rect 165804 21496 165856 21548
rect 520280 21496 520332 21548
rect 165896 21428 165948 21480
rect 523132 21428 523184 21480
rect 85580 21360 85632 21412
rect 131764 21360 131816 21412
rect 166080 21360 166132 21412
rect 527180 21360 527232 21412
rect 362224 20612 362276 20664
rect 365076 20612 365128 20664
rect 396724 20612 396776 20664
rect 398932 20612 398984 20664
rect 299296 20340 299348 20392
rect 326528 20340 326580 20392
rect 145104 20272 145156 20324
rect 262220 20272 262272 20324
rect 313280 20272 313332 20324
rect 322204 20272 322256 20324
rect 323492 20272 323544 20324
rect 358084 20272 358136 20324
rect 369860 20272 369912 20324
rect 379520 20272 379572 20324
rect 145012 20204 145064 20256
rect 255320 20204 255372 20256
rect 255964 20204 256016 20256
rect 456800 20204 456852 20256
rect 143816 20136 143868 20188
rect 241520 20136 241572 20188
rect 242164 20136 242216 20188
rect 449900 20136 449952 20188
rect 157524 20068 157576 20120
rect 415400 20068 415452 20120
rect 164424 20000 164476 20052
rect 506572 20000 506624 20052
rect 164516 19932 164568 19984
rect 509240 19932 509292 19984
rect 356704 19252 356756 19304
rect 359556 19252 359608 19304
rect 369124 18980 369176 19032
rect 378692 18980 378744 19032
rect 359464 18912 359516 18964
rect 377404 18912 377456 18964
rect 143724 18844 143776 18896
rect 234620 18844 234672 18896
rect 275284 18844 275336 18896
rect 288440 18844 288492 18896
rect 292764 18844 292816 18896
rect 302056 18844 302108 18896
rect 347044 18844 347096 18896
rect 388536 18844 388588 18896
rect 164240 18776 164292 18828
rect 498292 18776 498344 18828
rect 164332 18708 164384 18760
rect 502340 18708 502392 18760
rect 168472 18640 168524 18692
rect 553400 18640 553452 18692
rect 81440 18572 81492 18624
rect 131672 18572 131724 18624
rect 168564 18572 168616 18624
rect 556252 18572 556304 18624
rect 351828 18028 351880 18080
rect 354772 18028 354824 18080
rect 400864 17960 400916 18012
rect 402980 17960 403032 18012
rect 365168 17892 365220 17944
rect 373448 17892 373500 17944
rect 379520 17892 379572 17944
rect 382280 17892 382332 17944
rect 369952 17348 370004 17400
rect 375380 17348 375432 17400
rect 342260 17212 342312 17264
rect 348700 17212 348752 17264
rect 392584 17212 392636 17264
rect 397184 17212 397236 17264
rect 324320 17008 324372 17060
rect 327080 17008 327132 17060
rect 143632 16124 143684 16176
rect 237656 16124 237708 16176
rect 288440 16124 288492 16176
rect 298744 16124 298796 16176
rect 302884 16124 302936 16176
rect 313924 16124 313976 16176
rect 326528 16124 326580 16176
rect 337016 16124 337068 16176
rect 152096 16056 152148 16108
rect 342904 16056 342956 16108
rect 344284 16056 344336 16108
rect 357348 16056 357400 16108
rect 358084 16056 358136 16108
rect 385868 16056 385920 16108
rect 153476 15988 153528 16040
rect 361120 15988 361172 16040
rect 385684 15988 385736 16040
rect 390560 15988 390612 16040
rect 157432 15920 157484 15972
rect 415492 15920 415544 15972
rect 157340 15852 157392 15904
rect 420184 15852 420236 15904
rect 302056 15240 302108 15292
rect 304264 15240 304316 15292
rect 380164 15172 380216 15224
rect 382924 15172 382976 15224
rect 305644 14832 305696 14884
rect 309600 14832 309652 14884
rect 149428 14764 149480 14816
rect 311440 14764 311492 14816
rect 159640 14696 159692 14748
rect 382372 14764 382424 14816
rect 382280 14696 382332 14748
rect 402520 14696 402572 14748
rect 159272 14628 159324 14680
rect 429200 14628 429252 14680
rect 159364 14560 159416 14612
rect 436744 14560 436796 14612
rect 159180 14492 159232 14544
rect 439136 14492 439188 14544
rect 162952 14424 163004 14476
rect 492312 14424 492364 14476
rect 377404 13812 377456 13864
rect 380900 13812 380952 13864
rect 304264 13744 304316 13796
rect 307024 13744 307076 13796
rect 385868 13744 385920 13796
rect 392584 13744 392636 13796
rect 153292 13132 153344 13184
rect 357532 13132 357584 13184
rect 153384 13064 153436 13116
rect 365812 13064 365864 13116
rect 375380 13064 375432 13116
rect 381728 13064 381780 13116
rect 323584 12384 323636 12436
rect 326252 12384 326304 12436
rect 348700 12384 348752 12436
rect 357072 12384 357124 12436
rect 381636 12384 381688 12436
rect 384396 12384 384448 12436
rect 390560 12384 390612 12436
rect 395344 12384 395396 12436
rect 397184 12384 397236 12436
rect 403716 12384 403768 12436
rect 304356 12316 304408 12368
rect 312544 12316 312596 12368
rect 326436 12316 326488 12368
rect 332692 12316 332744 12368
rect 152004 12248 152056 12300
rect 345296 12248 345348 12300
rect 357348 12248 357400 12300
rect 373356 12248 373408 12300
rect 373448 12248 373500 12300
rect 379520 12248 379572 12300
rect 151912 12180 151964 12232
rect 349252 12180 349304 12232
rect 354772 12180 354824 12232
rect 376024 12180 376076 12232
rect 162216 12112 162268 12164
rect 390652 12112 390704 12164
rect 159088 12044 159140 12096
rect 428464 12044 428516 12096
rect 158904 11976 158956 12028
rect 432052 11976 432104 12028
rect 158812 11908 158864 11960
rect 435088 11908 435140 11960
rect 160008 11840 160060 11892
rect 440332 11840 440384 11892
rect 162032 11772 162084 11824
rect 468208 11772 468260 11824
rect 169760 11704 169812 11756
rect 574652 11704 574704 11756
rect 364984 11636 365036 11688
rect 367744 11636 367796 11688
rect 378692 11636 378744 11688
rect 381268 11636 381320 11688
rect 117320 10548 117372 10600
rect 134248 10548 134300 10600
rect 106464 10480 106516 10532
rect 133052 10480 133104 10532
rect 78128 10412 78180 10464
rect 129096 10412 129148 10464
rect 149336 10412 149388 10464
rect 309784 10412 309836 10464
rect 25320 10344 25372 10396
rect 93124 10344 93176 10396
rect 99840 10344 99892 10396
rect 132960 10344 133012 10396
rect 149244 10344 149296 10396
rect 313832 10344 313884 10396
rect 35992 10276 36044 10328
rect 127440 10276 127492 10328
rect 167000 10276 167052 10328
rect 542728 10276 542780 10328
rect 147772 9596 147824 9648
rect 296076 9596 296128 9648
rect 309600 9596 309652 9648
rect 313096 9596 313148 9648
rect 315304 9596 315356 9648
rect 465172 9596 465224 9648
rect 160192 9528 160244 9580
rect 445024 9528 445076 9580
rect 165712 9460 165764 9512
rect 449900 9460 449952 9512
rect 160284 9392 160336 9444
rect 446220 9392 446272 9444
rect 160468 9324 160520 9376
rect 448612 9324 448664 9376
rect 60832 9256 60884 9308
rect 128360 9256 128412 9308
rect 161204 9256 161256 9308
rect 449808 9256 449860 9308
rect 59636 9188 59688 9240
rect 130108 9188 130160 9240
rect 160560 9188 160612 9240
rect 452108 9188 452160 9240
rect 53748 9120 53800 9172
rect 128728 9120 128780 9172
rect 160376 9120 160428 9172
rect 453304 9120 453356 9172
rect 52552 9052 52604 9104
rect 128636 9052 128688 9104
rect 160652 9052 160704 9104
rect 455696 9052 455748 9104
rect 45468 8984 45520 9036
rect 128544 8984 128596 9036
rect 161848 8984 161900 9036
rect 463976 8984 464028 9036
rect 9956 8916 10008 8968
rect 126152 8916 126204 8968
rect 161940 8916 161992 8968
rect 467472 8916 467524 8968
rect 327724 8848 327776 8900
rect 330392 8848 330444 8900
rect 357072 8848 357124 8900
rect 362316 8848 362368 8900
rect 322204 8304 322256 8356
rect 327080 8304 327132 8356
rect 116400 8032 116452 8084
rect 134156 8032 134208 8084
rect 105728 7964 105780 8016
rect 132868 7964 132920 8016
rect 98644 7896 98696 7948
rect 132776 7896 132828 7948
rect 142252 7896 142304 7948
rect 222752 7896 222804 7948
rect 84476 7828 84528 7880
rect 131580 7828 131632 7880
rect 143540 7828 143592 7880
rect 242992 7828 243044 7880
rect 48964 7760 49016 7812
rect 129188 7760 129240 7812
rect 144920 7760 144972 7812
rect 260656 7760 260708 7812
rect 34796 7692 34848 7744
rect 127348 7692 127400 7744
rect 147036 7692 147088 7744
rect 278320 7692 278372 7744
rect 373264 7692 373316 7744
rect 381176 7692 381228 7744
rect 381544 7692 381596 7744
rect 391848 7692 391900 7744
rect 24216 7624 24268 7676
rect 122104 7624 122156 7676
rect 149060 7624 149112 7676
rect 307944 7624 307996 7676
rect 365076 7624 365128 7676
rect 376484 7624 376536 7676
rect 380900 7624 380952 7676
rect 393044 7624 393096 7676
rect 27712 7556 27764 7608
rect 127256 7556 127308 7608
rect 165620 7556 165672 7608
rect 449164 7556 449216 7608
rect 381268 6876 381320 6928
rect 384764 6876 384816 6928
rect 140780 6808 140832 6860
rect 203892 6808 203944 6860
rect 162308 6740 162360 6792
rect 235816 6740 235868 6792
rect 160928 6672 160980 6724
rect 271236 6672 271288 6724
rect 104532 6604 104584 6656
rect 132684 6604 132736 6656
rect 146944 6604 146996 6656
rect 270040 6604 270092 6656
rect 80888 6536 80940 6588
rect 131488 6536 131540 6588
rect 146852 6536 146904 6588
rect 273628 6536 273680 6588
rect 77392 6468 77444 6520
rect 131396 6468 131448 6520
rect 146760 6468 146812 6520
rect 276020 6468 276072 6520
rect 313924 6468 313976 6520
rect 322756 6468 322808 6520
rect 66720 6400 66772 6452
rect 130016 6400 130068 6452
rect 146576 6400 146628 6452
rect 277124 6400 277176 6452
rect 307024 6400 307076 6452
rect 329196 6400 329248 6452
rect 44272 6332 44324 6384
rect 128820 6332 128872 6384
rect 146668 6332 146720 6384
rect 279516 6332 279568 6384
rect 298744 6332 298796 6384
rect 320916 6332 320968 6384
rect 392584 6332 392636 6384
rect 398104 6332 398156 6384
rect 33600 6264 33652 6316
rect 127164 6264 127216 6316
rect 151820 6264 151872 6316
rect 348056 6264 348108 6316
rect 373356 6264 373408 6316
rect 378048 6264 378100 6316
rect 381728 6264 381780 6316
rect 395252 6264 395304 6316
rect 19432 6196 19484 6248
rect 124956 6196 125008 6248
rect 161756 6196 161808 6248
rect 471060 6196 471112 6248
rect 18236 6128 18288 6180
rect 126060 6128 126112 6180
rect 137100 6128 137152 6180
rect 145932 6128 145984 6180
rect 171048 6128 171100 6180
rect 576308 6128 576360 6180
rect 313096 5516 313148 5568
rect 314660 5516 314712 5568
rect 376024 5516 376076 5568
rect 378876 5516 378928 5568
rect 384304 5516 384356 5568
rect 387156 5516 387208 5568
rect 114008 5312 114060 5364
rect 134064 5312 134116 5364
rect 101036 5244 101088 5296
rect 133236 5244 133288 5296
rect 136916 5244 136968 5296
rect 154212 5244 154264 5296
rect 93952 5176 94004 5228
rect 133144 5176 133196 5228
rect 137008 5176 137060 5228
rect 157800 5176 157852 5228
rect 63224 5108 63276 5160
rect 129924 5108 129976 5160
rect 138296 5108 138348 5160
rect 169576 5108 169628 5160
rect 30104 5040 30156 5092
rect 127808 5040 127860 5092
rect 136824 5040 136876 5092
rect 148324 5040 148376 5092
rect 154396 5040 154448 5092
rect 213092 5040 213144 5092
rect 15936 4972 15988 5024
rect 113824 4972 113876 5024
rect 142160 4972 142212 5024
rect 216864 4972 216916 5024
rect 436836 4972 436888 5024
rect 28908 4904 28960 4956
rect 127900 4904 127952 4956
rect 148692 4904 148744 4956
rect 294880 4904 294932 4956
rect 479340 4904 479392 4956
rect 6460 4836 6512 4888
rect 10324 4836 10376 4888
rect 13544 4836 13596 4888
rect 125968 4836 126020 4888
rect 138204 4836 138256 4888
rect 162492 4836 162544 4888
rect 162860 4836 162912 4888
rect 487620 4836 487672 4888
rect 8760 4768 8812 4820
rect 125876 4768 125928 4820
rect 138112 4768 138164 4820
rect 166080 4768 166132 4820
rect 169484 4768 169536 4820
rect 562048 4768 562100 4820
rect 136732 4428 136784 4480
rect 144736 4428 144788 4480
rect 184940 4156 184992 4208
rect 186136 4156 186188 4208
rect 201500 4156 201552 4208
rect 202696 4156 202748 4208
rect 242900 4156 242952 4208
rect 244096 4156 244148 4208
rect 251180 4156 251232 4208
rect 252376 4156 252428 4208
rect 572 4088 624 4140
rect 7564 4088 7616 4140
rect 11152 4088 11204 4140
rect 126428 4088 126480 4140
rect 144368 4088 144420 4140
rect 153016 4088 153068 4140
rect 172336 4088 172388 4140
rect 288992 4088 289044 4140
rect 87972 3952 88024 4004
rect 124864 4020 124916 4072
rect 125876 4020 125928 4072
rect 134524 4020 134576 4072
rect 146484 4020 146536 4072
rect 268844 4020 268896 4072
rect 124680 3952 124732 4004
rect 134616 3952 134668 4004
rect 138940 3952 138992 4004
rect 143540 3952 143592 4004
rect 146392 3952 146444 4004
rect 272432 3952 272484 4004
rect 314660 3952 314712 4004
rect 324412 3952 324464 4004
rect 86868 3884 86920 3936
rect 131212 3884 131264 3936
rect 144460 3884 144512 3936
rect 156604 3884 156656 3936
rect 163780 3884 163832 3936
rect 303160 3884 303212 3936
rect 312544 3884 312596 3936
rect 322112 3884 322164 3936
rect 83280 3816 83332 3868
rect 131948 3816 132000 3868
rect 142804 3816 142856 3868
rect 163688 3816 163740 3868
rect 173624 3816 173676 3868
rect 212172 3816 212224 3868
rect 213092 3816 213144 3868
rect 364616 3816 364668 3868
rect 367744 3816 367796 3868
rect 377680 3816 377732 3868
rect 388444 3816 388496 3868
rect 396540 3816 396592 3868
rect 398104 3816 398156 3868
rect 408408 3816 408460 3868
rect 79692 3748 79744 3800
rect 131304 3748 131356 3800
rect 140228 3748 140280 3800
rect 164884 3748 164936 3800
rect 172428 3748 172480 3800
rect 356336 3748 356388 3800
rect 359556 3748 359608 3800
rect 368204 3748 368256 3800
rect 382924 3748 382976 3800
rect 388260 3748 388312 3800
rect 388536 3748 388588 3800
rect 398840 3748 398892 3800
rect 449164 3748 449216 3800
rect 521844 3748 521896 3800
rect 69112 3680 69164 3732
rect 126244 3680 126296 3732
rect 65524 3612 65576 3664
rect 130660 3680 130712 3732
rect 142988 3680 143040 3732
rect 155408 3680 155460 3732
rect 159824 3680 159876 3732
rect 437940 3680 437992 3732
rect 449900 3680 449952 3732
rect 525432 3680 525484 3732
rect 126980 3612 127032 3664
rect 130292 3612 130344 3664
rect 140136 3612 140188 3664
rect 170772 3612 170824 3664
rect 176660 3612 176712 3664
rect 177856 3612 177908 3664
rect 177948 3612 178000 3664
rect 461584 3612 461636 3664
rect 17040 3544 17092 3596
rect 125784 3544 125836 3596
rect 129372 3544 129424 3596
rect 130476 3544 130528 3596
rect 131764 3544 131816 3596
rect 135812 3544 135864 3596
rect 138664 3544 138716 3596
rect 151820 3544 151872 3596
rect 161664 3544 161716 3596
rect 462780 3544 462832 3596
rect 481640 3544 481692 3596
rect 482468 3544 482520 3596
rect 506480 3544 506532 3596
rect 507308 3544 507360 3596
rect 12348 3476 12400 3528
rect 126612 3476 126664 3528
rect 135260 3476 135312 3528
rect 136548 3476 136600 3528
rect 162768 3476 162820 3528
rect 466276 3476 466328 3528
rect 474004 3476 474056 3528
rect 518348 3544 518400 3596
rect 574744 3544 574796 3596
rect 514760 3476 514812 3528
rect 515588 3476 515640 3528
rect 539600 3476 539652 3528
rect 540428 3476 540480 3528
rect 564440 3476 564492 3528
rect 565268 3476 565320 3528
rect 35900 3408 35952 3460
rect 36820 3408 36872 3460
rect 118700 3408 118752 3460
rect 119896 3408 119948 3460
rect 135904 3408 135956 3460
rect 138848 3408 138900 3460
rect 139032 3408 139084 3460
rect 168380 3408 168432 3460
rect 172060 3408 172112 3460
rect 179052 3408 179104 3460
rect 135720 3340 135772 3392
rect 141240 3340 141292 3392
rect 173256 3340 173308 3392
rect 177948 3340 178000 3392
rect 137836 3272 137888 3324
rect 150624 3272 150676 3324
rect 154488 3272 154540 3324
rect 173164 3272 173216 3324
rect 173440 3272 173492 3324
rect 181444 3408 181496 3460
rect 181536 3408 181588 3460
rect 519544 3408 519596 3460
rect 581000 3408 581052 3460
rect 132960 3136 133012 3188
rect 135444 3136 135496 3188
rect 135536 3136 135588 3188
rect 140044 3136 140096 3188
rect 171876 3136 171928 3188
rect 285404 3340 285456 3392
rect 307760 3340 307812 3392
rect 309048 3340 309100 3392
rect 316040 3340 316092 3392
rect 317328 3340 317380 3392
rect 332692 3340 332744 3392
rect 333888 3340 333940 3392
rect 340972 3340 341024 3392
rect 342168 3340 342220 3392
rect 365812 3340 365864 3392
rect 367008 3340 367060 3392
rect 374092 3340 374144 3392
rect 375288 3340 375340 3392
rect 382372 3340 382424 3392
rect 383568 3340 383620 3392
rect 398932 3340 398984 3392
rect 400128 3340 400180 3392
rect 415492 3340 415544 3392
rect 416688 3340 416740 3392
rect 423772 3340 423824 3392
rect 424968 3340 425020 3392
rect 431960 3340 432012 3392
rect 433248 3340 433300 3392
rect 440332 3340 440384 3392
rect 441528 3340 441580 3392
rect 456800 3340 456852 3392
rect 458088 3340 458140 3392
rect 322756 3272 322808 3324
rect 325608 3272 325660 3324
rect 403716 3272 403768 3324
rect 406016 3272 406068 3324
rect 395344 3204 395396 3256
rect 401324 3204 401376 3256
rect 384396 3136 384448 3188
rect 389456 3136 389508 3188
rect 173716 3068 173768 3120
rect 182548 3068 182600 3120
rect 326436 3068 326488 3120
rect 331588 3068 331640 3120
rect 135628 3000 135680 3052
rect 137652 3000 137704 3052
rect 378048 3000 378100 3052
rect 382372 3000 382424 3052
rect 165068 2932 165120 2984
rect 171968 2932 172020 2984
rect 327080 2932 327132 2984
rect 335084 2932 335136 2984
rect 357440 2456 357492 2508
rect 358728 2456 358780 2508
rect 349160 1232 349212 1284
rect 350448 1232 350500 1284
<< metal2 >>
rect 6932 703582 7972 703610
rect 2778 684312 2834 684321
rect 2778 684247 2834 684256
rect 2792 683738 2820 684247
rect 2780 683732 2832 683738
rect 2780 683674 2832 683680
rect 4804 683732 4856 683738
rect 4804 683674 4856 683680
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3054 566944 3110 566953
rect 3054 566879 3110 566888
rect 3068 565894 3096 566879
rect 3056 565888 3108 565894
rect 3056 565830 3108 565836
rect 3238 449576 3294 449585
rect 3238 449511 3294 449520
rect 2962 423600 3018 423609
rect 2962 423535 3018 423544
rect 2976 422346 3004 423535
rect 2964 422340 3016 422346
rect 2964 422282 3016 422288
rect 3054 410544 3110 410553
rect 3054 410479 3110 410488
rect 3068 409902 3096 410479
rect 3056 409896 3108 409902
rect 3056 409838 3108 409844
rect 3054 397488 3110 397497
rect 3054 397423 3110 397432
rect 3068 78849 3096 397423
rect 3252 78985 3280 449511
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 3344 371278 3372 371311
rect 3332 371272 3384 371278
rect 3332 371214 3384 371220
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3344 357474 3372 358391
rect 3332 357468 3384 357474
rect 3332 357410 3384 357416
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3344 318850 3372 319223
rect 3332 318844 3384 318850
rect 3332 318786 3384 318792
rect 3330 306232 3386 306241
rect 3330 306167 3386 306176
rect 3344 305046 3372 306167
rect 3332 305040 3384 305046
rect 3332 304982 3384 304988
rect 3330 267200 3386 267209
rect 3330 267135 3386 267144
rect 3344 266422 3372 267135
rect 3332 266416 3384 266422
rect 3332 266358 3384 266364
rect 3330 254144 3386 254153
rect 3330 254079 3386 254088
rect 3344 253978 3372 254079
rect 3332 253972 3384 253978
rect 3332 253914 3384 253920
rect 3330 241088 3386 241097
rect 3330 241023 3386 241032
rect 3344 240174 3372 241023
rect 3332 240168 3384 240174
rect 3332 240110 3384 240116
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3344 213994 3372 214911
rect 3332 213988 3384 213994
rect 3332 213930 3384 213936
rect 3330 201920 3386 201929
rect 3330 201855 3386 201864
rect 3344 201550 3372 201855
rect 3332 201544 3384 201550
rect 3332 201486 3384 201492
rect 3330 188864 3386 188873
rect 3330 188799 3386 188808
rect 3344 187746 3372 188799
rect 3332 187740 3384 187746
rect 3332 187682 3384 187688
rect 3332 139460 3384 139466
rect 3332 139402 3384 139408
rect 3344 134994 3372 139402
rect 3436 135114 3464 658135
rect 3516 632120 3568 632126
rect 3514 632088 3516 632097
rect 3568 632088 3570 632097
rect 3514 632023 3570 632032
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 618322 3556 619103
rect 3516 618316 3568 618322
rect 3516 618258 3568 618264
rect 3606 606112 3662 606121
rect 3606 606047 3662 606056
rect 3514 580000 3570 580009
rect 3514 579935 3570 579944
rect 3528 579698 3556 579935
rect 3516 579692 3568 579698
rect 3516 579634 3568 579640
rect 3514 527912 3570 527921
rect 3514 527847 3516 527856
rect 3568 527847 3570 527856
rect 3516 527818 3568 527824
rect 3514 514856 3570 514865
rect 3514 514791 3516 514800
rect 3568 514791 3570 514800
rect 3516 514762 3568 514768
rect 3514 475688 3570 475697
rect 3514 475623 3570 475632
rect 3528 474774 3556 475623
rect 3516 474768 3568 474774
rect 3516 474710 3568 474716
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3528 166326 3556 462567
rect 3516 166320 3568 166326
rect 3516 166262 3568 166268
rect 3516 162920 3568 162926
rect 3514 162888 3516 162897
rect 3568 162888 3570 162897
rect 3514 162823 3570 162832
rect 3514 149832 3570 149841
rect 3514 149767 3570 149776
rect 3528 149122 3556 149767
rect 3516 149116 3568 149122
rect 3516 149058 3568 149064
rect 3516 137828 3568 137834
rect 3516 137770 3568 137776
rect 3528 136785 3556 137770
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3424 135108 3476 135114
rect 3424 135050 3476 135056
rect 3344 134966 3556 134994
rect 3424 134904 3476 134910
rect 3424 134846 3476 134852
rect 3332 111784 3384 111790
rect 3332 111726 3384 111732
rect 3344 110673 3372 111726
rect 3330 110664 3386 110673
rect 3330 110599 3386 110608
rect 3436 79121 3464 134846
rect 3528 97617 3556 134966
rect 3514 97608 3570 97617
rect 3514 97543 3570 97552
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 3528 84250 3556 84623
rect 3516 84244 3568 84250
rect 3516 84186 3568 84192
rect 3620 79257 3648 606047
rect 3790 553888 3846 553897
rect 3790 553823 3846 553832
rect 3698 345400 3754 345409
rect 3698 345335 3754 345344
rect 3712 79626 3740 345335
rect 3700 79620 3752 79626
rect 3700 79562 3752 79568
rect 3804 79393 3832 553823
rect 3974 501800 4030 501809
rect 3974 501735 4030 501744
rect 3882 293176 3938 293185
rect 3882 293111 3938 293120
rect 3790 79384 3846 79393
rect 3896 79354 3924 293111
rect 3988 79529 4016 501735
rect 4816 118658 4844 683674
rect 4804 118652 4856 118658
rect 4804 118594 4856 118600
rect 6932 80034 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 7564 632120 7616 632126
rect 7564 632062 7616 632068
rect 7576 120086 7604 632062
rect 17224 579692 17276 579698
rect 17224 579634 17276 579640
rect 8944 527876 8996 527882
rect 8944 527818 8996 527824
rect 7656 136740 7708 136746
rect 7656 136682 7708 136688
rect 7564 120080 7616 120086
rect 7564 120022 7616 120028
rect 6920 80028 6972 80034
rect 6920 79970 6972 79976
rect 3974 79520 4030 79529
rect 3974 79455 4030 79464
rect 3790 79319 3846 79328
rect 3884 79348 3936 79354
rect 3884 79290 3936 79296
rect 3606 79248 3662 79257
rect 3606 79183 3662 79192
rect 3422 79112 3478 79121
rect 3422 79047 3478 79056
rect 3238 78976 3294 78985
rect 3238 78911 3294 78920
rect 3054 78840 3110 78849
rect 3054 78775 3110 78784
rect 6920 76560 6972 76566
rect 6920 76502 6972 76508
rect 2778 75304 2834 75313
rect 2778 75239 2834 75248
rect 1398 75168 1454 75177
rect 1398 75103 1454 75112
rect 572 4140 624 4146
rect 572 4082 624 4088
rect 584 480 612 4082
rect 542 -960 654 480
rect 1412 354 1440 75103
rect 2792 16574 2820 75239
rect 4160 74112 4212 74118
rect 4160 74054 4212 74060
rect 3424 71664 3476 71670
rect 3422 71632 3424 71641
rect 3476 71632 3478 71641
rect 3422 71567 3478 71576
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3424 32564 3476 32570
rect 3424 32506 3476 32512
rect 3436 32473 3464 32506
rect 3422 32464 3478 32473
rect 3422 32399 3478 32408
rect 3332 24336 3384 24342
rect 3332 24278 3384 24284
rect 3344 19417 3372 24278
rect 3424 23248 3476 23254
rect 3424 23190 3476 23196
rect 3330 19408 3386 19417
rect 3330 19343 3386 19352
rect 2792 16546 2912 16574
rect 2884 480 2912 16546
rect 3436 6497 3464 23190
rect 4172 16574 4200 74054
rect 6932 16574 6960 76502
rect 7564 36576 7616 36582
rect 7564 36518 7616 36524
rect 4172 16546 5304 16574
rect 6932 16546 7512 16574
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 4066 4856 4122 4865
rect 4066 4791 4122 4800
rect 4080 480 4108 4791
rect 5276 480 5304 16546
rect 6460 4888 6512 4894
rect 6460 4830 6512 4836
rect 6472 480 6500 4830
rect 7484 3482 7512 16546
rect 7576 4146 7604 36518
rect 7668 32570 7696 136682
rect 8956 122806 8984 527818
rect 10324 474768 10376 474774
rect 10324 474710 10376 474716
rect 9036 135312 9088 135318
rect 9036 135254 9088 135260
rect 8944 122800 8996 122806
rect 8944 122742 8996 122748
rect 9048 71670 9076 135254
rect 10336 124166 10364 474710
rect 13084 422340 13136 422346
rect 13084 422282 13136 422288
rect 13096 126954 13124 422282
rect 14464 318844 14516 318850
rect 14464 318786 14516 318792
rect 14476 129742 14504 318786
rect 14464 129736 14516 129742
rect 14464 129678 14516 129684
rect 13084 126948 13136 126954
rect 13084 126890 13136 126896
rect 10324 124160 10376 124166
rect 10324 124102 10376 124108
rect 17236 121446 17264 579634
rect 18604 266416 18656 266422
rect 18604 266358 18656 266364
rect 18616 131102 18644 266358
rect 21364 162920 21416 162926
rect 21364 162862 21416 162868
rect 21376 133890 21404 162862
rect 23492 145586 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 31024 213988 31076 213994
rect 31024 213930 31076 213936
rect 23480 145580 23532 145586
rect 23480 145522 23532 145528
rect 22744 133952 22796 133958
rect 22744 133894 22796 133900
rect 21364 133884 21416 133890
rect 21364 133826 21416 133832
rect 18604 131096 18656 131102
rect 18604 131038 18656 131044
rect 17224 121440 17276 121446
rect 17224 121382 17276 121388
rect 22756 111790 22784 133894
rect 31036 132462 31064 213930
rect 31024 132456 31076 132462
rect 31024 132398 31076 132404
rect 40052 117298 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 40040 117292 40092 117298
rect 40040 117234 40092 117240
rect 22744 111784 22796 111790
rect 22744 111726 22796 111732
rect 10324 77988 10376 77994
rect 10324 77930 10376 77936
rect 9036 71664 9088 71670
rect 9036 71606 9088 71612
rect 7656 32564 7708 32570
rect 7656 32506 7708 32512
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7484 3454 7696 3482
rect 7668 480 7696 3454
rect 8772 480 8800 4762
rect 9968 480 9996 8910
rect 10336 4894 10364 77930
rect 71792 77217 71820 702986
rect 89180 700330 89208 703520
rect 89168 700324 89220 700330
rect 89168 700266 89220 700272
rect 105464 699718 105492 703520
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106924 699712 106976 699718
rect 106924 699654 106976 699660
rect 84844 371272 84896 371278
rect 84844 371214 84896 371220
rect 82084 240168 82136 240174
rect 82084 240110 82136 240116
rect 82096 79762 82124 240110
rect 84856 128314 84884 371214
rect 84844 128308 84896 128314
rect 84844 128250 84896 128256
rect 106936 115938 106964 699654
rect 120724 616888 120776 616894
rect 120724 616830 120776 616836
rect 118700 431248 118752 431254
rect 118700 431190 118752 431196
rect 118608 404388 118660 404394
rect 118608 404330 118660 404336
rect 118516 351960 118568 351966
rect 118516 351902 118568 351908
rect 118240 142928 118292 142934
rect 118240 142870 118292 142876
rect 118148 141568 118200 141574
rect 118148 141510 118200 141516
rect 118056 141500 118108 141506
rect 118056 141442 118108 141448
rect 117318 137592 117374 137601
rect 117318 137527 117374 137536
rect 117332 136746 117360 137527
rect 117320 136740 117372 136746
rect 117320 136682 117372 136688
rect 117318 136096 117374 136105
rect 117318 136031 117374 136040
rect 117332 135318 117360 136031
rect 117320 135312 117372 135318
rect 117320 135254 117372 135260
rect 117318 134600 117374 134609
rect 117318 134535 117374 134544
rect 117332 133958 117360 134535
rect 117320 133952 117372 133958
rect 117320 133894 117372 133900
rect 117412 133884 117464 133890
rect 117412 133826 117464 133832
rect 117424 133113 117452 133826
rect 117410 133104 117466 133113
rect 117410 133039 117466 133048
rect 117320 132456 117372 132462
rect 117320 132398 117372 132404
rect 117332 131617 117360 132398
rect 117318 131608 117374 131617
rect 117318 131543 117374 131552
rect 117320 131096 117372 131102
rect 117320 131038 117372 131044
rect 117332 130121 117360 131038
rect 117318 130112 117374 130121
rect 117318 130047 117374 130056
rect 117320 129736 117372 129742
rect 117320 129678 117372 129684
rect 117332 128625 117360 129678
rect 117318 128616 117374 128625
rect 117318 128551 117374 128560
rect 117320 128308 117372 128314
rect 117320 128250 117372 128256
rect 117332 127129 117360 128250
rect 117318 127120 117374 127129
rect 117318 127055 117374 127064
rect 117320 126948 117372 126954
rect 117320 126890 117372 126896
rect 117332 125633 117360 126890
rect 117318 125624 117374 125633
rect 117318 125559 117374 125568
rect 117320 124160 117372 124166
rect 117318 124128 117320 124137
rect 117372 124128 117374 124137
rect 117318 124063 117374 124072
rect 117320 122800 117372 122806
rect 117320 122742 117372 122748
rect 117332 122641 117360 122742
rect 117318 122632 117374 122641
rect 117318 122567 117374 122576
rect 117320 121440 117372 121446
rect 117320 121382 117372 121388
rect 117332 121145 117360 121382
rect 117318 121136 117374 121145
rect 117318 121071 117374 121080
rect 117320 120080 117372 120086
rect 117320 120022 117372 120028
rect 117332 119649 117360 120022
rect 117318 119640 117374 119649
rect 117318 119575 117374 119584
rect 117320 118652 117372 118658
rect 117320 118594 117372 118600
rect 117332 118153 117360 118594
rect 117318 118144 117374 118153
rect 117318 118079 117374 118088
rect 117320 117292 117372 117298
rect 117320 117234 117372 117240
rect 117332 116657 117360 117234
rect 117318 116648 117374 116657
rect 117318 116583 117374 116592
rect 106924 115932 106976 115938
rect 106924 115874 106976 115880
rect 117320 115932 117372 115938
rect 117320 115874 117372 115880
rect 117332 115161 117360 115874
rect 117318 115152 117374 115161
rect 117318 115087 117374 115096
rect 118068 113665 118096 141442
rect 118054 113656 118110 113665
rect 118054 113591 118110 113600
rect 118160 91225 118188 141510
rect 118252 92721 118280 142870
rect 118332 139596 118384 139602
rect 118332 139538 118384 139544
rect 118238 92712 118294 92721
rect 118238 92647 118294 92656
rect 118146 91216 118202 91225
rect 118146 91151 118202 91160
rect 118344 89729 118372 139538
rect 118424 139528 118476 139534
rect 118424 139470 118476 139476
rect 118330 89720 118386 89729
rect 118330 89655 118386 89664
rect 118436 88233 118464 139470
rect 118528 94217 118556 351902
rect 118620 95713 118648 404330
rect 118712 103193 118740 431190
rect 119344 187740 119396 187746
rect 119344 187682 119396 187688
rect 119068 145648 119120 145654
rect 119068 145590 119120 145596
rect 118976 142860 119028 142866
rect 118976 142802 119028 142808
rect 118884 141432 118936 141438
rect 118884 141374 118936 141380
rect 118792 140072 118844 140078
rect 118792 140014 118844 140020
rect 118804 104689 118832 140014
rect 118896 106185 118924 141374
rect 118988 107681 119016 142802
rect 119080 112169 119108 145590
rect 119160 144220 119212 144226
rect 119160 144162 119212 144168
rect 119066 112160 119122 112169
rect 119066 112095 119122 112104
rect 119172 110673 119200 144162
rect 119252 140140 119304 140146
rect 119252 140082 119304 140088
rect 119158 110664 119214 110673
rect 119158 110599 119214 110608
rect 119264 109177 119292 140082
rect 119250 109168 119306 109177
rect 119250 109103 119306 109112
rect 118974 107672 119030 107681
rect 118974 107607 119030 107616
rect 118882 106176 118938 106185
rect 118882 106111 118938 106120
rect 118790 104680 118846 104689
rect 118790 104615 118846 104624
rect 118698 103184 118754 103193
rect 118698 103119 118754 103128
rect 118606 95704 118662 95713
rect 118606 95639 118662 95648
rect 118514 94208 118570 94217
rect 118514 94143 118570 94152
rect 118422 88224 118478 88233
rect 118422 88159 118478 88168
rect 118422 86728 118478 86737
rect 118422 86663 118478 86672
rect 118330 82240 118386 82249
rect 118330 82175 118386 82184
rect 82084 79756 82136 79762
rect 82084 79698 82136 79704
rect 116584 78260 116636 78266
rect 116584 78202 116636 78208
rect 113824 78192 113876 78198
rect 113824 78134 113876 78140
rect 93124 78056 93176 78062
rect 93124 77998 93176 78004
rect 71778 77208 71834 77217
rect 71778 77143 71834 77152
rect 70400 76764 70452 76770
rect 70400 76706 70452 76712
rect 37278 76664 37334 76673
rect 37278 76599 37334 76608
rect 69020 76628 69072 76634
rect 20718 76528 20774 76537
rect 20718 76463 20774 76472
rect 13820 51740 13872 51746
rect 13820 51682 13872 51688
rect 13832 16574 13860 51682
rect 20732 16574 20760 76463
rect 26240 75200 26292 75206
rect 26240 75142 26292 75148
rect 22100 22840 22152 22846
rect 22100 22782 22152 22788
rect 22112 16574 22140 22782
rect 13832 16546 14320 16574
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 10324 4888 10376 4894
rect 10324 4830 10376 4836
rect 13544 4888 13596 4894
rect 13544 4830 13596 4836
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 11164 480 11192 4082
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 12360 480 12388 3470
rect 13556 480 13584 4830
rect 1646 354 1758 480
rect 1412 326 1758 354
rect 1646 -960 1758 326
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 19432 6248 19484 6254
rect 19432 6190 19484 6196
rect 18236 6180 18288 6186
rect 18236 6122 18288 6128
rect 15936 5024 15988 5030
rect 15936 4966 15988 4972
rect 15948 480 15976 4966
rect 17040 3596 17092 3602
rect 17040 3538 17092 3544
rect 17052 480 17080 3538
rect 18248 480 18276 6122
rect 19444 480 19472 6190
rect 20626 4992 20682 5001
rect 20626 4927 20682 4936
rect 20640 480 20668 4927
rect 21836 480 21864 16546
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 25320 10396 25372 10402
rect 25320 10338 25372 10344
rect 24216 7676 24268 7682
rect 24216 7618 24268 7624
rect 24228 480 24256 7618
rect 25332 480 25360 10338
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 75142
rect 30380 73908 30432 73914
rect 30380 73850 30432 73856
rect 30392 16574 30420 73850
rect 31760 32428 31812 32434
rect 31760 32370 31812 32376
rect 31772 16574 31800 32370
rect 35900 22908 35952 22914
rect 35900 22850 35952 22856
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 27712 7608 27764 7614
rect 27712 7550 27764 7556
rect 27724 480 27752 7550
rect 30104 5092 30156 5098
rect 30104 5034 30156 5040
rect 28908 4956 28960 4962
rect 28908 4898 28960 4904
rect 28920 480 28948 4898
rect 30116 480 30144 5034
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 34796 7744 34848 7750
rect 34796 7686 34848 7692
rect 33600 6316 33652 6322
rect 33600 6258 33652 6264
rect 33612 480 33640 6258
rect 34808 480 34836 7686
rect 35912 3466 35940 22850
rect 37292 16574 37320 76599
rect 69020 76570 69072 76576
rect 51080 75472 51132 75478
rect 51080 75414 51132 75420
rect 49700 75336 49752 75342
rect 49700 75278 49752 75284
rect 46940 75268 46992 75274
rect 46940 75210 46992 75216
rect 45560 37936 45612 37942
rect 45560 37878 45612 37884
rect 38660 35216 38712 35222
rect 38660 35158 38712 35164
rect 38672 16574 38700 35158
rect 42798 19952 42854 19961
rect 42798 19887 42854 19896
rect 37292 16546 38424 16574
rect 38672 16546 39160 16574
rect 35992 10328 36044 10334
rect 35992 10270 36044 10276
rect 35900 3460 35952 3466
rect 35900 3402 35952 3408
rect 36004 480 36032 10270
rect 36820 3460 36872 3466
rect 36820 3402 36872 3408
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 36832 354 36860 3402
rect 38396 480 38424 16546
rect 37158 354 37270 480
rect 36832 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 41878 8936 41934 8945
rect 41878 8871 41934 8880
rect 40682 6216 40738 6225
rect 40682 6151 40738 6160
rect 40696 480 40724 6151
rect 41892 480 41920 8871
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 39550 -960 39662 326
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 42812 354 42840 19887
rect 45572 16574 45600 37878
rect 46952 16574 46980 75210
rect 49712 16574 49740 75278
rect 45572 16546 46704 16574
rect 46952 16546 47440 16574
rect 49712 16546 50200 16574
rect 45468 9036 45520 9042
rect 45468 8978 45520 8984
rect 44272 6384 44324 6390
rect 44272 6326 44324 6332
rect 44284 480 44312 6326
rect 45480 480 45508 8978
rect 46676 480 46704 16546
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 48964 7812 49016 7818
rect 48964 7754 49016 7760
rect 48976 480 49004 7754
rect 50172 480 50200 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 47830 -960 47942 326
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51092 354 51120 75414
rect 60740 73976 60792 73982
rect 57978 73944 58034 73953
rect 60740 73918 60792 73924
rect 57978 73879 58034 73888
rect 53838 73808 53894 73817
rect 53838 73743 53894 73752
rect 53852 16574 53880 73743
rect 57992 16574 58020 73879
rect 60752 16574 60780 73918
rect 67640 44872 67692 44878
rect 67640 44814 67692 44820
rect 63500 22976 63552 22982
rect 63500 22918 63552 22924
rect 63512 16574 63540 22918
rect 53852 16546 54984 16574
rect 57992 16546 58480 16574
rect 60752 16546 61608 16574
rect 63512 16546 64368 16574
rect 53748 9172 53800 9178
rect 53748 9114 53800 9120
rect 52552 9104 52604 9110
rect 52552 9046 52604 9052
rect 52564 480 52592 9046
rect 53760 480 53788 9114
rect 54956 480 54984 16546
rect 57242 9208 57298 9217
rect 57242 9143 57298 9152
rect 56046 9072 56102 9081
rect 56046 9007 56102 9016
rect 56060 480 56088 9007
rect 57256 480 57284 9143
rect 58452 480 58480 16546
rect 60832 9308 60884 9314
rect 60832 9250 60884 9256
rect 59636 9240 59688 9246
rect 59636 9182 59688 9188
rect 59648 480 59676 9182
rect 60844 480 60872 9250
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61580 354 61608 16546
rect 63224 5160 63276 5166
rect 63224 5102 63276 5108
rect 63236 480 63264 5102
rect 64340 480 64368 16546
rect 66720 6452 66772 6458
rect 66720 6394 66772 6400
rect 65524 3664 65576 3670
rect 65524 3606 65576 3612
rect 65536 480 65564 3606
rect 66732 480 66760 6394
rect 61998 354 62110 480
rect 61580 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67652 354 67680 44814
rect 69032 16574 69060 76570
rect 70412 16574 70440 76706
rect 89718 75576 89774 75585
rect 89718 75511 89774 75520
rect 75918 75440 75974 75449
rect 75918 75375 75974 75384
rect 71778 74080 71834 74089
rect 71778 74015 71834 74024
rect 71792 16574 71820 74015
rect 69032 16546 69888 16574
rect 70412 16546 71544 16574
rect 71792 16546 72648 16574
rect 69112 3732 69164 3738
rect 69112 3674 69164 3680
rect 69124 480 69152 3674
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 16546
rect 71516 480 71544 16546
rect 72620 480 72648 16546
rect 74998 10296 75054 10305
rect 74998 10231 75054 10240
rect 73802 6352 73858 6361
rect 73802 6287 73858 6296
rect 73816 480 73844 6287
rect 75012 480 75040 10231
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 75932 354 75960 75375
rect 88340 55888 88392 55894
rect 88340 55830 88392 55836
rect 85580 21412 85632 21418
rect 85580 21354 85632 21360
rect 81440 18624 81492 18630
rect 81440 18566 81492 18572
rect 81452 16574 81480 18566
rect 85592 16574 85620 21354
rect 88352 16574 88380 55830
rect 89732 16574 89760 75511
rect 91098 44840 91154 44849
rect 91098 44775 91154 44784
rect 91112 16574 91140 44775
rect 81452 16546 81664 16574
rect 85592 16546 85712 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 78128 10464 78180 10470
rect 78128 10406 78180 10412
rect 77392 6520 77444 6526
rect 77392 6462 77444 6468
rect 77404 480 77432 6462
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78140 354 78168 10406
rect 80888 6588 80940 6594
rect 80888 6530 80940 6536
rect 79692 3800 79744 3806
rect 79692 3742 79744 3748
rect 79704 480 79732 3742
rect 80900 480 80928 6530
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 78558 -960 78670 326
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 84476 7880 84528 7886
rect 84476 7822 84528 7828
rect 83280 3868 83332 3874
rect 83280 3810 83332 3816
rect 83292 480 83320 3810
rect 84488 480 84516 7822
rect 85684 480 85712 16546
rect 87972 4004 88024 4010
rect 87972 3946 88024 3952
rect 86868 3936 86920 3942
rect 86868 3878 86920 3884
rect 86880 480 86908 3878
rect 87984 480 88012 3946
rect 89180 480 89208 16546
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 92478 10432 92534 10441
rect 93136 10402 93164 77998
rect 102140 76832 102192 76838
rect 102140 76774 102192 76780
rect 111798 76800 111854 76809
rect 93860 76696 93912 76702
rect 93860 76638 93912 76644
rect 93872 16574 93900 76638
rect 96620 72480 96672 72486
rect 96620 72422 96672 72428
rect 95240 57248 95292 57254
rect 95240 57190 95292 57196
rect 95252 16574 95280 57190
rect 96632 16574 96660 72422
rect 93872 16546 94728 16574
rect 95252 16546 95832 16574
rect 96632 16546 97488 16574
rect 92478 10367 92534 10376
rect 93124 10396 93176 10402
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 10367
rect 93124 10338 93176 10344
rect 93952 5228 94004 5234
rect 93952 5170 94004 5176
rect 93964 480 93992 5170
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94700 354 94728 16546
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95804 354 95832 16546
rect 97460 480 97488 16546
rect 99840 10396 99892 10402
rect 99840 10338 99892 10344
rect 98644 7948 98696 7954
rect 98644 7890 98696 7896
rect 98656 480 98684 7890
rect 99852 480 99880 10338
rect 102152 6914 102180 76774
rect 111798 76735 111854 76744
rect 107660 75404 107712 75410
rect 107660 75346 107712 75352
rect 102232 61396 102284 61402
rect 102232 61338 102284 61344
rect 102244 16574 102272 61338
rect 107672 16574 107700 75346
rect 111812 16574 111840 76735
rect 102244 16546 103376 16574
rect 107672 16546 108160 16574
rect 111812 16546 112392 16574
rect 102152 6886 102272 6914
rect 101036 5296 101088 5302
rect 101036 5238 101088 5244
rect 101048 480 101076 5238
rect 102244 480 102272 6886
rect 103348 480 103376 16546
rect 106464 10532 106516 10538
rect 106464 10474 106516 10480
rect 105728 8016 105780 8022
rect 105728 7958 105780 7964
rect 104532 6656 104584 6662
rect 104532 6598 104584 6604
rect 104544 480 104572 6598
rect 105740 480 105768 7958
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106476 354 106504 10474
rect 108132 480 108160 16546
rect 110510 10568 110566 10577
rect 110510 10503 110566 10512
rect 109314 7576 109370 7585
rect 109314 7511 109370 7520
rect 109328 480 109356 7511
rect 110524 480 110552 10503
rect 111614 7712 111670 7721
rect 111614 7647 111670 7656
rect 111628 480 111656 7647
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 113836 5030 113864 78134
rect 114560 72548 114612 72554
rect 114560 72490 114612 72496
rect 114572 16574 114600 72490
rect 116596 37942 116624 78202
rect 116584 37936 116636 37942
rect 116584 37878 116636 37884
rect 118344 22778 118372 82175
rect 118436 80617 118464 86663
rect 118606 85232 118662 85241
rect 118606 85167 118662 85176
rect 118514 83736 118570 83745
rect 118514 83671 118570 83680
rect 118422 80608 118478 80617
rect 118422 80543 118478 80552
rect 118528 46918 118556 83671
rect 118620 80481 118648 85167
rect 118606 80472 118662 80481
rect 118606 80407 118662 80416
rect 119356 78577 119384 187682
rect 120736 102105 120764 616830
rect 120816 563100 120868 563106
rect 120816 563042 120868 563048
rect 120722 102096 120778 102105
rect 120722 102031 120778 102040
rect 120828 100745 120856 563042
rect 120908 510672 120960 510678
rect 120908 510614 120960 510620
rect 120814 100736 120870 100745
rect 120814 100671 120870 100680
rect 120920 98705 120948 510614
rect 121000 456816 121052 456822
rect 121000 456758 121052 456764
rect 120906 98696 120962 98705
rect 120906 98631 120962 98640
rect 121012 97209 121040 456758
rect 126244 244316 126296 244322
rect 126244 244258 126296 244264
rect 122104 205692 122156 205698
rect 122104 205634 122156 205640
rect 122116 139602 122144 205634
rect 122196 165640 122248 165646
rect 122196 165582 122248 165588
rect 122104 139596 122156 139602
rect 122104 139538 122156 139544
rect 122208 139534 122236 165582
rect 126256 141574 126284 244258
rect 136652 141574 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 702434 154160 703520
rect 170324 702434 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 153212 702406 154160 702434
rect 169772 702406 170352 702434
rect 146944 298172 146996 298178
rect 146944 298114 146996 298120
rect 146956 142934 146984 298114
rect 153212 142934 153240 702406
rect 146944 142928 146996 142934
rect 146944 142870 146996 142876
rect 153200 142928 153252 142934
rect 153200 142870 153252 142876
rect 126244 141568 126296 141574
rect 126244 141510 126296 141516
rect 136640 141568 136692 141574
rect 136640 141510 136692 141516
rect 169772 141506 169800 702406
rect 196624 700664 196676 700670
rect 196624 700606 196676 700612
rect 193864 700596 193916 700602
rect 193864 700538 193916 700544
rect 192484 700528 192536 700534
rect 192484 700470 192536 700476
rect 189724 700460 189776 700466
rect 189724 700402 189776 700408
rect 188344 700392 188396 700398
rect 188344 700334 188396 700340
rect 180800 700324 180852 700330
rect 180800 700266 180852 700272
rect 185584 700324 185636 700330
rect 185584 700266 185636 700272
rect 179420 565888 179472 565894
rect 179420 565830 179472 565836
rect 178684 253972 178736 253978
rect 178684 253914 178736 253920
rect 169760 141500 169812 141506
rect 169760 141442 169812 141448
rect 122196 139528 122248 139534
rect 122196 139470 122248 139476
rect 178696 139398 178724 253914
rect 178776 201544 178828 201550
rect 178776 201486 178828 201492
rect 178684 139392 178736 139398
rect 178684 139334 178736 139340
rect 178788 139330 178816 201486
rect 178776 139324 178828 139330
rect 178776 139266 178828 139272
rect 121092 137828 121144 137834
rect 121092 137770 121144 137776
rect 120998 97200 121054 97209
rect 120998 97135 121054 97144
rect 120724 84244 120776 84250
rect 120724 84186 120776 84192
rect 120736 79286 120764 84186
rect 120908 80844 120960 80850
rect 120908 80786 120960 80792
rect 120920 79762 120948 80786
rect 120908 79756 120960 79762
rect 120908 79698 120960 79704
rect 120724 79280 120776 79286
rect 120724 79222 120776 79228
rect 121104 79218 121132 137770
rect 179432 116657 179460 565830
rect 180064 536852 180116 536858
rect 180064 536794 180116 536800
rect 179512 409896 179564 409902
rect 179512 409838 179564 409844
rect 179524 120737 179552 409838
rect 179696 166320 179748 166326
rect 179696 166262 179748 166268
rect 179604 149116 179656 149122
rect 179604 149058 179656 149064
rect 179616 126857 179644 149058
rect 179602 126848 179658 126857
rect 179602 126783 179658 126792
rect 179510 120728 179566 120737
rect 179510 120663 179566 120672
rect 179708 119377 179736 166262
rect 179788 145580 179840 145586
rect 179788 145522 179840 145528
rect 179694 119368 179750 119377
rect 179694 119303 179750 119312
rect 179418 116648 179474 116657
rect 179418 116583 179474 116592
rect 179800 112577 179828 145522
rect 179878 130520 179934 130529
rect 179878 130455 179934 130464
rect 179786 112568 179842 112577
rect 179786 112503 179842 112512
rect 178592 80776 178644 80782
rect 178592 80718 178644 80724
rect 122104 80640 122156 80646
rect 122104 80582 122156 80588
rect 174728 80640 174780 80646
rect 174728 80582 174780 80588
rect 174820 80640 174872 80646
rect 174820 80582 174872 80588
rect 175004 80640 175056 80646
rect 175004 80582 175056 80588
rect 122116 80034 122144 80582
rect 174452 80436 174504 80442
rect 174452 80378 174504 80384
rect 124678 80200 124734 80209
rect 124678 80135 124734 80144
rect 122104 80028 122156 80034
rect 122104 79970 122156 79976
rect 124404 79348 124456 79354
rect 124404 79290 124456 79296
rect 121092 79212 121144 79218
rect 121092 79154 121144 79160
rect 122196 78600 122248 78606
rect 119342 78568 119398 78577
rect 122196 78542 122248 78548
rect 119342 78503 119398 78512
rect 120724 78328 120776 78334
rect 120724 78270 120776 78276
rect 118700 76900 118752 76906
rect 118700 76842 118752 76848
rect 118516 46912 118568 46918
rect 118516 46854 118568 46860
rect 118332 22772 118384 22778
rect 118332 22714 118384 22720
rect 114572 16546 114784 16574
rect 114008 5364 114060 5370
rect 114008 5306 114060 5312
rect 113824 5024 113876 5030
rect 113824 4966 113876 4972
rect 114020 480 114048 5306
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 117320 10600 117372 10606
rect 117320 10542 117372 10548
rect 116400 8084 116452 8090
rect 116400 8026 116452 8032
rect 116412 480 116440 8026
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 10542
rect 118712 3466 118740 76842
rect 118792 74044 118844 74050
rect 118792 73986 118844 73992
rect 118700 3460 118752 3466
rect 118700 3402 118752 3408
rect 118804 480 118832 73986
rect 120080 59628 120132 59634
rect 120080 59570 120132 59576
rect 120092 16574 120120 59570
rect 120736 32434 120764 78270
rect 122104 77512 122156 77518
rect 122104 77454 122156 77460
rect 121460 75540 121512 75546
rect 121460 75482 121512 75488
rect 120724 32428 120776 32434
rect 120724 32370 120776 32376
rect 120092 16546 120672 16574
rect 119896 3460 119948 3466
rect 119896 3402 119948 3408
rect 119908 480 119936 3402
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 121472 6914 121500 75482
rect 122116 7682 122144 77454
rect 122208 35222 122236 78542
rect 123484 77716 123536 77722
rect 123484 77658 123536 77664
rect 122840 77036 122892 77042
rect 122840 76978 122892 76984
rect 122196 35216 122248 35222
rect 122196 35158 122248 35164
rect 122852 16574 122880 76978
rect 123496 59634 123524 77658
rect 124416 75002 124444 79290
rect 124692 75274 124720 80135
rect 124784 80022 125580 80050
rect 124680 75268 124732 75274
rect 124680 75210 124732 75216
rect 124404 74996 124456 75002
rect 124404 74938 124456 74944
rect 124784 70394 124812 80022
rect 125232 79960 125284 79966
rect 125232 79902 125284 79908
rect 125140 79688 125192 79694
rect 124954 79656 125010 79665
rect 125140 79630 125192 79636
rect 124954 79591 125010 79600
rect 124864 77240 124916 77246
rect 124864 77182 124916 77188
rect 124232 70366 124812 70394
rect 123484 59628 123536 59634
rect 123484 59570 123536 59576
rect 124232 36582 124260 70366
rect 124220 36576 124272 36582
rect 124220 36518 124272 36524
rect 122852 16546 123064 16574
rect 122104 7676 122156 7682
rect 122104 7618 122156 7624
rect 121472 6886 122328 6914
rect 122300 480 122328 6886
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124876 4078 124904 77182
rect 124968 6254 124996 79591
rect 125048 77308 125100 77314
rect 125048 77250 125100 77256
rect 125060 51746 125088 77250
rect 125152 76566 125180 79630
rect 125140 76560 125192 76566
rect 125140 76502 125192 76508
rect 125140 76084 125192 76090
rect 125140 76026 125192 76032
rect 125152 55894 125180 76026
rect 125244 57254 125272 79902
rect 125506 79792 125562 79801
rect 125506 79727 125562 79736
rect 125658 79744 125686 80036
rect 125750 79971 125778 80036
rect 125736 79962 125792 79971
rect 125842 79966 125870 80036
rect 125934 79971 125962 80036
rect 125736 79897 125792 79906
rect 125830 79960 125882 79966
rect 125830 79902 125882 79908
rect 125920 79962 125976 79971
rect 125920 79897 125976 79906
rect 126026 79898 126054 80036
rect 126014 79892 126066 79898
rect 126014 79834 126066 79840
rect 126118 79830 126146 80036
rect 125876 79824 125928 79830
rect 125876 79766 125928 79772
rect 126106 79824 126158 79830
rect 126106 79766 126158 79772
rect 125324 79076 125376 79082
rect 125324 79018 125376 79024
rect 125336 61402 125364 79018
rect 125416 79008 125468 79014
rect 125416 78950 125468 78956
rect 125428 76770 125456 78950
rect 125520 77466 125548 79727
rect 125658 79716 125732 79744
rect 125704 78713 125732 79716
rect 125784 79620 125836 79626
rect 125784 79562 125836 79568
rect 125690 78704 125746 78713
rect 125796 78674 125824 79562
rect 125888 78713 125916 79766
rect 125968 79756 126020 79762
rect 125968 79698 126020 79704
rect 125874 78704 125930 78713
rect 125690 78639 125746 78648
rect 125784 78668 125836 78674
rect 125874 78639 125930 78648
rect 125784 78610 125836 78616
rect 125784 78532 125836 78538
rect 125784 78474 125836 78480
rect 125520 77438 125640 77466
rect 125416 76764 125468 76770
rect 125416 76706 125468 76712
rect 125612 74118 125640 77438
rect 125600 74112 125652 74118
rect 125600 74054 125652 74060
rect 125324 61396 125376 61402
rect 125324 61338 125376 61344
rect 125232 57248 125284 57254
rect 125232 57190 125284 57196
rect 125140 55888 125192 55894
rect 125140 55830 125192 55836
rect 125048 51740 125100 51746
rect 125048 51682 125100 51688
rect 124956 6248 125008 6254
rect 124956 6190 125008 6196
rect 124864 4072 124916 4078
rect 124864 4014 124916 4020
rect 124680 4004 124732 4010
rect 124680 3946 124732 3952
rect 124692 480 124720 3946
rect 125796 3602 125824 78474
rect 125980 77994 126008 79698
rect 126210 79642 126238 80036
rect 126302 79801 126330 80036
rect 126394 79971 126422 80036
rect 126380 79962 126436 79971
rect 126380 79897 126436 79906
rect 126288 79792 126344 79801
rect 126288 79727 126344 79736
rect 126164 79614 126238 79642
rect 126164 78792 126192 79614
rect 126486 79608 126514 80036
rect 126578 79966 126606 80036
rect 126670 79966 126698 80036
rect 126566 79960 126618 79966
rect 126566 79902 126618 79908
rect 126658 79960 126710 79966
rect 126658 79902 126710 79908
rect 126762 79830 126790 80036
rect 126854 79937 126882 80036
rect 126946 79966 126974 80036
rect 127038 79966 127066 80036
rect 127130 79971 127158 80036
rect 126934 79960 126986 79966
rect 126840 79928 126896 79937
rect 126934 79902 126986 79908
rect 127026 79960 127078 79966
rect 127026 79902 127078 79908
rect 127116 79962 127172 79971
rect 127116 79897 127172 79906
rect 126840 79863 126896 79872
rect 126750 79824 126802 79830
rect 126750 79766 126802 79772
rect 126888 79824 126940 79830
rect 126888 79766 126940 79772
rect 126980 79824 127032 79830
rect 126980 79766 127032 79772
rect 127070 79792 127126 79801
rect 126796 79688 126848 79694
rect 126796 79630 126848 79636
rect 126704 79620 126756 79626
rect 126486 79580 126560 79608
rect 126072 78764 126192 78792
rect 125968 77988 126020 77994
rect 125968 77930 126020 77936
rect 126072 75914 126100 78764
rect 126150 78704 126206 78713
rect 126150 78639 126206 78648
rect 126426 78704 126482 78713
rect 126426 78639 126482 78648
rect 125888 75886 126100 75914
rect 125888 4826 125916 75886
rect 125968 75200 126020 75206
rect 125968 75142 126020 75148
rect 125980 4894 126008 75142
rect 126060 75132 126112 75138
rect 126060 75074 126112 75080
rect 126072 6186 126100 75074
rect 126164 8974 126192 78639
rect 126336 73908 126388 73914
rect 126336 73850 126388 73856
rect 126244 73228 126296 73234
rect 126244 73170 126296 73176
rect 126152 8968 126204 8974
rect 126152 8910 126204 8916
rect 126060 6180 126112 6186
rect 126060 6122 126112 6128
rect 125968 4888 126020 4894
rect 125968 4830 126020 4836
rect 125876 4820 125928 4826
rect 125876 4762 125928 4768
rect 125876 4072 125928 4078
rect 125876 4014 125928 4020
rect 125784 3596 125836 3602
rect 125784 3538 125836 3544
rect 125888 480 125916 4014
rect 126256 3738 126284 73170
rect 126348 22982 126376 73850
rect 126336 22976 126388 22982
rect 126336 22918 126388 22924
rect 126440 4146 126468 78639
rect 126532 70394 126560 79580
rect 126704 79562 126756 79568
rect 126612 79552 126664 79558
rect 126612 79494 126664 79500
rect 126624 75206 126652 79494
rect 126716 77314 126744 79562
rect 126808 78198 126836 79630
rect 126796 78192 126848 78198
rect 126796 78134 126848 78140
rect 126796 77988 126848 77994
rect 126796 77930 126848 77936
rect 126704 77308 126756 77314
rect 126704 77250 126756 77256
rect 126612 75200 126664 75206
rect 126612 75142 126664 75148
rect 126808 73914 126836 77930
rect 126900 75138 126928 79766
rect 126992 79665 127020 79766
rect 127222 79778 127250 80036
rect 127314 79937 127342 80036
rect 127406 79966 127434 80036
rect 127498 79966 127526 80036
rect 127394 79960 127446 79966
rect 127300 79928 127356 79937
rect 127394 79902 127446 79908
rect 127486 79960 127538 79966
rect 127590 79937 127618 80036
rect 127682 79966 127710 80036
rect 127774 79966 127802 80036
rect 127866 79966 127894 80036
rect 127958 79971 127986 80036
rect 127670 79960 127722 79966
rect 127486 79902 127538 79908
rect 127576 79928 127632 79937
rect 127300 79863 127356 79872
rect 127670 79902 127722 79908
rect 127762 79960 127814 79966
rect 127762 79902 127814 79908
rect 127854 79960 127906 79966
rect 127854 79902 127906 79908
rect 127944 79962 128000 79971
rect 127944 79897 128000 79906
rect 127576 79863 127632 79872
rect 127808 79824 127860 79830
rect 127070 79727 127126 79736
rect 127176 79750 127250 79778
rect 127714 79792 127770 79801
rect 126978 79656 127034 79665
rect 126978 79591 127034 79600
rect 127084 78538 127112 79727
rect 127176 78826 127204 79750
rect 128050 79812 128078 80036
rect 128142 79971 128170 80036
rect 128128 79962 128184 79971
rect 128128 79897 128184 79906
rect 128234 79898 128262 80036
rect 128326 79966 128354 80036
rect 128418 79966 128446 80036
rect 128314 79960 128366 79966
rect 128314 79902 128366 79908
rect 128406 79960 128458 79966
rect 128406 79902 128458 79908
rect 128222 79892 128274 79898
rect 128222 79834 128274 79840
rect 128050 79784 128170 79812
rect 127808 79766 127860 79772
rect 127714 79727 127770 79736
rect 127530 79656 127586 79665
rect 127348 79620 127400 79626
rect 127530 79591 127586 79600
rect 127348 79562 127400 79568
rect 127176 78798 127296 78826
rect 127164 78736 127216 78742
rect 127164 78678 127216 78684
rect 127072 78532 127124 78538
rect 127072 78474 127124 78480
rect 126980 78396 127032 78402
rect 126980 78338 127032 78344
rect 126888 75132 126940 75138
rect 126888 75074 126940 75080
rect 126796 73908 126848 73914
rect 126796 73850 126848 73856
rect 126532 70366 126652 70394
rect 126428 4140 126480 4146
rect 126428 4082 126480 4088
rect 126244 3732 126296 3738
rect 126244 3674 126296 3680
rect 126624 3534 126652 70366
rect 126992 22914 127020 78338
rect 126980 22908 127032 22914
rect 126980 22850 127032 22856
rect 127176 6322 127204 78678
rect 127268 76537 127296 78798
rect 127360 77518 127388 79562
rect 127440 79552 127492 79558
rect 127440 79494 127492 79500
rect 127452 78062 127480 79494
rect 127440 78056 127492 78062
rect 127440 77998 127492 78004
rect 127348 77512 127400 77518
rect 127348 77454 127400 77460
rect 127254 76528 127310 76537
rect 127254 76463 127310 76472
rect 127440 76356 127492 76362
rect 127440 76298 127492 76304
rect 127256 74996 127308 75002
rect 127256 74938 127308 74944
rect 127268 7614 127296 74938
rect 127348 74724 127400 74730
rect 127348 74666 127400 74672
rect 127360 7750 127388 74666
rect 127452 10334 127480 76298
rect 127544 22846 127572 79591
rect 127624 79552 127676 79558
rect 127624 79494 127676 79500
rect 127636 75002 127664 79494
rect 127728 79354 127756 79727
rect 127716 79348 127768 79354
rect 127716 79290 127768 79296
rect 127624 74996 127676 75002
rect 127624 74938 127676 74944
rect 127532 22840 127584 22846
rect 127532 22782 127584 22788
rect 127622 22672 127678 22681
rect 127622 22607 127678 22616
rect 127636 16574 127664 22607
rect 127636 16546 127756 16574
rect 127440 10328 127492 10334
rect 127440 10270 127492 10276
rect 127348 7744 127400 7750
rect 127348 7686 127400 7692
rect 127256 7608 127308 7614
rect 127256 7550 127308 7556
rect 127164 6316 127216 6322
rect 127164 6258 127216 6264
rect 126980 3664 127032 3670
rect 126980 3606 127032 3612
rect 126612 3528 126664 3534
rect 126612 3470 126664 3476
rect 126992 480 127020 3606
rect 127728 3482 127756 16546
rect 127820 5098 127848 79766
rect 127900 79756 127952 79762
rect 127900 79698 127952 79704
rect 127808 5092 127860 5098
rect 127808 5034 127860 5040
rect 127912 4962 127940 79698
rect 127990 79656 128046 79665
rect 128142 79642 128170 79784
rect 128360 79756 128412 79762
rect 128360 79698 128412 79704
rect 128142 79614 128262 79642
rect 127990 79591 128046 79600
rect 128234 79608 128262 79614
rect 128004 78742 128032 79591
rect 128234 79580 128308 79608
rect 128084 79484 128136 79490
rect 128084 79426 128136 79432
rect 128176 79484 128228 79490
rect 128176 79426 128228 79432
rect 127992 78736 128044 78742
rect 127992 78678 128044 78684
rect 127990 78432 128046 78441
rect 127990 78367 128046 78376
rect 128004 73846 128032 78367
rect 128096 76362 128124 79426
rect 128084 76356 128136 76362
rect 128084 76298 128136 76304
rect 128188 74730 128216 79426
rect 128280 78334 128308 79580
rect 128372 78402 128400 79698
rect 128510 79676 128538 80036
rect 128602 79830 128630 80036
rect 128694 79937 128722 80036
rect 128680 79928 128736 79937
rect 128680 79863 128736 79872
rect 128590 79824 128642 79830
rect 128786 79812 128814 80036
rect 128590 79766 128642 79772
rect 128740 79784 128814 79812
rect 128878 79801 128906 80036
rect 128970 79971 128998 80036
rect 128956 79962 129012 79971
rect 129062 79966 129090 80036
rect 129154 79966 129182 80036
rect 128956 79897 129012 79906
rect 129050 79960 129102 79966
rect 129050 79902 129102 79908
rect 129142 79960 129194 79966
rect 129142 79902 129194 79908
rect 129246 79898 129274 80036
rect 129234 79892 129286 79898
rect 129234 79834 129286 79840
rect 128864 79792 128920 79801
rect 128636 79688 128688 79694
rect 128510 79648 128584 79676
rect 128556 79506 128584 79648
rect 128636 79630 128688 79636
rect 128464 79478 128584 79506
rect 128360 78396 128412 78402
rect 128360 78338 128412 78344
rect 128268 78328 128320 78334
rect 128268 78270 128320 78276
rect 128268 78124 128320 78130
rect 128268 78066 128320 78072
rect 128176 74724 128228 74730
rect 128176 74666 128228 74672
rect 128280 74186 128308 78066
rect 128464 76673 128492 79478
rect 128544 79416 128596 79422
rect 128544 79358 128596 79364
rect 128556 77994 128584 79358
rect 128648 78606 128676 79630
rect 128636 78600 128688 78606
rect 128636 78542 128688 78548
rect 128740 78441 128768 79784
rect 129186 79792 129242 79801
rect 128864 79727 128920 79736
rect 129004 79756 129056 79762
rect 129338 79744 129366 80036
rect 129430 79966 129458 80036
rect 129522 79971 129550 80036
rect 129418 79960 129470 79966
rect 129418 79902 129470 79908
rect 129508 79962 129564 79971
rect 129508 79897 129564 79906
rect 129614 79778 129642 80036
rect 129706 79937 129734 80036
rect 129798 79966 129826 80036
rect 129786 79960 129838 79966
rect 129692 79928 129748 79937
rect 129890 79937 129918 80036
rect 129786 79902 129838 79908
rect 129876 79928 129932 79937
rect 129692 79863 129748 79872
rect 129982 79898 130010 80036
rect 130074 79898 130102 80036
rect 130166 79898 130194 80036
rect 130258 79966 130286 80036
rect 130350 79971 130378 80036
rect 130246 79960 130298 79966
rect 130246 79902 130298 79908
rect 130336 79962 130392 79971
rect 129876 79863 129932 79872
rect 129970 79892 130022 79898
rect 129970 79834 130022 79840
rect 130062 79892 130114 79898
rect 130062 79834 130114 79840
rect 130154 79892 130206 79898
rect 130336 79897 130392 79906
rect 130154 79834 130206 79840
rect 130442 79812 130470 80036
rect 130534 79966 130562 80036
rect 130522 79960 130574 79966
rect 130522 79902 130574 79908
rect 130626 79898 130654 80036
rect 130614 79892 130666 79898
rect 130614 79834 130666 79840
rect 130396 79784 130470 79812
rect 129614 79750 129688 79778
rect 129186 79727 129242 79736
rect 129004 79698 129056 79704
rect 128820 79688 128872 79694
rect 128820 79630 128872 79636
rect 129016 79642 129044 79698
rect 128726 78432 128782 78441
rect 128726 78367 128782 78376
rect 128832 78266 128860 79630
rect 129016 79614 129136 79642
rect 128912 79484 128964 79490
rect 128912 79426 128964 79432
rect 128820 78260 128872 78266
rect 128820 78202 128872 78208
rect 128544 77988 128596 77994
rect 128544 77930 128596 77936
rect 128820 77512 128872 77518
rect 128820 77454 128872 77460
rect 128450 76664 128506 76673
rect 128450 76599 128506 76608
rect 128544 76016 128596 76022
rect 128544 75958 128596 75964
rect 128452 74996 128504 75002
rect 128452 74938 128504 74944
rect 128268 74180 128320 74186
rect 128268 74122 128320 74128
rect 127992 73840 128044 73846
rect 127992 73782 128044 73788
rect 128464 70394 128492 74938
rect 128372 70366 128492 70394
rect 128372 9314 128400 70366
rect 128360 9308 128412 9314
rect 128360 9250 128412 9256
rect 128556 9042 128584 75958
rect 128636 75676 128688 75682
rect 128636 75618 128688 75624
rect 128648 9110 128676 75618
rect 128832 70394 128860 77454
rect 128924 75002 128952 79426
rect 129004 78736 129056 78742
rect 129004 78678 129056 78684
rect 128912 74996 128964 75002
rect 128912 74938 128964 74944
rect 128740 70366 128860 70394
rect 128740 9178 128768 70366
rect 129016 64874 129044 78678
rect 129108 76022 129136 79614
rect 129200 78742 129228 79727
rect 129292 79716 129366 79744
rect 129188 78736 129240 78742
rect 129188 78678 129240 78684
rect 129186 77752 129242 77761
rect 129186 77687 129242 77696
rect 129096 76016 129148 76022
rect 129096 75958 129148 75964
rect 129200 75154 129228 77687
rect 128832 64846 129044 64874
rect 129108 75126 129228 75154
rect 128728 9172 128780 9178
rect 128728 9114 128780 9120
rect 128636 9104 128688 9110
rect 128636 9046 128688 9052
rect 128544 9036 128596 9042
rect 128544 8978 128596 8984
rect 128832 6390 128860 64846
rect 129108 10470 129136 75126
rect 129292 70394 129320 79716
rect 129464 79688 129516 79694
rect 129370 79656 129426 79665
rect 129464 79630 129516 79636
rect 129370 79591 129372 79600
rect 129424 79591 129426 79600
rect 129372 79562 129424 79568
rect 129370 78432 129426 78441
rect 129370 78367 129426 78376
rect 129384 75478 129412 78367
rect 129372 75472 129424 75478
rect 129372 75414 129424 75420
rect 129476 75342 129504 79630
rect 129660 78962 129688 79750
rect 129740 79688 129792 79694
rect 130016 79688 130068 79694
rect 129740 79630 129792 79636
rect 129830 79656 129886 79665
rect 129568 78934 129688 78962
rect 129568 75682 129596 78934
rect 129648 78804 129700 78810
rect 129648 78746 129700 78752
rect 129660 77081 129688 78746
rect 129752 78441 129780 79630
rect 130016 79630 130068 79636
rect 129830 79591 129886 79600
rect 129738 78432 129794 78441
rect 129738 78367 129794 78376
rect 129844 77518 129872 79591
rect 129924 79416 129976 79422
rect 129924 79358 129976 79364
rect 129936 78674 129964 79358
rect 129924 78668 129976 78674
rect 129924 78610 129976 78616
rect 130028 78305 130056 79630
rect 130108 79620 130160 79626
rect 130108 79562 130160 79568
rect 130200 79620 130252 79626
rect 130200 79562 130252 79568
rect 130120 78810 130148 79562
rect 130108 78804 130160 78810
rect 130108 78746 130160 78752
rect 130212 78690 130240 79562
rect 130120 78662 130240 78690
rect 130014 78296 130070 78305
rect 130014 78231 130070 78240
rect 129832 77512 129884 77518
rect 129832 77454 129884 77460
rect 129646 77072 129702 77081
rect 129646 77007 129702 77016
rect 129556 75676 129608 75682
rect 129556 75618 129608 75624
rect 129740 75472 129792 75478
rect 129740 75414 129792 75420
rect 129464 75336 129516 75342
rect 129464 75278 129516 75284
rect 129200 70366 129320 70394
rect 129096 10464 129148 10470
rect 129096 10406 129148 10412
rect 129200 7818 129228 70366
rect 129752 16574 129780 75414
rect 129924 75268 129976 75274
rect 129924 75210 129976 75216
rect 129752 16546 129872 16574
rect 129188 7812 129240 7818
rect 129188 7754 129240 7760
rect 128820 6384 128872 6390
rect 128820 6326 128872 6332
rect 127900 4956 127952 4962
rect 127900 4898 127952 4904
rect 129372 3596 129424 3602
rect 129372 3538 129424 3544
rect 127728 3454 128216 3482
rect 128188 480 128216 3454
rect 129384 480 129412 3538
rect 129844 3482 129872 16546
rect 129936 5166 129964 75210
rect 130016 75200 130068 75206
rect 130016 75142 130068 75148
rect 130028 6458 130056 75142
rect 130120 9246 130148 78662
rect 130198 78432 130254 78441
rect 130198 78367 130254 78376
rect 130212 73982 130240 78367
rect 130292 77172 130344 77178
rect 130292 77114 130344 77120
rect 130200 73976 130252 73982
rect 130200 73918 130252 73924
rect 130304 70394 130332 77114
rect 130396 75274 130424 79784
rect 130718 79744 130746 80036
rect 130810 79966 130838 80036
rect 130902 79966 130930 80036
rect 130798 79960 130850 79966
rect 130798 79902 130850 79908
rect 130890 79960 130942 79966
rect 130890 79902 130942 79908
rect 130994 79898 131022 80036
rect 130982 79892 131034 79898
rect 130982 79834 131034 79840
rect 131086 79778 131114 80036
rect 131178 79966 131206 80036
rect 131270 79966 131298 80036
rect 131166 79960 131218 79966
rect 131166 79902 131218 79908
rect 131258 79960 131310 79966
rect 131258 79902 131310 79908
rect 130936 79756 130988 79762
rect 130672 79716 130746 79744
rect 130856 79716 130936 79744
rect 130476 79688 130528 79694
rect 130476 79630 130528 79636
rect 130488 75914 130516 79630
rect 130568 79552 130620 79558
rect 130568 79494 130620 79500
rect 130580 77178 130608 79494
rect 130568 77172 130620 77178
rect 130568 77114 130620 77120
rect 130488 75886 130608 75914
rect 130476 75744 130528 75750
rect 130476 75686 130528 75692
rect 130384 75268 130436 75274
rect 130384 75210 130436 75216
rect 130382 75168 130438 75177
rect 130382 75103 130438 75112
rect 130212 70366 130332 70394
rect 130212 44878 130240 70366
rect 130200 44872 130252 44878
rect 130200 44814 130252 44820
rect 130108 9240 130160 9246
rect 130108 9182 130160 9188
rect 130396 6914 130424 75103
rect 130304 6886 130424 6914
rect 130016 6452 130068 6458
rect 130016 6394 130068 6400
rect 129924 5160 129976 5166
rect 129924 5102 129976 5108
rect 130304 3670 130332 6886
rect 130292 3664 130344 3670
rect 130292 3606 130344 3612
rect 130488 3602 130516 75686
rect 130580 16574 130608 75886
rect 130672 75206 130700 79716
rect 130752 79552 130804 79558
rect 130752 79494 130804 79500
rect 130764 76634 130792 79494
rect 130752 76628 130804 76634
rect 130752 76570 130804 76576
rect 130660 75200 130712 75206
rect 130660 75142 130712 75148
rect 130856 73234 130884 79716
rect 130936 79698 130988 79704
rect 131040 79750 131114 79778
rect 130936 79484 130988 79490
rect 130936 79426 130988 79432
rect 130948 78305 130976 79426
rect 131040 78878 131068 79750
rect 131362 79744 131390 80036
rect 131454 79966 131482 80036
rect 131546 79966 131574 80036
rect 131442 79960 131494 79966
rect 131442 79902 131494 79908
rect 131534 79960 131586 79966
rect 131638 79937 131666 80036
rect 131534 79902 131586 79908
rect 131624 79928 131680 79937
rect 131624 79863 131680 79872
rect 131442 79824 131494 79830
rect 131316 79716 131390 79744
rect 131440 79792 131442 79801
rect 131494 79792 131496 79801
rect 131730 79744 131758 80036
rect 131822 79830 131850 80036
rect 131914 79830 131942 80036
rect 132006 79966 132034 80036
rect 131994 79960 132046 79966
rect 131994 79902 132046 79908
rect 131810 79824 131862 79830
rect 131810 79766 131862 79772
rect 131902 79824 131954 79830
rect 132098 79812 132126 80036
rect 132190 79966 132218 80036
rect 132178 79960 132230 79966
rect 132178 79902 132230 79908
rect 132282 79898 132310 80036
rect 132374 79937 132402 80036
rect 132360 79928 132416 79937
rect 132270 79892 132322 79898
rect 132360 79863 132416 79872
rect 132270 79834 132322 79840
rect 132098 79784 132218 79812
rect 131902 79766 131954 79772
rect 131440 79727 131496 79736
rect 131684 79716 131758 79744
rect 131120 79688 131172 79694
rect 131120 79630 131172 79636
rect 131210 79656 131266 79665
rect 131028 78872 131080 78878
rect 131028 78814 131080 78820
rect 131132 78441 131160 79630
rect 131210 79591 131266 79600
rect 131118 78432 131174 78441
rect 131118 78367 131174 78376
rect 130934 78296 130990 78305
rect 130934 78231 130990 78240
rect 131224 77246 131252 79591
rect 131316 78033 131344 79716
rect 131684 79626 131712 79716
rect 132040 79688 132092 79694
rect 132190 79676 132218 79784
rect 132466 79778 132494 80036
rect 132558 79971 132586 80036
rect 132544 79962 132600 79971
rect 132544 79897 132600 79906
rect 132650 79898 132678 80036
rect 132638 79892 132690 79898
rect 132638 79834 132690 79840
rect 132742 79830 132770 80036
rect 132316 79756 132368 79762
rect 132316 79698 132368 79704
rect 132420 79750 132494 79778
rect 132730 79824 132782 79830
rect 132730 79766 132782 79772
rect 132040 79630 132092 79636
rect 132144 79648 132218 79676
rect 131396 79620 131448 79626
rect 131396 79562 131448 79568
rect 131672 79620 131724 79626
rect 131672 79562 131724 79568
rect 131764 79620 131816 79626
rect 131764 79562 131816 79568
rect 131302 78024 131358 78033
rect 131302 77959 131358 77968
rect 131212 77240 131264 77246
rect 131212 77182 131264 77188
rect 131212 75336 131264 75342
rect 131212 75278 131264 75284
rect 130844 73228 130896 73234
rect 130844 73170 130896 73176
rect 130580 16546 130700 16574
rect 130672 3738 130700 16546
rect 131224 3942 131252 75278
rect 131304 75200 131356 75206
rect 131304 75142 131356 75148
rect 131212 3936 131264 3942
rect 131212 3878 131264 3884
rect 131316 3806 131344 75142
rect 131408 6526 131436 79562
rect 131580 79552 131632 79558
rect 131580 79494 131632 79500
rect 131488 75268 131540 75274
rect 131488 75210 131540 75216
rect 131500 6594 131528 75210
rect 131592 75206 131620 79494
rect 131672 79484 131724 79490
rect 131672 79426 131724 79432
rect 131580 75200 131632 75206
rect 131580 75142 131632 75148
rect 131580 75064 131632 75070
rect 131580 75006 131632 75012
rect 131592 7886 131620 75006
rect 131684 18630 131712 79426
rect 131776 78112 131804 79562
rect 131776 78084 131896 78112
rect 131764 77988 131816 77994
rect 131764 77930 131816 77936
rect 131776 21418 131804 77930
rect 131868 75274 131896 78084
rect 132052 75914 132080 79630
rect 131960 75886 132080 75914
rect 131856 75268 131908 75274
rect 131856 75210 131908 75216
rect 131764 21412 131816 21418
rect 131764 21354 131816 21360
rect 131672 18624 131724 18630
rect 131672 18566 131724 18572
rect 131580 7880 131632 7886
rect 131580 7822 131632 7828
rect 131488 6588 131540 6594
rect 131488 6530 131540 6536
rect 131396 6520 131448 6526
rect 131396 6462 131448 6468
rect 131960 3874 131988 75886
rect 132144 75070 132172 79648
rect 132224 79552 132276 79558
rect 132224 79494 132276 79500
rect 132236 77994 132264 79494
rect 132224 77988 132276 77994
rect 132224 77930 132276 77936
rect 132328 75342 132356 79698
rect 132420 76090 132448 79750
rect 132834 79744 132862 80036
rect 132926 79966 132954 80036
rect 133018 79966 133046 80036
rect 132914 79960 132966 79966
rect 132914 79902 132966 79908
rect 133006 79960 133058 79966
rect 133006 79902 133058 79908
rect 132960 79824 133012 79830
rect 132960 79766 133012 79772
rect 132834 79716 132908 79744
rect 132500 79688 132552 79694
rect 132500 79630 132552 79636
rect 132684 79688 132736 79694
rect 132684 79630 132736 79636
rect 132512 76702 132540 79630
rect 132592 78804 132644 78810
rect 132592 78746 132644 78752
rect 132500 76696 132552 76702
rect 132500 76638 132552 76644
rect 132408 76084 132460 76090
rect 132408 76026 132460 76032
rect 132316 75336 132368 75342
rect 132316 75278 132368 75284
rect 132132 75064 132184 75070
rect 132132 75006 132184 75012
rect 132604 72486 132632 78746
rect 132696 78033 132724 79630
rect 132776 79620 132828 79626
rect 132776 79562 132828 79568
rect 132788 78946 132816 79562
rect 132776 78940 132828 78946
rect 132776 78882 132828 78888
rect 132776 78736 132828 78742
rect 132776 78678 132828 78684
rect 132682 78024 132738 78033
rect 132682 77959 132738 77968
rect 132684 75268 132736 75274
rect 132684 75210 132736 75216
rect 132592 72480 132644 72486
rect 132592 72422 132644 72428
rect 132696 6662 132724 75210
rect 132788 7954 132816 78678
rect 132880 78674 132908 79716
rect 132868 78668 132920 78674
rect 132868 78610 132920 78616
rect 132868 77444 132920 77450
rect 132868 77386 132920 77392
rect 132880 8022 132908 77386
rect 132972 75834 133000 79766
rect 133110 79744 133138 80036
rect 133202 79778 133230 80036
rect 133294 79898 133322 80036
rect 133386 79966 133414 80036
rect 133478 79966 133506 80036
rect 133570 79966 133598 80036
rect 133374 79960 133426 79966
rect 133374 79902 133426 79908
rect 133466 79960 133518 79966
rect 133466 79902 133518 79908
rect 133558 79960 133610 79966
rect 133558 79902 133610 79908
rect 133282 79892 133334 79898
rect 133282 79834 133334 79840
rect 133512 79824 133564 79830
rect 133202 79750 133276 79778
rect 133662 79812 133690 80036
rect 133512 79766 133564 79772
rect 133616 79784 133690 79812
rect 133064 79716 133138 79744
rect 133064 78810 133092 79716
rect 133144 79552 133196 79558
rect 133144 79494 133196 79500
rect 133052 78804 133104 78810
rect 133052 78746 133104 78752
rect 133052 78668 133104 78674
rect 133052 78610 133104 78616
rect 133064 75914 133092 78610
rect 133156 77897 133184 79494
rect 133248 78742 133276 79750
rect 133420 79756 133472 79762
rect 133420 79698 133472 79704
rect 133328 79688 133380 79694
rect 133328 79630 133380 79636
rect 133236 78736 133288 78742
rect 133236 78678 133288 78684
rect 133236 77988 133288 77994
rect 133236 77930 133288 77936
rect 133142 77888 133198 77897
rect 133142 77823 133198 77832
rect 133064 75886 133184 75914
rect 132972 75806 133092 75834
rect 132960 75132 133012 75138
rect 132960 75074 133012 75080
rect 132972 10402 133000 75074
rect 133064 10538 133092 75806
rect 133052 10532 133104 10538
rect 133052 10474 133104 10480
rect 132960 10396 133012 10402
rect 132960 10338 133012 10344
rect 132868 8016 132920 8022
rect 132868 7958 132920 7964
rect 132776 7948 132828 7954
rect 132776 7890 132828 7896
rect 132684 6656 132736 6662
rect 132684 6598 132736 6604
rect 133156 5234 133184 75886
rect 133248 5302 133276 77930
rect 133340 75138 133368 79630
rect 133432 77994 133460 79698
rect 133420 77988 133472 77994
rect 133420 77930 133472 77936
rect 133524 76838 133552 79766
rect 133512 76832 133564 76838
rect 133512 76774 133564 76780
rect 133616 75274 133644 79784
rect 133754 79744 133782 80036
rect 133846 79966 133874 80036
rect 133834 79960 133886 79966
rect 133834 79902 133886 79908
rect 133938 79898 133966 80036
rect 133926 79892 133978 79898
rect 133926 79834 133978 79840
rect 133708 79716 133782 79744
rect 133878 79792 133934 79801
rect 134030 79744 134058 80036
rect 134122 79966 134150 80036
rect 134214 79966 134242 80036
rect 134110 79960 134162 79966
rect 134110 79902 134162 79908
rect 134202 79960 134254 79966
rect 134306 79937 134334 80036
rect 134202 79902 134254 79908
rect 134292 79928 134348 79937
rect 134292 79863 134348 79872
rect 134398 79812 134426 80036
rect 134352 79784 134426 79812
rect 134352 79744 134380 79784
rect 134490 79744 134518 80036
rect 133878 79727 133934 79736
rect 133708 77450 133736 79716
rect 133788 79620 133840 79626
rect 133788 79562 133840 79568
rect 133696 77444 133748 77450
rect 133696 77386 133748 77392
rect 133800 75410 133828 79562
rect 133892 76809 133920 79727
rect 133984 79716 134058 79744
rect 134260 79716 134380 79744
rect 134444 79716 134518 79744
rect 134582 79744 134610 80036
rect 134674 79937 134702 80036
rect 134660 79928 134716 79937
rect 134660 79863 134716 79872
rect 134766 79778 134794 80036
rect 134858 79898 134886 80036
rect 134950 79971 134978 80036
rect 134936 79962 134992 79971
rect 134846 79892 134898 79898
rect 134936 79897 134992 79906
rect 134846 79834 134898 79840
rect 134720 79750 134794 79778
rect 135042 79778 135070 80036
rect 135134 79966 135162 80036
rect 135226 79966 135254 80036
rect 135318 79966 135346 80036
rect 135410 79966 135438 80036
rect 135502 79971 135530 80036
rect 135122 79960 135174 79966
rect 135122 79902 135174 79908
rect 135214 79960 135266 79966
rect 135214 79902 135266 79908
rect 135306 79960 135358 79966
rect 135306 79902 135358 79908
rect 135398 79960 135450 79966
rect 135398 79902 135450 79908
rect 135488 79962 135544 79971
rect 135488 79897 135544 79906
rect 135594 79898 135622 80036
rect 135582 79892 135634 79898
rect 135582 79834 135634 79840
rect 135686 79830 135714 80036
rect 135778 79898 135806 80036
rect 135870 79971 135898 80036
rect 135856 79962 135912 79971
rect 135766 79892 135818 79898
rect 135856 79897 135912 79906
rect 135766 79834 135818 79840
rect 135352 79824 135404 79830
rect 135350 79792 135352 79801
rect 135674 79824 135726 79830
rect 135404 79792 135406 79801
rect 134892 79756 134944 79762
rect 134582 79716 134656 79744
rect 133878 76800 133934 76809
rect 133878 76735 133934 76744
rect 133880 76016 133932 76022
rect 133880 75958 133932 75964
rect 133788 75404 133840 75410
rect 133788 75346 133840 75352
rect 133604 75268 133656 75274
rect 133604 75210 133656 75216
rect 133328 75132 133380 75138
rect 133328 75074 133380 75080
rect 133236 5296 133288 5302
rect 133236 5238 133288 5244
rect 133144 5228 133196 5234
rect 133144 5170 133196 5176
rect 131948 3868 132000 3874
rect 131948 3810 132000 3816
rect 131304 3800 131356 3806
rect 131304 3742 131356 3748
rect 130660 3732 130712 3738
rect 130660 3674 130712 3680
rect 130476 3596 130528 3602
rect 130476 3538 130528 3544
rect 131764 3596 131816 3602
rect 131764 3538 131816 3544
rect 129844 3454 130608 3482
rect 130580 480 130608 3454
rect 131776 480 131804 3538
rect 132960 3188 133012 3194
rect 132960 3130 133012 3136
rect 132972 480 133000 3130
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 133892 354 133920 75958
rect 133984 75313 134012 79716
rect 134064 79620 134116 79626
rect 134064 79562 134116 79568
rect 134076 77897 134104 79562
rect 134156 79552 134208 79558
rect 134156 79494 134208 79500
rect 134168 78033 134196 79494
rect 134154 78024 134210 78033
rect 134154 77959 134210 77968
rect 134062 77888 134118 77897
rect 134062 77823 134118 77832
rect 134260 75914 134288 79716
rect 134338 79656 134394 79665
rect 134338 79591 134394 79600
rect 134076 75886 134288 75914
rect 133970 75304 134026 75313
rect 133970 75239 134026 75248
rect 134076 5370 134104 75886
rect 134156 75404 134208 75410
rect 134156 75346 134208 75352
rect 134168 8090 134196 75346
rect 134352 70394 134380 79591
rect 134444 72554 134472 79716
rect 134524 79620 134576 79626
rect 134524 79562 134576 79568
rect 134432 72548 134484 72554
rect 134432 72490 134484 72496
rect 134260 70366 134380 70394
rect 134260 10606 134288 70366
rect 134248 10600 134300 10606
rect 134248 10542 134300 10548
rect 134156 8084 134208 8090
rect 134156 8026 134208 8032
rect 134064 5364 134116 5370
rect 134064 5306 134116 5312
rect 134536 4078 134564 79562
rect 134628 75410 134656 79716
rect 134616 75404 134668 75410
rect 134616 75346 134668 75352
rect 134616 75268 134668 75274
rect 134616 75210 134668 75216
rect 134524 4072 134576 4078
rect 134524 4014 134576 4020
rect 134628 4010 134656 75210
rect 134720 74050 134748 79750
rect 135042 79750 135116 79778
rect 134892 79698 134944 79704
rect 134798 79656 134854 79665
rect 134798 79591 134854 79600
rect 134812 77722 134840 79591
rect 134800 77716 134852 77722
rect 134800 77658 134852 77664
rect 134904 77042 134932 79698
rect 134984 79688 135036 79694
rect 134984 79630 135036 79636
rect 134892 77036 134944 77042
rect 134892 76978 134944 76984
rect 134996 76906 135024 79630
rect 134984 76900 135036 76906
rect 134984 76842 135036 76848
rect 135088 75546 135116 79750
rect 135350 79727 135406 79736
rect 135534 79792 135590 79801
rect 135962 79778 135990 80036
rect 136054 79966 136082 80036
rect 136146 79966 136174 80036
rect 136042 79960 136094 79966
rect 136042 79902 136094 79908
rect 136134 79960 136186 79966
rect 136134 79902 136186 79908
rect 136238 79778 136266 80036
rect 136330 79966 136358 80036
rect 136318 79960 136370 79966
rect 136422 79937 136450 80036
rect 136318 79902 136370 79908
rect 136408 79928 136464 79937
rect 136408 79863 136464 79872
rect 135674 79766 135726 79772
rect 135824 79762 135990 79778
rect 135534 79727 135590 79736
rect 135812 79756 135990 79762
rect 135168 79688 135220 79694
rect 135168 79630 135220 79636
rect 135350 79656 135406 79665
rect 135076 75540 135128 75546
rect 135076 75482 135128 75488
rect 135180 75274 135208 79630
rect 135260 79620 135312 79626
rect 135548 79626 135576 79727
rect 135864 79750 135990 79756
rect 136192 79750 136266 79778
rect 135812 79698 135864 79704
rect 135720 79688 135772 79694
rect 135904 79688 135956 79694
rect 135720 79630 135772 79636
rect 135824 79636 135904 79642
rect 135824 79630 135956 79636
rect 135996 79688 136048 79694
rect 135996 79630 136048 79636
rect 135350 79591 135406 79600
rect 135536 79620 135588 79626
rect 135260 79562 135312 79568
rect 135272 75750 135300 79562
rect 135260 75744 135312 75750
rect 135260 75686 135312 75692
rect 135168 75268 135220 75274
rect 135168 75210 135220 75216
rect 134708 74044 134760 74050
rect 134708 73986 134760 73992
rect 135364 70394 135392 79591
rect 135536 79562 135588 79568
rect 135628 79484 135680 79490
rect 135628 79426 135680 79432
rect 135536 79416 135588 79422
rect 135536 79358 135588 79364
rect 135548 79082 135576 79358
rect 135536 79076 135588 79082
rect 135536 79018 135588 79024
rect 135534 78432 135590 78441
rect 135534 78367 135590 78376
rect 135442 78296 135498 78305
rect 135442 78231 135498 78240
rect 135456 75313 135484 78231
rect 135548 76022 135576 78367
rect 135536 76016 135588 76022
rect 135536 75958 135588 75964
rect 135536 75336 135588 75342
rect 135442 75304 135498 75313
rect 135536 75278 135588 75284
rect 135442 75239 135498 75248
rect 135364 70366 135484 70394
rect 134616 4004 134668 4010
rect 134616 3946 134668 3952
rect 135260 3528 135312 3534
rect 135260 3470 135312 3476
rect 135272 480 135300 3470
rect 135456 3194 135484 70366
rect 135548 3194 135576 75278
rect 135444 3188 135496 3194
rect 135444 3130 135496 3136
rect 135536 3188 135588 3194
rect 135536 3130 135588 3136
rect 135640 3058 135668 79426
rect 135732 75478 135760 79630
rect 135824 79614 135944 79630
rect 135720 75472 135772 75478
rect 135720 75414 135772 75420
rect 135720 75200 135772 75206
rect 135720 75142 135772 75148
rect 135732 3398 135760 75142
rect 135824 3602 135852 79614
rect 135904 79552 135956 79558
rect 135904 79494 135956 79500
rect 135812 3596 135864 3602
rect 135812 3538 135864 3544
rect 135916 3466 135944 79494
rect 136008 75914 136036 79630
rect 136088 79620 136140 79626
rect 136088 79562 136140 79568
rect 136100 76090 136128 79562
rect 136192 79490 136220 79750
rect 136514 79744 136542 80036
rect 136606 79971 136634 80036
rect 136592 79962 136648 79971
rect 136698 79966 136726 80036
rect 136790 79966 136818 80036
rect 136592 79897 136648 79906
rect 136686 79960 136738 79966
rect 136686 79902 136738 79908
rect 136778 79960 136830 79966
rect 136778 79902 136830 79908
rect 136882 79898 136910 80036
rect 136974 79971 137002 80036
rect 136960 79962 137016 79971
rect 137066 79966 137094 80036
rect 137158 79966 137186 80036
rect 137250 79966 137278 80036
rect 137342 79966 137370 80036
rect 137434 79966 137462 80036
rect 136870 79892 136922 79898
rect 136960 79897 137016 79906
rect 137054 79960 137106 79966
rect 137054 79902 137106 79908
rect 137146 79960 137198 79966
rect 137146 79902 137198 79908
rect 137238 79960 137290 79966
rect 137238 79902 137290 79908
rect 137330 79960 137382 79966
rect 137330 79902 137382 79908
rect 137422 79960 137474 79966
rect 137422 79902 137474 79908
rect 136870 79834 136922 79840
rect 136732 79824 136784 79830
rect 136732 79766 136784 79772
rect 136468 79716 136542 79744
rect 136270 79656 136326 79665
rect 136270 79591 136326 79600
rect 136180 79484 136232 79490
rect 136180 79426 136232 79432
rect 136180 79348 136232 79354
rect 136180 79290 136232 79296
rect 136192 79150 136220 79290
rect 136180 79144 136232 79150
rect 136180 79086 136232 79092
rect 136088 76084 136140 76090
rect 136088 76026 136140 76032
rect 136008 75886 136128 75914
rect 135996 75268 136048 75274
rect 135996 75210 136048 75216
rect 136008 23458 136036 75210
rect 135996 23452 136048 23458
rect 135996 23394 136048 23400
rect 136100 6914 136128 75886
rect 136284 75342 136312 79591
rect 136468 77294 136496 79716
rect 136546 78432 136602 78441
rect 136546 78367 136602 78376
rect 136376 77266 136496 77294
rect 136272 75336 136324 75342
rect 136272 75278 136324 75284
rect 136376 75206 136404 77266
rect 136456 76084 136508 76090
rect 136456 76026 136508 76032
rect 136364 75200 136416 75206
rect 136364 75142 136416 75148
rect 136468 16574 136496 76026
rect 136560 75274 136588 78367
rect 136548 75268 136600 75274
rect 136548 75210 136600 75216
rect 136468 16546 136588 16574
rect 136100 6886 136496 6914
rect 135904 3460 135956 3466
rect 135904 3402 135956 3408
rect 135720 3392 135772 3398
rect 135720 3334 135772 3340
rect 135628 3052 135680 3058
rect 135628 2994 135680 3000
rect 136468 480 136496 6886
rect 136560 3534 136588 16546
rect 136744 4486 136772 79766
rect 137376 79756 137428 79762
rect 137376 79698 137428 79704
rect 136916 79688 136968 79694
rect 136916 79630 136968 79636
rect 136824 79620 136876 79626
rect 136824 79562 136876 79568
rect 136836 5098 136864 79562
rect 136928 75154 136956 79630
rect 137100 79620 137152 79626
rect 137100 79562 137152 79568
rect 137192 79620 137244 79626
rect 137192 79562 137244 79568
rect 137008 79552 137060 79558
rect 137008 79494 137060 79500
rect 137020 77246 137048 79494
rect 137008 77240 137060 77246
rect 137008 77182 137060 77188
rect 137112 75274 137140 79562
rect 137100 75268 137152 75274
rect 137100 75210 137152 75216
rect 136928 75126 137140 75154
rect 136916 75064 136968 75070
rect 136916 75006 136968 75012
rect 136928 5302 136956 75006
rect 137008 74996 137060 75002
rect 137008 74938 137060 74944
rect 136916 5296 136968 5302
rect 136916 5238 136968 5244
rect 137020 5234 137048 74938
rect 137112 6186 137140 75126
rect 137204 67590 137232 79562
rect 137388 78878 137416 79698
rect 137526 79676 137554 80036
rect 137618 79966 137646 80036
rect 137606 79960 137658 79966
rect 137606 79902 137658 79908
rect 137710 79898 137738 80036
rect 137802 79898 137830 80036
rect 137894 79966 137922 80036
rect 137986 79971 138014 80036
rect 137882 79960 137934 79966
rect 137882 79902 137934 79908
rect 137972 79962 138028 79971
rect 137698 79892 137750 79898
rect 137698 79834 137750 79840
rect 137790 79892 137842 79898
rect 137972 79897 138028 79906
rect 137790 79834 137842 79840
rect 137928 79824 137980 79830
rect 138078 79801 138106 80036
rect 138170 79971 138198 80036
rect 138156 79962 138212 79971
rect 138156 79897 138212 79906
rect 138262 79898 138290 80036
rect 138354 79966 138382 80036
rect 138342 79960 138394 79966
rect 138342 79902 138394 79908
rect 138250 79892 138302 79898
rect 138250 79834 138302 79840
rect 138446 79812 138474 80036
rect 138538 79830 138566 80036
rect 138630 79937 138658 80036
rect 138616 79928 138672 79937
rect 138722 79898 138750 80036
rect 138814 79966 138842 80036
rect 138906 79966 138934 80036
rect 138998 79966 139026 80036
rect 138802 79960 138854 79966
rect 138802 79902 138854 79908
rect 138894 79960 138946 79966
rect 138894 79902 138946 79908
rect 138986 79960 139038 79966
rect 138986 79902 139038 79908
rect 138616 79863 138672 79872
rect 138710 79892 138762 79898
rect 138710 79834 138762 79840
rect 137928 79766 137980 79772
rect 138064 79792 138120 79801
rect 137744 79688 137796 79694
rect 137526 79648 137600 79676
rect 137468 79552 137520 79558
rect 137468 79494 137520 79500
rect 137376 78872 137428 78878
rect 137376 78814 137428 78820
rect 137480 78690 137508 79494
rect 137388 78662 137508 78690
rect 137284 75268 137336 75274
rect 137284 75210 137336 75216
rect 137296 69766 137324 75210
rect 137388 73438 137416 78662
rect 137572 75070 137600 79648
rect 137744 79630 137796 79636
rect 137560 75064 137612 75070
rect 137560 75006 137612 75012
rect 137756 75002 137784 79630
rect 137836 78872 137888 78878
rect 137836 78814 137888 78820
rect 137744 74996 137796 75002
rect 137744 74938 137796 74944
rect 137376 73432 137428 73438
rect 137376 73374 137428 73380
rect 137284 69760 137336 69766
rect 137284 69702 137336 69708
rect 137192 67584 137244 67590
rect 137192 67526 137244 67532
rect 137100 6180 137152 6186
rect 137100 6122 137152 6128
rect 137008 5228 137060 5234
rect 137008 5170 137060 5176
rect 136824 5092 136876 5098
rect 136824 5034 136876 5040
rect 136732 4480 136784 4486
rect 136732 4422 136784 4428
rect 136548 3528 136600 3534
rect 136548 3470 136600 3476
rect 137848 3330 137876 78814
rect 137940 78441 137968 79766
rect 138294 79792 138350 79801
rect 138064 79727 138120 79736
rect 138216 79750 138294 79778
rect 138112 79688 138164 79694
rect 138112 79630 138164 79636
rect 137926 78432 137982 78441
rect 137926 78367 137982 78376
rect 138124 75914 138152 79630
rect 138032 75886 138152 75914
rect 138032 71058 138060 75886
rect 138112 75268 138164 75274
rect 138112 75210 138164 75216
rect 138020 71052 138072 71058
rect 138020 70994 138072 71000
rect 138124 4826 138152 75210
rect 138216 4894 138244 79750
rect 138294 79727 138350 79736
rect 138400 79784 138474 79812
rect 138526 79824 138578 79830
rect 138400 79608 138428 79784
rect 139090 79778 139118 80036
rect 139182 79937 139210 80036
rect 139168 79928 139224 79937
rect 139274 79898 139302 80036
rect 139366 79966 139394 80036
rect 139458 79971 139486 80036
rect 139354 79960 139406 79966
rect 139354 79902 139406 79908
rect 139444 79962 139500 79971
rect 139550 79966 139578 80036
rect 139168 79863 139224 79872
rect 139262 79892 139314 79898
rect 139444 79897 139500 79906
rect 139538 79960 139590 79966
rect 139538 79902 139590 79908
rect 139262 79834 139314 79840
rect 138526 79766 138578 79772
rect 138664 79756 138716 79762
rect 138664 79698 138716 79704
rect 139044 79750 139118 79778
rect 139492 79824 139544 79830
rect 139642 79812 139670 80036
rect 139734 79966 139762 80036
rect 139826 79966 139854 80036
rect 139722 79960 139774 79966
rect 139722 79902 139774 79908
rect 139814 79960 139866 79966
rect 139814 79902 139866 79908
rect 139918 79812 139946 80036
rect 139596 79801 139670 79812
rect 139492 79766 139544 79772
rect 139582 79792 139670 79801
rect 138308 79580 138428 79608
rect 138480 79620 138532 79626
rect 138308 75274 138336 79580
rect 138480 79562 138532 79568
rect 138388 79484 138440 79490
rect 138388 79426 138440 79432
rect 138296 75268 138348 75274
rect 138296 75210 138348 75216
rect 138296 75132 138348 75138
rect 138296 75074 138348 75080
rect 138308 5166 138336 75074
rect 138400 62082 138428 79426
rect 138492 67114 138520 79562
rect 138572 79552 138624 79558
rect 138572 79494 138624 79500
rect 138584 75914 138612 79494
rect 138676 77294 138704 79698
rect 138846 79656 138902 79665
rect 138846 79591 138902 79600
rect 138676 77266 138796 77294
rect 138584 75886 138704 75914
rect 138676 70394 138704 75886
rect 138768 75138 138796 77266
rect 138860 75274 138888 79591
rect 139044 78305 139072 79750
rect 139124 79688 139176 79694
rect 139122 79656 139124 79665
rect 139400 79688 139452 79694
rect 139176 79656 139178 79665
rect 139400 79630 139452 79636
rect 139122 79591 139178 79600
rect 139308 79620 139360 79626
rect 139308 79562 139360 79568
rect 139124 79552 139176 79558
rect 139124 79494 139176 79500
rect 139030 78296 139086 78305
rect 139030 78231 139086 78240
rect 138940 77240 138992 77246
rect 138940 77182 138992 77188
rect 138848 75268 138900 75274
rect 138848 75210 138900 75216
rect 138756 75132 138808 75138
rect 138756 75074 138808 75080
rect 138584 70366 138704 70394
rect 138584 69698 138612 70366
rect 138572 69692 138624 69698
rect 138572 69634 138624 69640
rect 138664 67584 138716 67590
rect 138664 67526 138716 67532
rect 138480 67108 138532 67114
rect 138480 67050 138532 67056
rect 138388 62076 138440 62082
rect 138388 62018 138440 62024
rect 138296 5160 138348 5166
rect 138296 5102 138348 5108
rect 138204 4888 138256 4894
rect 138204 4830 138256 4836
rect 138112 4820 138164 4826
rect 138112 4762 138164 4768
rect 138676 3602 138704 67526
rect 138952 4010 138980 77182
rect 139032 75268 139084 75274
rect 139032 75210 139084 75216
rect 138940 4004 138992 4010
rect 138940 3946 138992 3952
rect 138664 3596 138716 3602
rect 138664 3538 138716 3544
rect 139044 3466 139072 75210
rect 139136 74526 139164 79494
rect 139320 77110 139348 79562
rect 139412 78441 139440 79630
rect 139398 78432 139454 78441
rect 139398 78367 139454 78376
rect 139400 78192 139452 78198
rect 139400 78134 139452 78140
rect 139308 77104 139360 77110
rect 139308 77046 139360 77052
rect 139124 74520 139176 74526
rect 139124 74462 139176 74468
rect 139412 25838 139440 78134
rect 139504 25974 139532 79766
rect 139638 79784 139670 79792
rect 139780 79784 139946 79812
rect 139582 79727 139638 79736
rect 139584 79688 139636 79694
rect 139584 79630 139636 79636
rect 139674 79656 139730 79665
rect 139492 25968 139544 25974
rect 139492 25910 139544 25916
rect 139596 25906 139624 79630
rect 139674 79591 139730 79600
rect 139688 77586 139716 79591
rect 139676 77580 139728 77586
rect 139676 77522 139728 77528
rect 139676 75200 139728 75206
rect 139676 75142 139728 75148
rect 139688 32774 139716 75142
rect 139780 44878 139808 79784
rect 140010 79744 140038 80036
rect 139964 79716 140038 79744
rect 140102 79744 140130 80036
rect 140194 79966 140222 80036
rect 140182 79960 140234 79966
rect 140182 79902 140234 79908
rect 140286 79898 140314 80036
rect 140378 79898 140406 80036
rect 140274 79892 140326 79898
rect 140274 79834 140326 79840
rect 140366 79892 140418 79898
rect 140366 79834 140418 79840
rect 140470 79744 140498 80036
rect 140562 79937 140590 80036
rect 140654 79966 140682 80036
rect 140746 79971 140774 80036
rect 140642 79960 140694 79966
rect 140548 79928 140604 79937
rect 140642 79902 140694 79908
rect 140732 79962 140788 79971
rect 140732 79897 140788 79906
rect 140838 79898 140866 80036
rect 140930 79971 140958 80036
rect 140916 79962 140972 79971
rect 141022 79966 141050 80036
rect 140548 79863 140604 79872
rect 140826 79892 140878 79898
rect 140916 79897 140972 79906
rect 141010 79960 141062 79966
rect 141010 79902 141062 79908
rect 140826 79834 140878 79840
rect 140964 79824 141016 79830
rect 140964 79766 141016 79772
rect 140102 79716 140176 79744
rect 139964 79608 139992 79716
rect 139872 79580 139992 79608
rect 140044 79620 140096 79626
rect 139872 63170 139900 79580
rect 140044 79562 140096 79568
rect 139952 79416 140004 79422
rect 139952 79358 140004 79364
rect 139964 79082 139992 79358
rect 139952 79076 140004 79082
rect 139952 79018 140004 79024
rect 139950 77888 140006 77897
rect 139950 77823 140006 77832
rect 139964 75886 139992 77823
rect 139952 75880 140004 75886
rect 139952 75822 140004 75828
rect 139952 75268 140004 75274
rect 139952 75210 140004 75216
rect 139964 67046 139992 75210
rect 140056 70242 140084 79562
rect 140148 78198 140176 79716
rect 140424 79716 140498 79744
rect 140780 79756 140832 79762
rect 140228 79688 140280 79694
rect 140228 79630 140280 79636
rect 140136 78192 140188 78198
rect 140136 78134 140188 78140
rect 140240 75274 140268 79630
rect 140320 79552 140372 79558
rect 140320 79494 140372 79500
rect 140228 75268 140280 75274
rect 140228 75210 140280 75216
rect 140332 75206 140360 79494
rect 140424 78305 140452 79716
rect 140780 79698 140832 79704
rect 140872 79756 140924 79762
rect 140872 79698 140924 79704
rect 140596 79688 140648 79694
rect 140596 79630 140648 79636
rect 140410 78296 140466 78305
rect 140410 78231 140466 78240
rect 140502 78160 140558 78169
rect 140502 78095 140558 78104
rect 140516 78062 140544 78095
rect 140504 78056 140556 78062
rect 140608 78033 140636 79630
rect 140686 78160 140742 78169
rect 140686 78095 140742 78104
rect 140504 77998 140556 78004
rect 140594 78024 140650 78033
rect 140594 77959 140650 77968
rect 140504 77104 140556 77110
rect 140504 77046 140556 77052
rect 140320 75200 140372 75206
rect 140320 75142 140372 75148
rect 140136 74520 140188 74526
rect 140136 74462 140188 74468
rect 140044 70236 140096 70242
rect 140044 70178 140096 70184
rect 139952 67040 140004 67046
rect 139952 66982 140004 66988
rect 139860 63164 139912 63170
rect 139860 63106 139912 63112
rect 139768 44872 139820 44878
rect 139768 44814 139820 44820
rect 139676 32768 139728 32774
rect 139676 32710 139728 32716
rect 139584 25900 139636 25906
rect 139584 25842 139636 25848
rect 139400 25832 139452 25838
rect 139400 25774 139452 25780
rect 140148 3670 140176 74462
rect 140516 70394 140544 77046
rect 140700 75914 140728 78095
rect 140792 77518 140820 79698
rect 140780 77512 140832 77518
rect 140780 77454 140832 77460
rect 140700 75886 140820 75914
rect 140424 70366 140544 70394
rect 140228 69692 140280 69698
rect 140228 69634 140280 69640
rect 140240 3806 140268 69634
rect 140424 26042 140452 70366
rect 140412 26036 140464 26042
rect 140412 25978 140464 25984
rect 140792 6866 140820 75886
rect 140884 25770 140912 79698
rect 140976 79506 141004 79766
rect 141114 79744 141142 80036
rect 141206 79898 141234 80036
rect 141194 79892 141246 79898
rect 141194 79834 141246 79840
rect 141298 79744 141326 80036
rect 141390 79971 141418 80036
rect 141376 79962 141432 79971
rect 141376 79897 141432 79906
rect 141068 79716 141142 79744
rect 141252 79716 141326 79744
rect 141068 79608 141096 79716
rect 141068 79580 141188 79608
rect 140976 79478 141096 79506
rect 140964 78804 141016 78810
rect 140964 78746 141016 78752
rect 140976 27402 141004 78746
rect 141068 75274 141096 79478
rect 141160 78606 141188 79580
rect 141148 78600 141200 78606
rect 141148 78542 141200 78548
rect 141252 77294 141280 79716
rect 141482 79676 141510 80036
rect 141574 79898 141602 80036
rect 141562 79892 141614 79898
rect 141562 79834 141614 79840
rect 141666 79744 141694 80036
rect 141758 79966 141786 80036
rect 141850 79966 141878 80036
rect 141942 79966 141970 80036
rect 142034 79971 142062 80036
rect 141746 79960 141798 79966
rect 141746 79902 141798 79908
rect 141838 79960 141890 79966
rect 141838 79902 141890 79908
rect 141930 79960 141982 79966
rect 141930 79902 141982 79908
rect 142020 79962 142076 79971
rect 142020 79897 142076 79906
rect 141792 79824 141844 79830
rect 142126 79801 142154 80036
rect 141792 79766 141844 79772
rect 142112 79792 142168 79801
rect 141436 79648 141510 79676
rect 141620 79716 141694 79744
rect 141332 79552 141384 79558
rect 141332 79494 141384 79500
rect 141160 77266 141280 77294
rect 141056 75268 141108 75274
rect 141056 75210 141108 75216
rect 141056 75132 141108 75138
rect 141056 75074 141108 75080
rect 140964 27396 141016 27402
rect 140964 27338 141016 27344
rect 141068 27334 141096 75074
rect 141160 32706 141188 77266
rect 141344 75914 141372 79494
rect 141436 78810 141464 79648
rect 141620 78826 141648 79716
rect 141700 79620 141752 79626
rect 141700 79562 141752 79568
rect 141424 78804 141476 78810
rect 141424 78746 141476 78752
rect 141528 78798 141648 78826
rect 141528 75914 141556 78798
rect 141712 78282 141740 79562
rect 141620 78254 141740 78282
rect 141620 77994 141648 78254
rect 141804 78146 141832 79766
rect 142112 79727 142168 79736
rect 142218 79744 142246 80036
rect 142310 79937 142338 80036
rect 142402 79966 142430 80036
rect 142390 79960 142442 79966
rect 142296 79928 142352 79937
rect 142390 79902 142442 79908
rect 142494 79898 142522 80036
rect 142296 79863 142352 79872
rect 142482 79892 142534 79898
rect 142482 79834 142534 79840
rect 142586 79744 142614 80036
rect 142218 79716 142292 79744
rect 142066 79656 142122 79665
rect 141976 79620 142028 79626
rect 142066 79591 142122 79600
rect 142160 79620 142212 79626
rect 141976 79562 142028 79568
rect 141988 78690 142016 79562
rect 141712 78118 141832 78146
rect 141896 78662 142016 78690
rect 141608 77988 141660 77994
rect 141608 77930 141660 77936
rect 141252 75886 141372 75914
rect 141436 75886 141556 75914
rect 141252 33930 141280 75886
rect 141332 75268 141384 75274
rect 141332 75210 141384 75216
rect 141344 33998 141372 75210
rect 141436 60178 141464 75886
rect 141712 73778 141740 78118
rect 141792 77988 141844 77994
rect 141792 77930 141844 77936
rect 141804 75138 141832 77930
rect 141792 75132 141844 75138
rect 141792 75074 141844 75080
rect 141700 73772 141752 73778
rect 141700 73714 141752 73720
rect 141896 70394 141924 78662
rect 141976 78600 142028 78606
rect 141976 78542 142028 78548
rect 141988 77450 142016 78542
rect 142080 78198 142108 79591
rect 142160 79562 142212 79568
rect 142068 78192 142120 78198
rect 142068 78134 142120 78140
rect 141976 77444 142028 77450
rect 141976 77386 142028 77392
rect 141528 70366 141924 70394
rect 141528 69630 141556 70366
rect 141516 69624 141568 69630
rect 141516 69566 141568 69572
rect 141424 60172 141476 60178
rect 141424 60114 141476 60120
rect 141332 33992 141384 33998
rect 141332 33934 141384 33940
rect 141240 33924 141292 33930
rect 141240 33866 141292 33872
rect 141148 32700 141200 32706
rect 141148 32642 141200 32648
rect 141056 27328 141108 27334
rect 141056 27270 141108 27276
rect 140872 25764 140924 25770
rect 140872 25706 140924 25712
rect 140780 6860 140832 6866
rect 140780 6802 140832 6808
rect 142172 5030 142200 79562
rect 142264 77994 142292 79716
rect 142356 79716 142614 79744
rect 142252 77988 142304 77994
rect 142252 77930 142304 77936
rect 142252 75200 142304 75206
rect 142252 75142 142304 75148
rect 142264 7954 142292 75142
rect 142356 27198 142384 79716
rect 142678 79676 142706 80036
rect 142770 79812 142798 80036
rect 142862 79937 142890 80036
rect 142848 79928 142904 79937
rect 142954 79898 142982 80036
rect 142848 79863 142904 79872
rect 142942 79892 142994 79898
rect 142942 79834 142994 79840
rect 142770 79784 142844 79812
rect 142540 79648 142706 79676
rect 142436 79552 142488 79558
rect 142436 79494 142488 79500
rect 142448 78266 142476 79494
rect 142436 78260 142488 78266
rect 142436 78202 142488 78208
rect 142434 78024 142490 78033
rect 142434 77959 142490 77968
rect 142448 27266 142476 77959
rect 142540 33862 142568 79648
rect 142620 79552 142672 79558
rect 142620 79494 142672 79500
rect 142632 76702 142660 79494
rect 142712 78260 142764 78266
rect 142712 78202 142764 78208
rect 142620 76696 142672 76702
rect 142620 76638 142672 76644
rect 142620 75268 142672 75274
rect 142620 75210 142672 75216
rect 142632 63102 142660 75210
rect 142724 65822 142752 78202
rect 142816 66978 142844 79784
rect 143046 79778 143074 80036
rect 143138 79966 143166 80036
rect 143126 79960 143178 79966
rect 143230 79937 143258 80036
rect 143322 79966 143350 80036
rect 143414 79971 143442 80036
rect 143310 79960 143362 79966
rect 143126 79902 143178 79908
rect 143216 79928 143272 79937
rect 143310 79902 143362 79908
rect 143400 79962 143456 79971
rect 143506 79966 143534 80036
rect 143400 79897 143456 79906
rect 143494 79960 143546 79966
rect 143494 79902 143546 79908
rect 143598 79898 143626 80036
rect 143216 79863 143272 79872
rect 143586 79892 143638 79898
rect 143586 79834 143638 79840
rect 143690 79830 143718 80036
rect 143782 79971 143810 80036
rect 143768 79962 143824 79971
rect 143874 79966 143902 80036
rect 143768 79897 143824 79906
rect 143862 79960 143914 79966
rect 143862 79902 143914 79908
rect 143000 79750 143074 79778
rect 143172 79824 143224 79830
rect 143172 79766 143224 79772
rect 143356 79824 143408 79830
rect 143356 79766 143408 79772
rect 143678 79824 143730 79830
rect 143678 79766 143730 79772
rect 142894 79656 142950 79665
rect 142894 79591 142950 79600
rect 142908 75206 142936 79591
rect 143000 75274 143028 79750
rect 143080 79688 143132 79694
rect 143184 79665 143212 79766
rect 143080 79630 143132 79636
rect 143170 79656 143226 79665
rect 143092 76906 143120 79630
rect 143170 79591 143226 79600
rect 143264 79552 143316 79558
rect 143264 79494 143316 79500
rect 143172 79484 143224 79490
rect 143172 79426 143224 79432
rect 143184 77790 143212 79426
rect 143172 77784 143224 77790
rect 143172 77726 143224 77732
rect 143080 76900 143132 76906
rect 143080 76842 143132 76848
rect 143276 75914 143304 79494
rect 143368 78441 143396 79766
rect 143966 79744 143994 80036
rect 144058 79966 144086 80036
rect 144046 79960 144098 79966
rect 144046 79902 144098 79908
rect 144150 79812 144178 80036
rect 144242 79966 144270 80036
rect 144334 79966 144362 80036
rect 144230 79960 144282 79966
rect 144230 79902 144282 79908
rect 144322 79960 144374 79966
rect 144322 79902 144374 79908
rect 143920 79716 143994 79744
rect 144104 79784 144178 79812
rect 144276 79824 144328 79830
rect 143630 79656 143686 79665
rect 143540 79620 143592 79626
rect 143630 79591 143686 79600
rect 143540 79562 143592 79568
rect 143354 78432 143410 78441
rect 143354 78367 143410 78376
rect 143092 75886 143304 75914
rect 142988 75268 143040 75274
rect 142988 75210 143040 75216
rect 142896 75200 142948 75206
rect 142896 75142 142948 75148
rect 143092 74526 143120 75886
rect 143552 75154 143580 79562
rect 143644 75914 143672 79591
rect 143644 75886 143764 75914
rect 143552 75126 143672 75154
rect 143540 75064 143592 75070
rect 143540 75006 143592 75012
rect 143080 74520 143132 74526
rect 143080 74462 143132 74468
rect 142988 73432 143040 73438
rect 142988 73374 143040 73380
rect 142804 66972 142856 66978
rect 142804 66914 142856 66920
rect 142712 65816 142764 65822
rect 142712 65758 142764 65764
rect 142620 63096 142672 63102
rect 142620 63038 142672 63044
rect 142804 62076 142856 62082
rect 142804 62018 142856 62024
rect 142528 33856 142580 33862
rect 142528 33798 142580 33804
rect 142436 27260 142488 27266
rect 142436 27202 142488 27208
rect 142344 27192 142396 27198
rect 142344 27134 142396 27140
rect 142344 23452 142396 23458
rect 142344 23394 142396 23400
rect 142356 16574 142384 23394
rect 142356 16546 142476 16574
rect 142252 7948 142304 7954
rect 142252 7890 142304 7896
rect 142160 5024 142212 5030
rect 142160 4966 142212 4972
rect 140228 3800 140280 3806
rect 140228 3742 140280 3748
rect 140136 3664 140188 3670
rect 140136 3606 140188 3612
rect 138848 3460 138900 3466
rect 138848 3402 138900 3408
rect 139032 3460 139084 3466
rect 139032 3402 139084 3408
rect 137836 3324 137888 3330
rect 137836 3266 137888 3272
rect 137652 3052 137704 3058
rect 137652 2994 137704 3000
rect 137664 480 137692 2994
rect 138860 480 138888 3402
rect 141240 3392 141292 3398
rect 141240 3334 141292 3340
rect 140044 3188 140096 3194
rect 140044 3130 140096 3136
rect 140056 480 140084 3130
rect 141252 480 141280 3334
rect 142448 480 142476 16546
rect 142816 3874 142844 62018
rect 142804 3868 142856 3874
rect 142804 3810 142856 3816
rect 143000 3738 143028 73374
rect 143552 7886 143580 75006
rect 143644 16182 143672 75126
rect 143736 18902 143764 75886
rect 143816 75336 143868 75342
rect 143816 75278 143868 75284
rect 143828 20194 143856 75278
rect 143920 27130 143948 79716
rect 144000 79552 144052 79558
rect 144000 79494 144052 79500
rect 144012 75914 144040 79494
rect 144104 77294 144132 79784
rect 144276 79766 144328 79772
rect 144104 77266 144224 77294
rect 144012 75886 144132 75914
rect 144000 75200 144052 75206
rect 144000 75142 144052 75148
rect 144012 28626 144040 75142
rect 144104 60110 144132 75886
rect 144196 65754 144224 77266
rect 144288 75342 144316 79766
rect 144426 79744 144454 80036
rect 144518 79966 144546 80036
rect 144506 79960 144558 79966
rect 144506 79902 144558 79908
rect 144506 79824 144558 79830
rect 144380 79716 144454 79744
rect 144504 79792 144506 79801
rect 144558 79792 144560 79801
rect 144504 79727 144560 79736
rect 144276 75336 144328 75342
rect 144276 75278 144328 75284
rect 144380 75070 144408 79716
rect 144610 79676 144638 80036
rect 144702 79966 144730 80036
rect 144794 79966 144822 80036
rect 144886 79971 144914 80036
rect 144690 79960 144742 79966
rect 144690 79902 144742 79908
rect 144782 79960 144834 79966
rect 144782 79902 144834 79908
rect 144872 79962 144928 79971
rect 144872 79897 144928 79906
rect 144978 79898 145006 80036
rect 144966 79892 145018 79898
rect 144966 79834 145018 79840
rect 144826 79792 144882 79801
rect 145070 79778 145098 80036
rect 145162 79898 145190 80036
rect 145150 79892 145202 79898
rect 145150 79834 145202 79840
rect 145254 79778 145282 80036
rect 145346 79898 145374 80036
rect 145438 79966 145466 80036
rect 145530 79966 145558 80036
rect 145622 79971 145650 80036
rect 145426 79960 145478 79966
rect 145426 79902 145478 79908
rect 145518 79960 145570 79966
rect 145518 79902 145570 79908
rect 145608 79962 145664 79971
rect 145714 79966 145742 80036
rect 145806 79966 145834 80036
rect 145334 79892 145386 79898
rect 145608 79897 145664 79906
rect 145702 79960 145754 79966
rect 145702 79902 145754 79908
rect 145794 79960 145846 79966
rect 145794 79902 145846 79908
rect 145334 79834 145386 79840
rect 145898 79812 145926 80036
rect 145990 79898 146018 80036
rect 145978 79892 146030 79898
rect 145978 79834 146030 79840
rect 145852 79801 145926 79812
rect 145838 79792 145926 79801
rect 144826 79727 144882 79736
rect 144920 79756 144972 79762
rect 144458 79656 144514 79665
rect 144610 79648 144684 79676
rect 144458 79591 144460 79600
rect 144512 79591 144514 79600
rect 144460 79562 144512 79568
rect 144552 79348 144604 79354
rect 144552 79290 144604 79296
rect 144460 78668 144512 78674
rect 144460 78610 144512 78616
rect 144472 75206 144500 78610
rect 144564 77194 144592 79290
rect 144656 78441 144684 79648
rect 144840 78674 144868 79727
rect 145070 79750 145144 79778
rect 145254 79750 145328 79778
rect 144920 79698 144972 79704
rect 144828 78668 144880 78674
rect 144828 78610 144880 78616
rect 144642 78432 144698 78441
rect 144642 78367 144698 78376
rect 144932 77738 144960 79698
rect 145012 79688 145064 79694
rect 145012 79630 145064 79636
rect 145024 78266 145052 79630
rect 145012 78260 145064 78266
rect 145012 78202 145064 78208
rect 145012 77852 145064 77858
rect 145012 77794 145064 77800
rect 144840 77710 144960 77738
rect 144840 77314 144868 77710
rect 144920 77648 144972 77654
rect 144920 77590 144972 77596
rect 144828 77308 144880 77314
rect 144828 77250 144880 77256
rect 144564 77166 144684 77194
rect 144552 76696 144604 76702
rect 144552 76638 144604 76644
rect 144460 75200 144512 75206
rect 144460 75142 144512 75148
rect 144368 75064 144420 75070
rect 144368 75006 144420 75012
rect 144564 70394 144592 76638
rect 144380 70366 144592 70394
rect 144656 70394 144684 77166
rect 144656 70366 144776 70394
rect 144184 65748 144236 65754
rect 144184 65690 144236 65696
rect 144092 60104 144144 60110
rect 144092 60046 144144 60052
rect 144000 28620 144052 28626
rect 144000 28562 144052 28568
rect 143908 27124 143960 27130
rect 143908 27066 143960 27072
rect 143816 20188 143868 20194
rect 143816 20130 143868 20136
rect 143724 18896 143776 18902
rect 143724 18838 143776 18844
rect 143632 16176 143684 16182
rect 143632 16118 143684 16124
rect 143540 7880 143592 7886
rect 143540 7822 143592 7828
rect 144380 4146 144408 70366
rect 144748 64874 144776 70366
rect 144472 64846 144776 64874
rect 144368 4140 144420 4146
rect 144368 4082 144420 4088
rect 143540 4004 143592 4010
rect 143540 3946 143592 3952
rect 142988 3732 143040 3738
rect 142988 3674 143040 3680
rect 143552 480 143580 3946
rect 144472 3942 144500 64846
rect 144932 7818 144960 77590
rect 145024 20262 145052 77794
rect 145116 75274 145144 79750
rect 145196 79688 145248 79694
rect 145196 79630 145248 79636
rect 145104 75268 145156 75274
rect 145104 75210 145156 75216
rect 145104 75132 145156 75138
rect 145104 75074 145156 75080
rect 145116 20330 145144 75074
rect 145208 28490 145236 79630
rect 145300 79082 145328 79750
rect 145564 79756 145616 79762
rect 145564 79698 145616 79704
rect 145656 79756 145708 79762
rect 145894 79784 145926 79792
rect 145838 79727 145894 79736
rect 145656 79698 145708 79704
rect 145380 79688 145432 79694
rect 145380 79630 145432 79636
rect 145470 79656 145526 79665
rect 145288 79076 145340 79082
rect 145288 79018 145340 79024
rect 145392 77858 145420 79630
rect 145470 79591 145526 79600
rect 145380 77852 145432 77858
rect 145380 77794 145432 77800
rect 145484 75914 145512 79591
rect 145392 75886 145512 75914
rect 145288 75268 145340 75274
rect 145288 75210 145340 75216
rect 145300 28558 145328 75210
rect 145288 28552 145340 28558
rect 145288 28494 145340 28500
rect 145196 28484 145248 28490
rect 145196 28426 145248 28432
rect 145392 28422 145420 75886
rect 145472 75268 145524 75274
rect 145472 75210 145524 75216
rect 145484 33794 145512 75210
rect 145576 66910 145604 79698
rect 145668 75274 145696 79698
rect 145840 79688 145892 79694
rect 145840 79630 145892 79636
rect 145932 79688 145984 79694
rect 146082 79676 146110 80036
rect 146174 79744 146202 80036
rect 146266 79971 146294 80036
rect 146252 79962 146308 79971
rect 146252 79897 146308 79906
rect 146358 79744 146386 80036
rect 146450 79830 146478 80036
rect 146542 79966 146570 80036
rect 146634 79966 146662 80036
rect 146530 79960 146582 79966
rect 146530 79902 146582 79908
rect 146622 79960 146674 79966
rect 146622 79902 146674 79908
rect 146726 79898 146754 80036
rect 146714 79892 146766 79898
rect 146714 79834 146766 79840
rect 146438 79824 146490 79830
rect 146818 79812 146846 80036
rect 146910 79966 146938 80036
rect 146898 79960 146950 79966
rect 146898 79902 146950 79908
rect 146818 79784 146892 79812
rect 146438 79766 146490 79772
rect 146174 79716 146248 79744
rect 145932 79630 145984 79636
rect 146036 79648 146110 79676
rect 146220 79665 146248 79716
rect 146312 79716 146386 79744
rect 146206 79656 146262 79665
rect 145748 78260 145800 78266
rect 145748 78202 145800 78208
rect 145656 75268 145708 75274
rect 145656 75210 145708 75216
rect 145760 74458 145788 78202
rect 145852 77654 145880 79630
rect 145840 77648 145892 77654
rect 145840 77590 145892 77596
rect 145944 75138 145972 79630
rect 146036 77625 146064 79648
rect 146206 79591 146262 79600
rect 146208 79552 146260 79558
rect 146208 79494 146260 79500
rect 146022 77616 146078 77625
rect 146022 77551 146078 77560
rect 146220 77178 146248 79494
rect 146312 78606 146340 79716
rect 146484 79688 146536 79694
rect 146484 79630 146536 79636
rect 146760 79688 146812 79694
rect 146760 79630 146812 79636
rect 146392 79620 146444 79626
rect 146392 79562 146444 79568
rect 146300 78600 146352 78606
rect 146300 78542 146352 78548
rect 146300 78056 146352 78062
rect 146300 77998 146352 78004
rect 146208 77172 146260 77178
rect 146208 77114 146260 77120
rect 145932 75132 145984 75138
rect 145932 75074 145984 75080
rect 145748 74452 145800 74458
rect 145748 74394 145800 74400
rect 145564 66904 145616 66910
rect 145564 66846 145616 66852
rect 145472 33788 145524 33794
rect 145472 33730 145524 33736
rect 145380 28416 145432 28422
rect 145380 28358 145432 28364
rect 145104 20324 145156 20330
rect 145104 20266 145156 20272
rect 145012 20256 145064 20262
rect 145012 20198 145064 20204
rect 144920 7812 144972 7818
rect 144920 7754 144972 7760
rect 145932 6180 145984 6186
rect 145932 6122 145984 6128
rect 144736 4480 144788 4486
rect 144736 4422 144788 4428
rect 144460 3936 144512 3942
rect 144460 3878 144512 3884
rect 144748 480 144776 4422
rect 145944 480 145972 6122
rect 146312 3482 146340 77998
rect 146404 76809 146432 79562
rect 146390 76800 146446 76809
rect 146390 76735 146446 76744
rect 146392 75268 146444 75274
rect 146392 75210 146444 75216
rect 146404 4010 146432 75210
rect 146496 4078 146524 79630
rect 146576 79620 146628 79626
rect 146576 79562 146628 79568
rect 146668 79620 146720 79626
rect 146668 79562 146720 79568
rect 146588 75138 146616 79562
rect 146680 75274 146708 79562
rect 146772 78538 146800 79630
rect 146760 78532 146812 78538
rect 146760 78474 146812 78480
rect 146668 75268 146720 75274
rect 146668 75210 146720 75216
rect 146760 75268 146812 75274
rect 146760 75210 146812 75216
rect 146576 75132 146628 75138
rect 146576 75074 146628 75080
rect 146668 75064 146720 75070
rect 146668 75006 146720 75012
rect 146576 74996 146628 75002
rect 146576 74938 146628 74944
rect 146588 6458 146616 74938
rect 146576 6452 146628 6458
rect 146576 6394 146628 6400
rect 146680 6390 146708 75006
rect 146772 6526 146800 75210
rect 146864 6594 146892 79784
rect 147002 79744 147030 80036
rect 146956 79716 147030 79744
rect 147094 79744 147122 80036
rect 147186 79898 147214 80036
rect 147278 79898 147306 80036
rect 147370 79966 147398 80036
rect 147462 79971 147490 80036
rect 147358 79960 147410 79966
rect 147358 79902 147410 79908
rect 147448 79962 147504 79971
rect 147174 79892 147226 79898
rect 147174 79834 147226 79840
rect 147266 79892 147318 79898
rect 147448 79897 147504 79906
rect 147266 79834 147318 79840
rect 147310 79792 147366 79801
rect 147094 79716 147260 79744
rect 147310 79727 147366 79736
rect 147554 79744 147582 80036
rect 147646 79937 147674 80036
rect 147632 79928 147688 79937
rect 147738 79898 147766 80036
rect 147632 79863 147688 79872
rect 147726 79892 147778 79898
rect 147726 79834 147778 79840
rect 147830 79801 147858 80036
rect 147922 79830 147950 80036
rect 148014 79830 148042 80036
rect 148106 79830 148134 80036
rect 148198 79971 148226 80036
rect 148184 79962 148240 79971
rect 148184 79897 148240 79906
rect 147910 79824 147962 79830
rect 147816 79792 147872 79801
rect 146956 75274 146984 79716
rect 147128 79620 147180 79626
rect 147128 79562 147180 79568
rect 147036 79552 147088 79558
rect 147036 79494 147088 79500
rect 146944 75268 146996 75274
rect 146944 75210 146996 75216
rect 146944 75132 146996 75138
rect 146944 75074 146996 75080
rect 146956 6662 146984 75074
rect 147048 7750 147076 79494
rect 147140 63034 147168 79562
rect 147232 75002 147260 79716
rect 147324 77110 147352 79727
rect 147554 79716 147720 79744
rect 147910 79766 147962 79772
rect 148002 79824 148054 79830
rect 148002 79766 148054 79772
rect 148094 79824 148146 79830
rect 148094 79766 148146 79772
rect 148290 79778 148318 80036
rect 148382 79898 148410 80036
rect 148370 79892 148422 79898
rect 148370 79834 148422 79840
rect 148290 79750 148364 79778
rect 147816 79727 147872 79736
rect 147496 79620 147548 79626
rect 147496 79562 147548 79568
rect 147588 79620 147640 79626
rect 147588 79562 147640 79568
rect 147312 77104 147364 77110
rect 147312 77046 147364 77052
rect 147508 75070 147536 79562
rect 147600 78441 147628 79562
rect 147586 78432 147642 78441
rect 147586 78367 147642 78376
rect 147692 76673 147720 79716
rect 147954 79656 148010 79665
rect 148138 79656 148194 79665
rect 147954 79591 148010 79600
rect 148048 79620 148100 79626
rect 147772 79552 147824 79558
rect 147772 79494 147824 79500
rect 147784 78674 147812 79494
rect 147864 79484 147916 79490
rect 147864 79426 147916 79432
rect 147772 78668 147824 78674
rect 147772 78610 147824 78616
rect 147678 76664 147734 76673
rect 147678 76599 147734 76608
rect 147772 75200 147824 75206
rect 147772 75142 147824 75148
rect 147496 75064 147548 75070
rect 147496 75006 147548 75012
rect 147220 74996 147272 75002
rect 147220 74938 147272 74944
rect 147128 63028 147180 63034
rect 147128 62970 147180 62976
rect 147784 9654 147812 75142
rect 147876 24682 147904 79426
rect 147968 78656 147996 79591
rect 148138 79591 148194 79600
rect 148048 79562 148100 79568
rect 148060 78810 148088 79562
rect 148152 78826 148180 79591
rect 148048 78804 148100 78810
rect 148152 78798 148272 78826
rect 148048 78746 148100 78752
rect 148140 78668 148192 78674
rect 147968 78628 148088 78656
rect 147954 78432 148010 78441
rect 147954 78367 148010 78376
rect 147968 77042 147996 78367
rect 147956 77036 148008 77042
rect 147956 76978 148008 76984
rect 147956 75268 148008 75274
rect 147956 75210 148008 75216
rect 147968 25702 147996 75210
rect 148060 29918 148088 78628
rect 148140 78610 148192 78616
rect 148152 35358 148180 78610
rect 148140 35352 148192 35358
rect 148140 35294 148192 35300
rect 148244 35290 148272 78798
rect 148336 61606 148364 79750
rect 148474 79676 148502 80036
rect 148566 79898 148594 80036
rect 148658 79971 148686 80036
rect 148644 79962 148700 79971
rect 148554 79892 148606 79898
rect 148644 79897 148700 79906
rect 148554 79834 148606 79840
rect 148750 79778 148778 80036
rect 148842 79937 148870 80036
rect 148828 79928 148884 79937
rect 148828 79863 148884 79872
rect 148750 79750 148824 79778
rect 148692 79688 148744 79694
rect 148474 79648 148548 79676
rect 148416 79552 148468 79558
rect 148416 79494 148468 79500
rect 148428 78946 148456 79494
rect 148416 78940 148468 78946
rect 148416 78882 148468 78888
rect 148416 77784 148468 77790
rect 148416 77726 148468 77732
rect 148428 70990 148456 77726
rect 148416 70984 148468 70990
rect 148416 70926 148468 70932
rect 148520 70394 148548 79648
rect 148692 79630 148744 79636
rect 148600 79620 148652 79626
rect 148600 79562 148652 79568
rect 148612 75274 148640 79562
rect 148600 75268 148652 75274
rect 148600 75210 148652 75216
rect 148704 75206 148732 79630
rect 148796 78033 148824 79750
rect 148934 79744 148962 80036
rect 149026 79966 149054 80036
rect 149014 79960 149066 79966
rect 149014 79902 149066 79908
rect 149118 79830 149146 80036
rect 149106 79824 149158 79830
rect 149106 79766 149158 79772
rect 148888 79716 148962 79744
rect 149210 79744 149238 80036
rect 149302 79937 149330 80036
rect 149288 79928 149344 79937
rect 149394 79898 149422 80036
rect 149486 79898 149514 80036
rect 149578 79937 149606 80036
rect 149564 79928 149620 79937
rect 149288 79863 149344 79872
rect 149382 79892 149434 79898
rect 149382 79834 149434 79840
rect 149474 79892 149526 79898
rect 149564 79863 149620 79872
rect 149474 79834 149526 79840
rect 149670 79744 149698 80036
rect 149762 79971 149790 80036
rect 149748 79962 149804 79971
rect 149748 79897 149804 79906
rect 149854 79898 149882 80036
rect 149946 79898 149974 80036
rect 149842 79892 149894 79898
rect 149842 79834 149894 79840
rect 149934 79892 149986 79898
rect 149934 79834 149986 79840
rect 150038 79830 150066 80036
rect 150130 79971 150158 80036
rect 150116 79962 150172 79971
rect 150116 79897 150172 79906
rect 150222 79835 150250 80036
rect 150314 79966 150342 80036
rect 150302 79960 150354 79966
rect 150302 79902 150354 79908
rect 150406 79898 150434 80036
rect 150498 79971 150526 80036
rect 150484 79962 150540 79971
rect 150590 79966 150618 80036
rect 150394 79892 150446 79898
rect 150484 79897 150540 79906
rect 150578 79960 150630 79966
rect 150578 79902 150630 79908
rect 150682 79898 150710 80036
rect 150774 79966 150802 80036
rect 150866 79966 150894 80036
rect 150958 79966 150986 80036
rect 150762 79960 150814 79966
rect 150762 79902 150814 79908
rect 150854 79960 150906 79966
rect 150854 79902 150906 79908
rect 150946 79960 150998 79966
rect 150946 79902 150998 79908
rect 150026 79824 150078 79830
rect 150026 79766 150078 79772
rect 150208 79826 150264 79835
rect 150394 79834 150446 79840
rect 150670 79892 150722 79898
rect 150670 79834 150722 79840
rect 150208 79761 150264 79770
rect 150854 79824 150906 79830
rect 150854 79766 150906 79772
rect 150440 79756 150492 79762
rect 149210 79716 149284 79744
rect 149670 79716 149744 79744
rect 148888 78305 148916 79716
rect 148968 79620 149020 79626
rect 148968 79562 149020 79568
rect 149060 79620 149112 79626
rect 149060 79562 149112 79568
rect 149152 79620 149204 79626
rect 149152 79562 149204 79568
rect 148980 78334 149008 79562
rect 148968 78328 149020 78334
rect 148874 78296 148930 78305
rect 148968 78270 149020 78276
rect 148874 78231 148930 78240
rect 149072 78169 149100 79562
rect 149058 78160 149114 78169
rect 149058 78095 149114 78104
rect 148782 78024 148838 78033
rect 148782 77959 148838 77968
rect 149060 76424 149112 76430
rect 149060 76366 149112 76372
rect 148692 75200 148744 75206
rect 148692 75142 148744 75148
rect 148520 70366 148732 70394
rect 148324 61600 148376 61606
rect 148324 61542 148376 61548
rect 148232 35284 148284 35290
rect 148232 35226 148284 35232
rect 148048 29912 148100 29918
rect 148048 29854 148100 29860
rect 147956 25696 148008 25702
rect 147956 25638 148008 25644
rect 147864 24676 147916 24682
rect 147864 24618 147916 24624
rect 147772 9648 147824 9654
rect 147772 9590 147824 9596
rect 147036 7744 147088 7750
rect 147036 7686 147088 7692
rect 146944 6656 146996 6662
rect 146944 6598 146996 6604
rect 146852 6588 146904 6594
rect 146852 6530 146904 6536
rect 146760 6520 146812 6526
rect 146760 6462 146812 6468
rect 146668 6384 146720 6390
rect 146668 6326 146720 6332
rect 148324 5092 148376 5098
rect 148324 5034 148376 5040
rect 146484 4072 146536 4078
rect 146484 4014 146536 4020
rect 146392 4004 146444 4010
rect 146392 3946 146444 3952
rect 146312 3454 147168 3482
rect 147140 480 147168 3454
rect 148336 480 148364 5034
rect 148704 4962 148732 70366
rect 149072 7682 149100 76366
rect 149164 75138 149192 79562
rect 149256 76242 149284 79716
rect 149520 79688 149572 79694
rect 149426 79656 149482 79665
rect 149336 79620 149388 79626
rect 149716 79676 149744 79716
rect 150440 79698 150492 79704
rect 150164 79688 150216 79694
rect 149716 79648 149790 79676
rect 149520 79630 149572 79636
rect 149426 79591 149482 79600
rect 149336 79562 149388 79568
rect 149348 77246 149376 79562
rect 149336 77240 149388 77246
rect 149336 77182 149388 77188
rect 149440 76362 149468 79591
rect 149532 76430 149560 79630
rect 149762 79608 149790 79648
rect 150070 79656 150126 79665
rect 149762 79580 149836 79608
rect 150164 79630 150216 79636
rect 150070 79591 150126 79600
rect 149612 79552 149664 79558
rect 149612 79494 149664 79500
rect 149624 78656 149652 79494
rect 149624 78628 149744 78656
rect 149610 78432 149666 78441
rect 149610 78367 149666 78376
rect 149520 76424 149572 76430
rect 149520 76366 149572 76372
rect 149428 76356 149480 76362
rect 149428 76298 149480 76304
rect 149256 76214 149560 76242
rect 149244 75336 149296 75342
rect 149244 75278 149296 75284
rect 149152 75132 149204 75138
rect 149152 75074 149204 75080
rect 149152 69760 149204 69766
rect 149152 69702 149204 69708
rect 149060 7676 149112 7682
rect 149060 7618 149112 7624
rect 149164 6914 149192 69702
rect 149256 10402 149284 75278
rect 149336 75268 149388 75274
rect 149336 75210 149388 75216
rect 149348 10470 149376 75210
rect 149428 75200 149480 75206
rect 149428 75142 149480 75148
rect 149440 14822 149468 75142
rect 149532 27062 149560 76214
rect 149624 60042 149652 78367
rect 149716 61538 149744 78628
rect 149808 75274 149836 79580
rect 149980 79552 150032 79558
rect 149980 79494 150032 79500
rect 149992 78441 150020 79494
rect 149978 78432 150034 78441
rect 149978 78367 150034 78376
rect 150084 78316 150112 79591
rect 149900 78288 150112 78316
rect 149796 75268 149848 75274
rect 149796 75210 149848 75216
rect 149900 75206 149928 78288
rect 150072 77240 150124 77246
rect 150072 77182 150124 77188
rect 149980 76356 150032 76362
rect 149980 76298 150032 76304
rect 149888 75200 149940 75206
rect 149888 75142 149940 75148
rect 149992 72690 150020 76298
rect 149980 72684 150032 72690
rect 149980 72626 150032 72632
rect 150084 72622 150112 77182
rect 150176 75342 150204 79630
rect 150256 79620 150308 79626
rect 150256 79562 150308 79568
rect 150268 78305 150296 79562
rect 150348 79552 150400 79558
rect 150348 79494 150400 79500
rect 150360 78402 150388 79494
rect 150452 78674 150480 79698
rect 150532 79688 150584 79694
rect 150866 79676 150894 79766
rect 151050 79744 151078 80036
rect 151142 79937 151170 80036
rect 151234 79966 151262 80036
rect 151222 79960 151274 79966
rect 151128 79928 151184 79937
rect 151222 79902 151274 79908
rect 151326 79898 151354 80036
rect 151418 79898 151446 80036
rect 151510 79966 151538 80036
rect 151498 79960 151550 79966
rect 151498 79902 151550 79908
rect 151128 79863 151184 79872
rect 151314 79892 151366 79898
rect 151314 79834 151366 79840
rect 151406 79892 151458 79898
rect 151406 79834 151458 79840
rect 151602 79812 151630 80036
rect 151694 79971 151722 80036
rect 151680 79962 151736 79971
rect 151680 79897 151736 79906
rect 151602 79784 151676 79812
rect 151786 79801 151814 80036
rect 151878 79966 151906 80036
rect 151970 79966 151998 80036
rect 151866 79960 151918 79966
rect 151866 79902 151918 79908
rect 151958 79960 152010 79966
rect 152062 79937 152090 80036
rect 151958 79902 152010 79908
rect 152048 79928 152104 79937
rect 152048 79863 152104 79872
rect 152154 79830 152182 80036
rect 152246 79898 152274 80036
rect 152234 79892 152286 79898
rect 152234 79834 152286 79840
rect 152142 79824 152194 79830
rect 151050 79716 151124 79744
rect 150532 79630 150584 79636
rect 150714 79656 150770 79665
rect 150440 78668 150492 78674
rect 150440 78610 150492 78616
rect 150348 78396 150400 78402
rect 150348 78338 150400 78344
rect 150254 78296 150310 78305
rect 150254 78231 150310 78240
rect 150544 77294 150572 79630
rect 150866 79648 150940 79676
rect 150714 79591 150770 79600
rect 150728 78520 150756 79591
rect 150808 79552 150860 79558
rect 150808 79494 150860 79500
rect 150636 78492 150756 78520
rect 150636 78130 150664 78492
rect 150716 78396 150768 78402
rect 150716 78338 150768 78344
rect 150624 78124 150676 78130
rect 150624 78066 150676 78072
rect 150544 77266 150664 77294
rect 150636 75750 150664 77266
rect 150624 75744 150676 75750
rect 150624 75686 150676 75692
rect 150164 75336 150216 75342
rect 150164 75278 150216 75284
rect 150728 73098 150756 78338
rect 150716 73092 150768 73098
rect 150716 73034 150768 73040
rect 150072 72616 150124 72622
rect 150072 72558 150124 72564
rect 150820 71534 150848 79494
rect 150912 72758 150940 79648
rect 150992 79620 151044 79626
rect 150992 79562 151044 79568
rect 151004 78878 151032 79562
rect 150992 78872 151044 78878
rect 150992 78814 151044 78820
rect 150992 78056 151044 78062
rect 150992 77998 151044 78004
rect 150900 72752 150952 72758
rect 150900 72694 150952 72700
rect 151004 71738 151032 77998
rect 151096 75682 151124 79716
rect 151452 79688 151504 79694
rect 151174 79656 151230 79665
rect 151452 79630 151504 79636
rect 151544 79688 151596 79694
rect 151544 79630 151596 79636
rect 151174 79591 151230 79600
rect 151268 79620 151320 79626
rect 151188 78062 151216 79591
rect 151268 79562 151320 79568
rect 151360 79620 151412 79626
rect 151360 79562 151412 79568
rect 151176 78056 151228 78062
rect 151176 77998 151228 78004
rect 151084 75676 151136 75682
rect 151084 75618 151136 75624
rect 151280 73166 151308 79562
rect 151372 75546 151400 79562
rect 151464 77790 151492 79630
rect 151452 77784 151504 77790
rect 151452 77726 151504 77732
rect 151360 75540 151412 75546
rect 151360 75482 151412 75488
rect 151556 74322 151584 79630
rect 151648 78169 151676 79784
rect 151772 79792 151828 79801
rect 152142 79766 152194 79772
rect 152338 79744 152366 80036
rect 152430 79937 152458 80036
rect 152522 79966 152550 80036
rect 152510 79960 152562 79966
rect 152416 79928 152472 79937
rect 152510 79902 152562 79908
rect 152614 79898 152642 80036
rect 152706 79966 152734 80036
rect 152798 79971 152826 80036
rect 152694 79960 152746 79966
rect 152694 79902 152746 79908
rect 152784 79962 152840 79971
rect 152416 79863 152472 79872
rect 152602 79892 152654 79898
rect 152784 79897 152840 79906
rect 152602 79834 152654 79840
rect 152890 79812 152918 80036
rect 152982 79966 153010 80036
rect 153074 79971 153102 80036
rect 152970 79960 153022 79966
rect 152970 79902 153022 79908
rect 153060 79962 153116 79971
rect 153166 79966 153194 80036
rect 153258 79966 153286 80036
rect 153350 79966 153378 80036
rect 153442 79966 153470 80036
rect 153060 79897 153116 79906
rect 153154 79960 153206 79966
rect 153154 79902 153206 79908
rect 153246 79960 153298 79966
rect 153246 79902 153298 79908
rect 153338 79960 153390 79966
rect 153338 79902 153390 79908
rect 153430 79960 153482 79966
rect 153430 79902 153482 79908
rect 152844 79784 152918 79812
rect 151772 79727 151828 79736
rect 152246 79716 152366 79744
rect 152556 79756 152608 79762
rect 151728 79688 151780 79694
rect 152004 79688 152056 79694
rect 151728 79630 151780 79636
rect 151818 79656 151874 79665
rect 151740 79014 151768 79630
rect 152004 79630 152056 79636
rect 152096 79688 152148 79694
rect 152246 79642 152274 79716
rect 152844 79744 152872 79784
rect 153534 79778 153562 80036
rect 152556 79698 152608 79704
rect 152798 79716 152872 79744
rect 153016 79756 153068 79762
rect 152568 79642 152596 79698
rect 152798 79676 152826 79716
rect 153016 79698 153068 79704
rect 153108 79756 153160 79762
rect 153108 79698 153160 79704
rect 153200 79756 153252 79762
rect 153200 79698 153252 79704
rect 153396 79750 153562 79778
rect 152096 79630 152148 79636
rect 151818 79591 151874 79600
rect 151912 79620 151964 79626
rect 151728 79008 151780 79014
rect 151728 78950 151780 78956
rect 151728 78872 151780 78878
rect 151728 78814 151780 78820
rect 151634 78160 151690 78169
rect 151634 78095 151690 78104
rect 151636 78056 151688 78062
rect 151636 77998 151688 78004
rect 151648 76430 151676 77998
rect 151636 76424 151688 76430
rect 151636 76366 151688 76372
rect 151740 75954 151768 78814
rect 151728 75948 151780 75954
rect 151728 75890 151780 75896
rect 151832 75018 151860 79591
rect 151912 79562 151964 79568
rect 151924 75206 151952 79562
rect 152016 75274 152044 79630
rect 152004 75268 152056 75274
rect 152004 75210 152056 75216
rect 151912 75200 151964 75206
rect 151912 75142 151964 75148
rect 151832 74990 152044 75018
rect 151912 74928 151964 74934
rect 151912 74870 151964 74876
rect 151820 74860 151872 74866
rect 151820 74802 151872 74808
rect 151544 74316 151596 74322
rect 151544 74258 151596 74264
rect 151268 73160 151320 73166
rect 151268 73102 151320 73108
rect 150992 71732 151044 71738
rect 150992 71674 151044 71680
rect 150808 71528 150860 71534
rect 150808 71470 150860 71476
rect 149704 61532 149756 61538
rect 149704 61474 149756 61480
rect 149612 60036 149664 60042
rect 149612 59978 149664 59984
rect 149520 27056 149572 27062
rect 149520 26998 149572 27004
rect 149428 14816 149480 14822
rect 149428 14758 149480 14764
rect 149336 10464 149388 10470
rect 149336 10406 149388 10412
rect 149244 10396 149296 10402
rect 149244 10338 149296 10344
rect 149164 6886 149560 6914
rect 148692 4956 148744 4962
rect 148692 4898 148744 4904
rect 149532 480 149560 6886
rect 151832 6322 151860 74802
rect 151924 12238 151952 74870
rect 152016 12306 152044 74990
rect 152108 16114 152136 79630
rect 152200 79614 152274 79642
rect 152476 79614 152596 79642
rect 152752 79648 152826 79676
rect 152200 21758 152228 79614
rect 152372 79076 152424 79082
rect 152372 79018 152424 79024
rect 152280 78736 152332 78742
rect 152280 78678 152332 78684
rect 152292 29714 152320 78678
rect 152384 78198 152412 79018
rect 152476 78742 152504 79614
rect 152556 79552 152608 79558
rect 152556 79494 152608 79500
rect 152464 78736 152516 78742
rect 152464 78678 152516 78684
rect 152372 78192 152424 78198
rect 152372 78134 152424 78140
rect 152372 77988 152424 77994
rect 152372 77930 152424 77936
rect 152384 77382 152412 77930
rect 152372 77376 152424 77382
rect 152372 77318 152424 77324
rect 152372 77240 152424 77246
rect 152372 77182 152424 77188
rect 152384 76906 152412 77182
rect 152372 76900 152424 76906
rect 152372 76842 152424 76848
rect 152464 75268 152516 75274
rect 152464 75210 152516 75216
rect 152372 75200 152424 75206
rect 152372 75142 152424 75148
rect 152384 29782 152412 75142
rect 152476 62966 152504 75210
rect 152568 64326 152596 79494
rect 152648 79416 152700 79422
rect 152648 79358 152700 79364
rect 152660 79150 152688 79358
rect 152648 79144 152700 79150
rect 152648 79086 152700 79092
rect 152648 79008 152700 79014
rect 152648 78950 152700 78956
rect 152660 77994 152688 78950
rect 152752 78441 152780 79648
rect 152832 79552 152884 79558
rect 152832 79494 152884 79500
rect 152924 79552 152976 79558
rect 152924 79494 152976 79500
rect 152738 78432 152794 78441
rect 152738 78367 152794 78376
rect 152648 77988 152700 77994
rect 152648 77930 152700 77936
rect 152844 77294 152872 79494
rect 152660 77266 152872 77294
rect 152936 77294 152964 79494
rect 153028 78305 153056 79698
rect 153120 78418 153148 79698
rect 153212 79082 153240 79698
rect 153292 79688 153344 79694
rect 153292 79630 153344 79636
rect 153200 79076 153252 79082
rect 153200 79018 153252 79024
rect 153198 78432 153254 78441
rect 153120 78390 153198 78418
rect 153198 78367 153254 78376
rect 153014 78296 153070 78305
rect 153014 78231 153070 78240
rect 153198 78160 153254 78169
rect 153198 78095 153254 78104
rect 152936 77266 153148 77294
rect 152660 74866 152688 77266
rect 153120 74934 153148 77266
rect 153108 74928 153160 74934
rect 153108 74870 153160 74876
rect 152648 74860 152700 74866
rect 152648 74802 152700 74808
rect 153212 72554 153240 78095
rect 153200 72548 153252 72554
rect 153200 72490 153252 72496
rect 152556 64320 152608 64326
rect 152556 64262 152608 64268
rect 152464 62960 152516 62966
rect 152464 62902 152516 62908
rect 152372 29776 152424 29782
rect 152372 29718 152424 29724
rect 152280 29708 152332 29714
rect 152280 29650 152332 29656
rect 152188 21752 152240 21758
rect 152188 21694 152240 21700
rect 152096 16108 152148 16114
rect 152096 16050 152148 16056
rect 153304 13190 153332 79630
rect 153396 79608 153424 79750
rect 153626 79744 153654 80036
rect 153718 79971 153746 80036
rect 153704 79962 153760 79971
rect 153704 79897 153760 79906
rect 153810 79744 153838 80036
rect 153902 79971 153930 80036
rect 153888 79962 153944 79971
rect 153888 79897 153944 79906
rect 153626 79716 153700 79744
rect 153396 79580 153470 79608
rect 153442 79506 153470 79580
rect 153396 79478 153470 79506
rect 153568 79552 153620 79558
rect 153568 79494 153620 79500
rect 153396 79014 153424 79478
rect 153476 79416 153528 79422
rect 153476 79358 153528 79364
rect 153384 79008 153436 79014
rect 153384 78950 153436 78956
rect 153384 78124 153436 78130
rect 153384 78066 153436 78072
rect 153292 13184 153344 13190
rect 153292 13126 153344 13132
rect 153396 13122 153424 78066
rect 153488 16046 153516 79358
rect 153580 35222 153608 79494
rect 153672 79422 153700 79716
rect 153764 79716 153838 79744
rect 153994 79744 154022 80036
rect 154086 79966 154114 80036
rect 154074 79960 154126 79966
rect 154178 79937 154206 80036
rect 154074 79902 154126 79908
rect 154164 79928 154220 79937
rect 154164 79863 154220 79872
rect 154270 79778 154298 80036
rect 154362 79937 154390 80036
rect 154348 79928 154404 79937
rect 154348 79863 154404 79872
rect 154454 79830 154482 80036
rect 154442 79824 154494 79830
rect 154120 79756 154172 79762
rect 153994 79716 154068 79744
rect 153660 79416 153712 79422
rect 153660 79358 153712 79364
rect 153764 78656 153792 79716
rect 153934 79656 153990 79665
rect 153934 79591 153990 79600
rect 153844 79008 153896 79014
rect 153844 78950 153896 78956
rect 153672 78628 153792 78656
rect 153672 61470 153700 78628
rect 153856 78588 153884 78950
rect 153764 78560 153884 78588
rect 153764 68542 153792 78560
rect 153844 77784 153896 77790
rect 153844 77726 153896 77732
rect 153856 70394 153884 77726
rect 153948 77194 153976 79591
rect 154040 77897 154068 79716
rect 154270 79750 154344 79778
rect 154442 79766 154494 79772
rect 154120 79698 154172 79704
rect 154132 78130 154160 79698
rect 154212 79688 154264 79694
rect 154210 79656 154212 79665
rect 154264 79656 154266 79665
rect 154210 79591 154266 79600
rect 154212 79552 154264 79558
rect 154212 79494 154264 79500
rect 154224 79150 154252 79494
rect 154212 79144 154264 79150
rect 154212 79086 154264 79092
rect 154316 78792 154344 79750
rect 154546 79676 154574 80036
rect 154638 79966 154666 80036
rect 154626 79960 154678 79966
rect 154626 79902 154678 79908
rect 154730 79744 154758 80036
rect 154822 79971 154850 80036
rect 154808 79962 154864 79971
rect 154808 79897 154864 79906
rect 154914 79898 154942 80036
rect 155006 79971 155034 80036
rect 154992 79962 155048 79971
rect 154902 79892 154954 79898
rect 154992 79897 155048 79906
rect 154902 79834 154954 79840
rect 155098 79830 155126 80036
rect 155086 79824 155138 79830
rect 154684 79716 154758 79744
rect 154946 79792 155002 79801
rect 155086 79766 155138 79772
rect 154946 79727 155002 79736
rect 154546 79648 154620 79676
rect 154316 78764 154528 78792
rect 154304 78668 154356 78674
rect 154304 78610 154356 78616
rect 154120 78124 154172 78130
rect 154120 78066 154172 78072
rect 154118 78024 154174 78033
rect 154118 77959 154174 77968
rect 154132 77926 154160 77959
rect 154120 77920 154172 77926
rect 154026 77888 154082 77897
rect 154120 77862 154172 77868
rect 154026 77823 154082 77832
rect 153948 77166 154252 77194
rect 154224 70394 154252 77166
rect 154316 74118 154344 78610
rect 154394 78296 154450 78305
rect 154394 78231 154450 78240
rect 154408 75914 154436 78231
rect 154500 78062 154528 78764
rect 154592 78169 154620 79648
rect 154578 78160 154634 78169
rect 154578 78095 154634 78104
rect 154488 78056 154540 78062
rect 154488 77998 154540 78004
rect 154684 77858 154712 79716
rect 154762 79656 154818 79665
rect 154762 79591 154818 79600
rect 154856 79620 154908 79626
rect 154672 77852 154724 77858
rect 154672 77794 154724 77800
rect 154408 75886 154620 75914
rect 154592 75614 154620 75886
rect 154580 75608 154632 75614
rect 154580 75550 154632 75556
rect 154670 75576 154726 75585
rect 154670 75511 154726 75520
rect 154304 74112 154356 74118
rect 154304 74054 154356 74060
rect 154684 71602 154712 75511
rect 154672 71596 154724 71602
rect 154672 71538 154724 71544
rect 154776 71262 154804 79591
rect 154856 79562 154908 79568
rect 154868 79014 154896 79562
rect 154856 79008 154908 79014
rect 154856 78950 154908 78956
rect 154856 75948 154908 75954
rect 154856 75890 154908 75896
rect 154868 71466 154896 75890
rect 154856 71460 154908 71466
rect 154856 71402 154908 71408
rect 154764 71256 154816 71262
rect 154764 71198 154816 71204
rect 154960 70394 154988 79727
rect 155040 79688 155092 79694
rect 155190 79676 155218 80036
rect 155282 79830 155310 80036
rect 155374 79830 155402 80036
rect 155466 79830 155494 80036
rect 155270 79824 155322 79830
rect 155270 79766 155322 79772
rect 155362 79824 155414 79830
rect 155362 79766 155414 79772
rect 155454 79824 155506 79830
rect 155454 79766 155506 79772
rect 155558 79744 155586 80036
rect 155650 79971 155678 80036
rect 155636 79962 155692 79971
rect 155636 79897 155692 79906
rect 155742 79812 155770 80036
rect 155834 79898 155862 80036
rect 155822 79892 155874 79898
rect 155822 79834 155874 79840
rect 155696 79801 155770 79812
rect 155682 79792 155770 79801
rect 155558 79716 155632 79744
rect 155738 79784 155770 79792
rect 155926 79812 155954 80036
rect 156018 79966 156046 80036
rect 156006 79960 156058 79966
rect 156110 79937 156138 80036
rect 156202 79966 156230 80036
rect 156190 79960 156242 79966
rect 156006 79902 156058 79908
rect 156096 79928 156152 79937
rect 156190 79902 156242 79908
rect 156096 79863 156152 79872
rect 156052 79824 156104 79830
rect 155926 79784 156000 79812
rect 155682 79727 155738 79736
rect 155040 79630 155092 79636
rect 155144 79648 155218 79676
rect 155408 79688 155460 79694
rect 155052 76770 155080 79630
rect 155144 79506 155172 79648
rect 155408 79630 155460 79636
rect 155316 79620 155368 79626
rect 155316 79562 155368 79568
rect 155144 79478 155264 79506
rect 155132 79416 155184 79422
rect 155132 79358 155184 79364
rect 155144 79150 155172 79358
rect 155132 79144 155184 79150
rect 155132 79086 155184 79092
rect 155040 76764 155092 76770
rect 155040 76706 155092 76712
rect 155236 76498 155264 79478
rect 155224 76492 155276 76498
rect 155224 76434 155276 76440
rect 155328 75914 155356 79562
rect 155420 78266 155448 79630
rect 155500 79620 155552 79626
rect 155500 79562 155552 79568
rect 155408 78260 155460 78266
rect 155408 78202 155460 78208
rect 155512 78130 155540 79562
rect 155500 78124 155552 78130
rect 155500 78066 155552 78072
rect 155500 77920 155552 77926
rect 155500 77862 155552 77868
rect 155328 75886 155448 75914
rect 155316 73160 155368 73166
rect 155316 73102 155368 73108
rect 153856 70366 154160 70394
rect 154224 70366 154436 70394
rect 153752 68536 153804 68542
rect 153752 68478 153804 68484
rect 153660 61464 153712 61470
rect 153660 61406 153712 61412
rect 153568 35216 153620 35222
rect 153568 35158 153620 35164
rect 154132 29850 154160 70366
rect 154120 29844 154172 29850
rect 154120 29786 154172 29792
rect 153476 16040 153528 16046
rect 153476 15982 153528 15988
rect 153384 13116 153436 13122
rect 153384 13058 153436 13064
rect 152004 12300 152056 12306
rect 152004 12242 152056 12248
rect 151912 12232 151964 12238
rect 151912 12174 151964 12180
rect 151820 6316 151872 6322
rect 151820 6258 151872 6264
rect 154212 5296 154264 5302
rect 154212 5238 154264 5244
rect 153016 4140 153068 4146
rect 153016 4082 153068 4088
rect 151820 3596 151872 3602
rect 151820 3538 151872 3544
rect 150624 3324 150676 3330
rect 150624 3266 150676 3272
rect 150636 480 150664 3266
rect 151832 480 151860 3538
rect 153028 480 153056 4082
rect 154224 480 154252 5238
rect 154408 5098 154436 70366
rect 154684 70366 154988 70394
rect 155328 70378 155356 73102
rect 155420 71330 155448 75886
rect 155512 71398 155540 77862
rect 155604 75914 155632 79716
rect 155868 79688 155920 79694
rect 155868 79630 155920 79636
rect 155684 79552 155736 79558
rect 155684 79494 155736 79500
rect 155696 76362 155724 79494
rect 155880 78538 155908 79630
rect 155868 78532 155920 78538
rect 155868 78474 155920 78480
rect 155868 78124 155920 78130
rect 155868 78066 155920 78072
rect 155684 76356 155736 76362
rect 155684 76298 155736 76304
rect 155604 75886 155724 75914
rect 155696 75410 155724 75886
rect 155684 75404 155736 75410
rect 155684 75346 155736 75352
rect 155776 73092 155828 73098
rect 155776 73034 155828 73040
rect 155500 71392 155552 71398
rect 155500 71334 155552 71340
rect 155408 71324 155460 71330
rect 155408 71266 155460 71272
rect 155316 70372 155368 70378
rect 154684 70106 154712 70366
rect 155316 70314 155368 70320
rect 155788 70310 155816 73034
rect 155776 70304 155828 70310
rect 155776 70246 155828 70252
rect 154672 70100 154724 70106
rect 154672 70042 154724 70048
rect 155880 70038 155908 78066
rect 155972 77722 156000 79784
rect 156052 79766 156104 79772
rect 155960 77716 156012 77722
rect 155960 77658 156012 77664
rect 156064 76974 156092 79766
rect 156144 79756 156196 79762
rect 156144 79698 156196 79704
rect 156156 78130 156184 79698
rect 156294 79676 156322 80036
rect 156386 79830 156414 80036
rect 156478 79971 156506 80036
rect 156464 79962 156520 79971
rect 156464 79897 156520 79906
rect 156374 79824 156426 79830
rect 156374 79766 156426 79772
rect 156570 79744 156598 80036
rect 156662 79937 156690 80036
rect 156754 79966 156782 80036
rect 156846 79966 156874 80036
rect 156742 79960 156794 79966
rect 156648 79928 156704 79937
rect 156742 79902 156794 79908
rect 156834 79960 156886 79966
rect 156938 79937 156966 80036
rect 156834 79902 156886 79908
rect 156924 79928 156980 79937
rect 156648 79863 156704 79872
rect 156924 79863 156980 79872
rect 157030 79812 157058 80036
rect 157122 79971 157150 80036
rect 157108 79962 157164 79971
rect 157214 79966 157242 80036
rect 157306 79966 157334 80036
rect 157398 79966 157426 80036
rect 157108 79897 157164 79906
rect 157202 79960 157254 79966
rect 157202 79902 157254 79908
rect 157294 79960 157346 79966
rect 157294 79902 157346 79908
rect 157386 79960 157438 79966
rect 157386 79902 157438 79908
rect 157490 79898 157518 80036
rect 157478 79892 157530 79898
rect 157478 79834 157530 79840
rect 157582 79830 157610 80036
rect 157156 79824 157208 79830
rect 157030 79784 157104 79812
rect 156880 79756 156932 79762
rect 156570 79716 156644 79744
rect 156248 79648 156322 79676
rect 156144 78124 156196 78130
rect 156144 78066 156196 78072
rect 156142 78024 156198 78033
rect 156142 77959 156198 77968
rect 156052 76968 156104 76974
rect 156052 76910 156104 76916
rect 156156 75478 156184 77959
rect 156144 75472 156196 75478
rect 156144 75414 156196 75420
rect 156248 74390 156276 79648
rect 156328 79552 156380 79558
rect 156328 79494 156380 79500
rect 156236 74384 156288 74390
rect 156236 74326 156288 74332
rect 156340 70394 156368 79494
rect 156420 78124 156472 78130
rect 156420 78066 156472 78072
rect 156432 73914 156460 78066
rect 156616 74254 156644 79716
rect 156880 79698 156932 79704
rect 156788 79688 156840 79694
rect 156786 79656 156788 79665
rect 156840 79656 156842 79665
rect 156696 79620 156748 79626
rect 156892 79642 156920 79698
rect 156892 79614 157012 79642
rect 156786 79591 156842 79600
rect 156696 79562 156748 79568
rect 156708 78713 156736 79562
rect 156788 79552 156840 79558
rect 156788 79494 156840 79500
rect 156694 78704 156750 78713
rect 156694 78639 156750 78648
rect 156696 78532 156748 78538
rect 156696 78474 156748 78480
rect 156708 75138 156736 78474
rect 156800 75818 156828 79494
rect 156788 75812 156840 75818
rect 156788 75754 156840 75760
rect 156696 75132 156748 75138
rect 156696 75074 156748 75080
rect 156604 74248 156656 74254
rect 156604 74190 156656 74196
rect 156878 74080 156934 74089
rect 156878 74015 156934 74024
rect 156420 73908 156472 73914
rect 156420 73850 156472 73856
rect 155972 70366 156368 70394
rect 155972 70174 156000 70366
rect 155960 70168 156012 70174
rect 155960 70110 156012 70116
rect 155868 70032 155920 70038
rect 155868 69974 155920 69980
rect 156892 69970 156920 74015
rect 156984 73982 157012 79614
rect 157076 77625 157104 79784
rect 157570 79824 157622 79830
rect 157156 79766 157208 79772
rect 157430 79792 157486 79801
rect 157168 78713 157196 79766
rect 157570 79766 157622 79772
rect 157430 79727 157486 79736
rect 157674 79744 157702 80036
rect 157766 79937 157794 80036
rect 157752 79928 157808 79937
rect 157752 79863 157808 79872
rect 157858 79812 157886 80036
rect 157812 79801 157886 79812
rect 157950 79801 157978 80036
rect 158042 79966 158070 80036
rect 158134 79966 158162 80036
rect 158030 79960 158082 79966
rect 158030 79902 158082 79908
rect 158122 79960 158174 79966
rect 158226 79937 158254 80036
rect 158122 79902 158174 79908
rect 158212 79928 158268 79937
rect 158212 79863 158268 79872
rect 157798 79792 157886 79801
rect 157248 79688 157300 79694
rect 157248 79630 157300 79636
rect 157154 78704 157210 78713
rect 157154 78639 157210 78648
rect 157062 77616 157118 77625
rect 157062 77551 157118 77560
rect 157260 74050 157288 79630
rect 157444 79286 157472 79727
rect 157674 79716 157748 79744
rect 157854 79784 157886 79792
rect 157936 79792 157992 79801
rect 157798 79727 157854 79736
rect 158318 79778 158346 80036
rect 157936 79727 157992 79736
rect 158076 79756 158128 79762
rect 157524 79688 157576 79694
rect 157524 79630 157576 79636
rect 157340 79280 157392 79286
rect 157340 79222 157392 79228
rect 157432 79280 157484 79286
rect 157432 79222 157484 79228
rect 157352 78878 157380 79222
rect 157432 78940 157484 78946
rect 157432 78882 157484 78888
rect 157340 78872 157392 78878
rect 157340 78814 157392 78820
rect 157444 78538 157472 78882
rect 157432 78532 157484 78538
rect 157432 78474 157484 78480
rect 157430 78432 157486 78441
rect 157430 78367 157486 78376
rect 157338 78296 157394 78305
rect 157338 78231 157394 78240
rect 157248 74044 157300 74050
rect 157248 73986 157300 73992
rect 156972 73976 157024 73982
rect 156972 73918 157024 73924
rect 156880 69964 156932 69970
rect 156880 69906 156932 69912
rect 157352 15910 157380 78231
rect 157444 76906 157472 78367
rect 157432 76900 157484 76906
rect 157432 76842 157484 76848
rect 157432 75336 157484 75342
rect 157432 75278 157484 75284
rect 157444 15978 157472 75278
rect 157536 75274 157564 79630
rect 157616 79620 157668 79626
rect 157616 79562 157668 79568
rect 157628 77926 157656 79562
rect 157720 78690 157748 79716
rect 158076 79698 158128 79704
rect 158180 79750 158346 79778
rect 157984 79620 158036 79626
rect 157984 79562 158036 79568
rect 157800 79552 157852 79558
rect 157800 79494 157852 79500
rect 157812 78946 157840 79494
rect 157996 79286 158024 79562
rect 157892 79280 157944 79286
rect 157892 79222 157944 79228
rect 157984 79280 158036 79286
rect 157984 79222 158036 79228
rect 157800 78940 157852 78946
rect 157800 78882 157852 78888
rect 157904 78792 157932 79222
rect 157904 78764 158024 78792
rect 157720 78662 157932 78690
rect 157706 78432 157762 78441
rect 157706 78367 157762 78376
rect 157616 77920 157668 77926
rect 157616 77862 157668 77868
rect 157524 75268 157576 75274
rect 157524 75210 157576 75216
rect 157616 75200 157668 75206
rect 157616 75142 157668 75148
rect 157524 75132 157576 75138
rect 157524 75074 157576 75080
rect 157536 20126 157564 75074
rect 157628 24614 157656 75142
rect 157720 25634 157748 78367
rect 157800 75268 157852 75274
rect 157800 75210 157852 75216
rect 157812 29646 157840 75210
rect 157904 61402 157932 78662
rect 157996 75138 158024 78764
rect 158088 75206 158116 79698
rect 158180 79422 158208 79750
rect 158410 79744 158438 80036
rect 158502 79903 158530 80036
rect 158488 79894 158544 79903
rect 158594 79898 158622 80036
rect 158488 79829 158544 79838
rect 158582 79892 158634 79898
rect 158582 79834 158634 79840
rect 158686 79744 158714 80036
rect 158778 79898 158806 80036
rect 158870 79966 158898 80036
rect 158858 79960 158910 79966
rect 158962 79937 158990 80036
rect 159054 79966 159082 80036
rect 159042 79960 159094 79966
rect 158858 79902 158910 79908
rect 158948 79928 159004 79937
rect 158766 79892 158818 79898
rect 159042 79902 159094 79908
rect 158948 79863 159004 79872
rect 158766 79834 158818 79840
rect 158904 79824 158956 79830
rect 158904 79766 158956 79772
rect 158410 79716 158484 79744
rect 158686 79716 158760 79744
rect 158260 79620 158312 79626
rect 158260 79562 158312 79568
rect 158168 79416 158220 79422
rect 158168 79358 158220 79364
rect 158166 78432 158222 78441
rect 158166 78367 158222 78376
rect 158180 75342 158208 78367
rect 158272 78198 158300 79562
rect 158352 79416 158404 79422
rect 158352 79358 158404 79364
rect 158260 78192 158312 78198
rect 158260 78134 158312 78140
rect 158260 77852 158312 77858
rect 158260 77794 158312 77800
rect 158168 75336 158220 75342
rect 158168 75278 158220 75284
rect 158076 75200 158128 75206
rect 158076 75142 158128 75148
rect 157984 75132 158036 75138
rect 157984 75074 158036 75080
rect 158272 70394 158300 77794
rect 158364 77081 158392 79358
rect 158456 78033 158484 79716
rect 158536 79688 158588 79694
rect 158536 79630 158588 79636
rect 158442 78024 158498 78033
rect 158442 77959 158498 77968
rect 158350 77072 158406 77081
rect 158350 77007 158406 77016
rect 158352 76900 158404 76906
rect 158352 76842 158404 76848
rect 158364 72486 158392 76842
rect 158548 75914 158576 79630
rect 158628 79620 158680 79626
rect 158628 79562 158680 79568
rect 158640 78810 158668 79562
rect 158628 78804 158680 78810
rect 158628 78746 158680 78752
rect 158732 78198 158760 79716
rect 158810 78296 158866 78305
rect 158810 78231 158866 78240
rect 158720 78192 158772 78198
rect 158720 78134 158772 78140
rect 158628 78056 158680 78062
rect 158628 77998 158680 78004
rect 158456 75886 158576 75914
rect 158456 75313 158484 75886
rect 158442 75304 158498 75313
rect 158442 75239 158498 75248
rect 158640 73846 158668 77998
rect 158628 73840 158680 73846
rect 158628 73782 158680 73788
rect 158352 72480 158404 72486
rect 158352 72422 158404 72428
rect 158180 70366 158300 70394
rect 158180 64874 158208 70366
rect 157996 64846 158208 64874
rect 157996 64258 158024 64846
rect 157984 64252 158036 64258
rect 157984 64194 158036 64200
rect 157892 61396 157944 61402
rect 157892 61338 157944 61344
rect 157800 29640 157852 29646
rect 157800 29582 157852 29588
rect 157708 25628 157760 25634
rect 157708 25570 157760 25576
rect 157616 24608 157668 24614
rect 157616 24550 157668 24556
rect 157524 20120 157576 20126
rect 157524 20062 157576 20068
rect 157432 15972 157484 15978
rect 157432 15914 157484 15920
rect 157340 15904 157392 15910
rect 157340 15846 157392 15852
rect 158824 11966 158852 78231
rect 158916 75274 158944 79766
rect 159146 79744 159174 80036
rect 159238 79898 159266 80036
rect 159330 79966 159358 80036
rect 159318 79960 159370 79966
rect 159318 79902 159370 79908
rect 159226 79892 159278 79898
rect 159226 79834 159278 79840
rect 159422 79835 159450 80036
rect 159514 79898 159542 80036
rect 159606 79898 159634 80036
rect 159502 79892 159554 79898
rect 159408 79826 159464 79835
rect 159502 79834 159554 79840
rect 159594 79892 159646 79898
rect 159594 79834 159646 79840
rect 159008 79716 159174 79744
rect 159270 79792 159326 79801
rect 159408 79761 159464 79770
rect 159698 79744 159726 80036
rect 159790 79937 159818 80036
rect 159776 79928 159832 79937
rect 159776 79863 159832 79872
rect 159882 79801 159910 80036
rect 159974 79937 160002 80036
rect 160066 79966 160094 80036
rect 160158 79966 160186 80036
rect 160054 79960 160106 79966
rect 159960 79928 160016 79937
rect 160054 79902 160106 79908
rect 160146 79960 160198 79966
rect 160146 79902 160198 79908
rect 159960 79863 160016 79872
rect 160146 79824 160198 79830
rect 159270 79727 159326 79736
rect 158904 75268 158956 75274
rect 158904 75210 158956 75216
rect 159008 70394 159036 79716
rect 159180 78940 159232 78946
rect 159180 78882 159232 78888
rect 159088 78804 159140 78810
rect 159088 78746 159140 78752
rect 159100 77294 159128 78746
rect 159192 78062 159220 78882
rect 159180 78056 159232 78062
rect 159180 77998 159232 78004
rect 159180 77784 159232 77790
rect 159180 77726 159232 77732
rect 159192 77518 159220 77726
rect 159180 77512 159232 77518
rect 159180 77454 159232 77460
rect 159100 77266 159220 77294
rect 159088 75268 159140 75274
rect 159088 75210 159140 75216
rect 158916 70366 159036 70394
rect 158916 12034 158944 70366
rect 159100 12102 159128 75210
rect 159192 14550 159220 77266
rect 159284 14686 159312 79727
rect 159652 79716 159726 79744
rect 159868 79792 159924 79801
rect 160146 79766 160198 79772
rect 159868 79727 159924 79736
rect 159456 79688 159508 79694
rect 159376 79648 159456 79676
rect 159272 14680 159324 14686
rect 159272 14622 159324 14628
rect 159376 14618 159404 79648
rect 159456 79630 159508 79636
rect 159456 79552 159508 79558
rect 159456 79494 159508 79500
rect 159468 76702 159496 79494
rect 159652 78810 159680 79716
rect 159916 79688 159968 79694
rect 160158 79676 160186 79766
rect 160250 79744 160278 80036
rect 160342 79898 160370 80036
rect 160434 79966 160462 80036
rect 160422 79960 160474 79966
rect 160422 79902 160474 79908
rect 160330 79892 160382 79898
rect 160330 79834 160382 79840
rect 160526 79812 160554 80036
rect 160618 79966 160646 80036
rect 160710 79971 160738 80036
rect 160606 79960 160658 79966
rect 160606 79902 160658 79908
rect 160696 79962 160752 79971
rect 160802 79966 160830 80036
rect 160894 79966 160922 80036
rect 160696 79897 160752 79906
rect 160790 79960 160842 79966
rect 160790 79902 160842 79908
rect 160882 79960 160934 79966
rect 160882 79902 160934 79908
rect 160882 79824 160934 79830
rect 160526 79784 160600 79812
rect 160250 79716 160324 79744
rect 159916 79630 159968 79636
rect 160006 79656 160062 79665
rect 159732 79416 159784 79422
rect 159732 79358 159784 79364
rect 159640 78804 159692 78810
rect 159640 78746 159692 78752
rect 159640 78260 159692 78266
rect 159640 78202 159692 78208
rect 159456 76696 159508 76702
rect 159456 76638 159508 76644
rect 159652 14754 159680 78202
rect 159744 78033 159772 79358
rect 159730 78024 159786 78033
rect 159730 77959 159786 77968
rect 159928 70394 159956 79630
rect 160158 79648 160232 79676
rect 160006 79591 160062 79600
rect 160020 79558 160048 79591
rect 160008 79552 160060 79558
rect 160008 79494 160060 79500
rect 160008 79416 160060 79422
rect 160008 79358 160060 79364
rect 160020 75274 160048 79358
rect 160100 79076 160152 79082
rect 160100 79018 160152 79024
rect 160112 78810 160140 79018
rect 160100 78804 160152 78810
rect 160100 78746 160152 78752
rect 160100 78464 160152 78470
rect 160100 78406 160152 78412
rect 160112 78130 160140 78406
rect 160100 78124 160152 78130
rect 160100 78066 160152 78072
rect 160008 75268 160060 75274
rect 160008 75210 160060 75216
rect 160006 75168 160062 75177
rect 160006 75103 160062 75112
rect 159836 70366 159956 70394
rect 159640 14748 159692 14754
rect 159640 14690 159692 14696
rect 159364 14612 159416 14618
rect 159364 14554 159416 14560
rect 159180 14544 159232 14550
rect 159180 14486 159232 14492
rect 159088 12096 159140 12102
rect 159088 12038 159140 12044
rect 158904 12028 158956 12034
rect 158904 11970 158956 11976
rect 158812 11960 158864 11966
rect 158812 11902 158864 11908
rect 157800 5228 157852 5234
rect 157800 5170 157852 5176
rect 154396 5092 154448 5098
rect 154396 5034 154448 5040
rect 154486 4992 154542 5001
rect 154486 4927 154542 4936
rect 154500 3330 154528 4927
rect 156604 3936 156656 3942
rect 156604 3878 156656 3884
rect 155408 3732 155460 3738
rect 155408 3674 155460 3680
rect 154488 3324 154540 3330
rect 154488 3266 154540 3272
rect 155420 480 155448 3674
rect 156616 480 156644 3878
rect 157812 480 157840 5170
rect 158902 4856 158958 4865
rect 158902 4791 158958 4800
rect 158916 480 158944 4791
rect 159836 3738 159864 70366
rect 160020 11898 160048 75103
rect 160098 19952 160154 19961
rect 160098 19887 160154 19896
rect 160008 11892 160060 11898
rect 160008 11834 160060 11840
rect 159824 3732 159876 3738
rect 159824 3674 159876 3680
rect 160112 480 160140 19887
rect 160204 9586 160232 79648
rect 160192 9580 160244 9586
rect 160192 9522 160244 9528
rect 160296 9450 160324 79716
rect 160468 79688 160520 79694
rect 160468 79630 160520 79636
rect 160376 78464 160428 78470
rect 160376 78406 160428 78412
rect 160284 9444 160336 9450
rect 160284 9386 160336 9392
rect 160388 9178 160416 78406
rect 160480 9382 160508 79630
rect 160572 79422 160600 79784
rect 160880 79792 160882 79801
rect 160934 79792 160936 79801
rect 160880 79727 160936 79736
rect 160986 79744 161014 80036
rect 161078 79971 161106 80036
rect 161064 79962 161120 79971
rect 161064 79897 161120 79906
rect 161170 79898 161198 80036
rect 161262 79898 161290 80036
rect 161354 79898 161382 80036
rect 161446 79971 161474 80036
rect 161432 79962 161488 79971
rect 161538 79966 161566 80036
rect 161630 79971 161658 80036
rect 161158 79892 161210 79898
rect 161158 79834 161210 79840
rect 161250 79892 161302 79898
rect 161250 79834 161302 79840
rect 161342 79892 161394 79898
rect 161432 79897 161488 79906
rect 161526 79960 161578 79966
rect 161526 79902 161578 79908
rect 161616 79962 161672 79971
rect 161616 79897 161672 79906
rect 161722 79898 161750 80036
rect 161814 79937 161842 80036
rect 161906 79966 161934 80036
rect 161894 79960 161946 79966
rect 161800 79928 161856 79937
rect 161342 79834 161394 79840
rect 161710 79892 161762 79898
rect 161894 79902 161946 79908
rect 161998 79898 162026 80036
rect 161800 79863 161856 79872
rect 161986 79892 162038 79898
rect 161710 79834 161762 79840
rect 161986 79834 162038 79840
rect 161526 79824 161578 79830
rect 162090 79778 162118 80036
rect 162182 79971 162210 80036
rect 162168 79962 162224 79971
rect 162168 79897 162224 79906
rect 162274 79778 162302 80036
rect 162366 79898 162394 80036
rect 162458 79966 162486 80036
rect 162550 79971 162578 80036
rect 162446 79960 162498 79966
rect 162446 79902 162498 79908
rect 162536 79962 162592 79971
rect 162354 79892 162406 79898
rect 162536 79897 162592 79906
rect 162354 79834 162406 79840
rect 161578 79772 161704 79778
rect 161526 79766 161704 79772
rect 161112 79756 161164 79762
rect 160986 79716 161060 79744
rect 160744 79688 160796 79694
rect 160650 79656 160706 79665
rect 160744 79630 160796 79636
rect 160650 79591 160706 79600
rect 160560 79416 160612 79422
rect 160560 79358 160612 79364
rect 160664 79098 160692 79591
rect 160572 79070 160692 79098
rect 160468 9376 160520 9382
rect 160468 9318 160520 9324
rect 160572 9246 160600 79070
rect 160652 79008 160704 79014
rect 160652 78950 160704 78956
rect 160560 9240 160612 9246
rect 160560 9182 160612 9188
rect 160376 9172 160428 9178
rect 160376 9114 160428 9120
rect 160664 9110 160692 78950
rect 160756 78470 160784 79630
rect 160928 79552 160980 79558
rect 160928 79494 160980 79500
rect 160836 79484 160888 79490
rect 160836 79426 160888 79432
rect 160848 78878 160876 79426
rect 160836 78872 160888 78878
rect 160836 78814 160888 78820
rect 160744 78464 160796 78470
rect 160744 78406 160796 78412
rect 160742 78160 160798 78169
rect 160742 78095 160798 78104
rect 160756 21690 160784 78095
rect 160940 77654 160968 79494
rect 161032 79014 161060 79716
rect 161538 79750 161704 79766
rect 161112 79698 161164 79704
rect 161020 79008 161072 79014
rect 161020 78950 161072 78956
rect 161020 78872 161072 78878
rect 161020 78814 161072 78820
rect 161032 78538 161060 78814
rect 161020 78532 161072 78538
rect 161020 78474 161072 78480
rect 160928 77648 160980 77654
rect 160928 77590 160980 77596
rect 161124 75313 161152 79698
rect 161204 79688 161256 79694
rect 161204 79630 161256 79636
rect 161572 79688 161624 79694
rect 161572 79630 161624 79636
rect 161216 77489 161244 79630
rect 161584 79422 161612 79630
rect 161388 79416 161440 79422
rect 161388 79358 161440 79364
rect 161572 79416 161624 79422
rect 161572 79358 161624 79364
rect 161296 78124 161348 78130
rect 161296 78066 161348 78072
rect 161202 77480 161258 77489
rect 161202 77415 161258 77424
rect 161308 77194 161336 78066
rect 161216 77166 161336 77194
rect 161110 75304 161166 75313
rect 160836 75268 160888 75274
rect 161110 75239 161166 75248
rect 160836 75210 160888 75216
rect 160848 32638 160876 75210
rect 161216 70394 161244 77166
rect 161400 70394 161428 79358
rect 161572 79212 161624 79218
rect 161572 79154 161624 79160
rect 161480 79076 161532 79082
rect 161480 79018 161532 79024
rect 161492 78985 161520 79018
rect 161478 78976 161534 78985
rect 161478 78911 161534 78920
rect 161584 78713 161612 79154
rect 161570 78704 161626 78713
rect 161570 78639 161626 78648
rect 161572 77988 161624 77994
rect 161572 77930 161624 77936
rect 161124 70366 161244 70394
rect 161308 70366 161428 70394
rect 161124 64874 161152 70366
rect 161308 64874 161336 70366
rect 160940 64846 161152 64874
rect 161216 64846 161336 64874
rect 160836 32632 160888 32638
rect 160836 32574 160888 32580
rect 160744 21684 160796 21690
rect 160744 21626 160796 21632
rect 160652 9104 160704 9110
rect 160652 9046 160704 9052
rect 160940 6730 160968 64846
rect 161216 9314 161244 64846
rect 161204 9308 161256 9314
rect 161204 9250 161256 9256
rect 160928 6724 160980 6730
rect 160928 6666 160980 6672
rect 161584 3913 161612 77930
rect 161570 3904 161626 3913
rect 161570 3839 161626 3848
rect 161676 3602 161704 79750
rect 161940 79756 161992 79762
rect 162090 79750 162210 79778
rect 162274 79762 162348 79778
rect 162274 79756 162360 79762
rect 162274 79750 162308 79756
rect 161940 79698 161992 79704
rect 161846 79656 161902 79665
rect 161756 79620 161808 79626
rect 161846 79591 161902 79600
rect 161756 79562 161808 79568
rect 161768 78266 161796 79562
rect 161756 78260 161808 78266
rect 161756 78202 161808 78208
rect 161754 75304 161810 75313
rect 161754 75239 161810 75248
rect 161768 6254 161796 75239
rect 161860 9042 161888 79591
rect 161848 9036 161900 9042
rect 161848 8978 161900 8984
rect 161952 8974 161980 79698
rect 162032 79688 162084 79694
rect 162182 79642 162210 79750
rect 162642 79744 162670 80036
rect 162734 79971 162762 80036
rect 162720 79962 162776 79971
rect 162720 79897 162776 79906
rect 162826 79778 162854 80036
rect 162308 79698 162360 79704
rect 162596 79716 162670 79744
rect 162780 79750 162854 79778
rect 162400 79688 162452 79694
rect 162032 79630 162084 79636
rect 162044 11830 162072 79630
rect 162136 79614 162210 79642
rect 162306 79656 162362 79665
rect 162400 79630 162452 79636
rect 162492 79688 162544 79694
rect 162596 79665 162624 79716
rect 162492 79630 162544 79636
rect 162582 79656 162638 79665
rect 162136 77994 162164 79614
rect 162306 79591 162308 79600
rect 162360 79591 162362 79600
rect 162308 79562 162360 79568
rect 162308 79416 162360 79422
rect 162308 79358 162360 79364
rect 162216 79008 162268 79014
rect 162216 78950 162268 78956
rect 162228 78606 162256 78950
rect 162216 78600 162268 78606
rect 162216 78542 162268 78548
rect 162320 78470 162348 79358
rect 162308 78464 162360 78470
rect 162308 78406 162360 78412
rect 162308 78192 162360 78198
rect 162308 78134 162360 78140
rect 162124 77988 162176 77994
rect 162124 77930 162176 77936
rect 162216 77920 162268 77926
rect 162216 77862 162268 77868
rect 162124 77716 162176 77722
rect 162124 77658 162176 77664
rect 162136 70394 162164 77658
rect 162228 75018 162256 77862
rect 162320 77722 162348 78134
rect 162412 77897 162440 79630
rect 162398 77888 162454 77897
rect 162398 77823 162454 77832
rect 162308 77716 162360 77722
rect 162308 77658 162360 77664
rect 162504 76294 162532 79630
rect 162582 79591 162638 79600
rect 162584 79552 162636 79558
rect 162584 79494 162636 79500
rect 162674 79520 162730 79529
rect 162596 78674 162624 79494
rect 162674 79455 162730 79464
rect 162688 79354 162716 79455
rect 162676 79348 162728 79354
rect 162676 79290 162728 79296
rect 162584 78668 162636 78674
rect 162584 78610 162636 78616
rect 162780 78402 162808 79750
rect 162918 79744 162946 80036
rect 163010 79898 163038 80036
rect 163102 79966 163130 80036
rect 163090 79960 163142 79966
rect 163090 79902 163142 79908
rect 162998 79892 163050 79898
rect 162998 79834 163050 79840
rect 163194 79812 163222 80036
rect 163286 79937 163314 80036
rect 163272 79928 163328 79937
rect 163272 79863 163328 79872
rect 163194 79784 163268 79812
rect 163240 79744 163268 79784
rect 162918 79716 163084 79744
rect 162860 79620 162912 79626
rect 162860 79562 162912 79568
rect 162768 78396 162820 78402
rect 162768 78338 162820 78344
rect 162766 78160 162822 78169
rect 162766 78095 162822 78104
rect 162582 77480 162638 77489
rect 162582 77415 162638 77424
rect 162492 76288 162544 76294
rect 162492 76230 162544 76236
rect 162596 75313 162624 77415
rect 162582 75304 162638 75313
rect 162582 75239 162638 75248
rect 162228 74990 162348 75018
rect 162136 70366 162256 70394
rect 162228 12170 162256 70366
rect 162216 12164 162268 12170
rect 162216 12106 162268 12112
rect 162032 11824 162084 11830
rect 162032 11766 162084 11772
rect 161940 8968 161992 8974
rect 161940 8910 161992 8916
rect 162320 6798 162348 74990
rect 162308 6792 162360 6798
rect 162308 6734 162360 6740
rect 161756 6248 161808 6254
rect 161756 6190 161808 6196
rect 162492 4888 162544 4894
rect 162492 4830 162544 4836
rect 161664 3596 161716 3602
rect 161664 3538 161716 3544
rect 161294 3496 161350 3505
rect 161294 3431 161350 3440
rect 161308 480 161336 3431
rect 162504 480 162532 4830
rect 162780 3534 162808 78095
rect 162872 4894 162900 79562
rect 163056 79558 163084 79716
rect 163148 79716 163268 79744
rect 163378 79744 163406 80036
rect 163470 79898 163498 80036
rect 163562 79898 163590 80036
rect 163654 79937 163682 80036
rect 163640 79928 163696 79937
rect 163458 79892 163510 79898
rect 163458 79834 163510 79840
rect 163550 79892 163602 79898
rect 163746 79898 163774 80036
rect 163838 79937 163866 80036
rect 163824 79928 163880 79937
rect 163640 79863 163696 79872
rect 163734 79892 163786 79898
rect 163550 79834 163602 79840
rect 163824 79863 163880 79872
rect 163734 79834 163786 79840
rect 163930 79812 163958 80036
rect 164022 79898 164050 80036
rect 164010 79892 164062 79898
rect 164010 79834 164062 79840
rect 163594 79792 163650 79801
rect 163378 79716 163498 79744
rect 163884 79784 163958 79812
rect 163594 79727 163650 79736
rect 163688 79756 163740 79762
rect 162952 79552 163004 79558
rect 162952 79494 163004 79500
rect 163044 79552 163096 79558
rect 163044 79494 163096 79500
rect 162964 78674 162992 79494
rect 163044 79416 163096 79422
rect 163044 79358 163096 79364
rect 162952 78668 163004 78674
rect 162952 78610 163004 78616
rect 163056 77294 163084 79358
rect 163148 78198 163176 79716
rect 163470 79676 163498 79716
rect 163318 79656 163374 79665
rect 163470 79648 163544 79676
rect 163318 79591 163374 79600
rect 163228 79552 163280 79558
rect 163228 79494 163280 79500
rect 163136 78192 163188 78198
rect 163136 78134 163188 78140
rect 163240 78130 163268 79494
rect 163332 78792 163360 79591
rect 163516 79422 163544 79648
rect 163504 79416 163556 79422
rect 163504 79358 163556 79364
rect 163332 78764 163452 78792
rect 163320 78668 163372 78674
rect 163320 78610 163372 78616
rect 163228 78124 163280 78130
rect 163228 78066 163280 78072
rect 163056 77266 163176 77294
rect 162952 75200 163004 75206
rect 162952 75142 163004 75148
rect 162964 14482 162992 75142
rect 163044 75132 163096 75138
rect 163044 75074 163096 75080
rect 163056 23118 163084 75074
rect 163148 32502 163176 77266
rect 163228 75268 163280 75274
rect 163228 75210 163280 75216
rect 163240 47598 163268 75210
rect 163332 62898 163360 78610
rect 163424 65686 163452 78764
rect 163608 75342 163636 79727
rect 163688 79698 163740 79704
rect 163596 75336 163648 75342
rect 163596 75278 163648 75284
rect 163700 75274 163728 79698
rect 163778 79656 163834 79665
rect 163778 79591 163834 79600
rect 163688 75268 163740 75274
rect 163688 75210 163740 75216
rect 163792 75206 163820 79591
rect 163780 75200 163832 75206
rect 163780 75142 163832 75148
rect 163884 75138 163912 79784
rect 164114 79778 164142 80036
rect 164206 79966 164234 80036
rect 164298 79966 164326 80036
rect 164194 79960 164246 79966
rect 164194 79902 164246 79908
rect 164286 79960 164338 79966
rect 164286 79902 164338 79908
rect 164068 79750 164142 79778
rect 164068 79506 164096 79750
rect 164390 79744 164418 80036
rect 164482 79898 164510 80036
rect 164574 79903 164602 80036
rect 164470 79892 164522 79898
rect 164470 79834 164522 79840
rect 164560 79894 164616 79903
rect 164560 79829 164616 79838
rect 164666 79744 164694 80036
rect 164252 79716 164418 79744
rect 164528 79716 164694 79744
rect 164148 79688 164200 79694
rect 164148 79630 164200 79636
rect 163976 79478 164096 79506
rect 163976 75313 164004 79478
rect 164056 79416 164108 79422
rect 164056 79358 164108 79364
rect 163962 75304 164018 75313
rect 163962 75239 164018 75248
rect 163872 75132 163924 75138
rect 163872 75074 163924 75080
rect 163688 74996 163740 75002
rect 163688 74938 163740 74944
rect 163700 70394 163728 74938
rect 164068 70582 164096 79358
rect 164160 75313 164188 79630
rect 164146 75304 164202 75313
rect 164146 75239 164202 75248
rect 164056 70576 164108 70582
rect 164056 70518 164108 70524
rect 163700 70366 163820 70394
rect 163412 65680 163464 65686
rect 163412 65622 163464 65628
rect 163320 62892 163372 62898
rect 163320 62834 163372 62840
rect 163228 47592 163280 47598
rect 163228 47534 163280 47540
rect 163136 32496 163188 32502
rect 163136 32438 163188 32444
rect 163044 23112 163096 23118
rect 163044 23054 163096 23060
rect 162952 14476 163004 14482
rect 162952 14418 163004 14424
rect 162860 4888 162912 4894
rect 162860 4830 162912 4836
rect 163792 3942 163820 70366
rect 164252 18834 164280 79716
rect 164528 79642 164556 79716
rect 164758 79676 164786 80036
rect 164850 79966 164878 80036
rect 164942 79966 164970 80036
rect 164838 79960 164890 79966
rect 164838 79902 164890 79908
rect 164930 79960 164982 79966
rect 164930 79902 164982 79908
rect 165034 79778 165062 80036
rect 165126 79937 165154 80036
rect 165112 79928 165168 79937
rect 165112 79863 165168 79872
rect 165218 79812 165246 80036
rect 164344 79614 164556 79642
rect 164712 79648 164786 79676
rect 164896 79750 165062 79778
rect 165172 79784 165246 79812
rect 164608 79620 164660 79626
rect 164240 18828 164292 18834
rect 164240 18770 164292 18776
rect 164344 18766 164372 79614
rect 164608 79562 164660 79568
rect 164516 79552 164568 79558
rect 164516 79494 164568 79500
rect 164424 79484 164476 79490
rect 164424 79426 164476 79432
rect 164436 75993 164464 79426
rect 164528 78062 164556 79494
rect 164516 78056 164568 78062
rect 164516 77998 164568 78004
rect 164422 75984 164478 75993
rect 164422 75919 164478 75928
rect 164424 75268 164476 75274
rect 164424 75210 164476 75216
rect 164436 20058 164464 75210
rect 164516 75200 164568 75206
rect 164516 75142 164568 75148
rect 164424 20052 164476 20058
rect 164424 19994 164476 20000
rect 164528 19990 164556 75142
rect 164620 31074 164648 79562
rect 164712 32434 164740 79648
rect 164792 79552 164844 79558
rect 164792 79494 164844 79500
rect 164804 69902 164832 79494
rect 164896 75002 164924 79750
rect 164976 79688 165028 79694
rect 164976 79630 165028 79636
rect 165066 79656 165122 79665
rect 164988 75274 165016 79630
rect 165066 79591 165122 79600
rect 164976 75268 165028 75274
rect 164976 75210 165028 75216
rect 164884 74996 164936 75002
rect 164884 74938 164936 74944
rect 165080 71194 165108 79591
rect 165172 75206 165200 79784
rect 165310 79778 165338 80036
rect 165402 79898 165430 80036
rect 165494 79898 165522 80036
rect 165586 79898 165614 80036
rect 165678 79966 165706 80036
rect 165770 79966 165798 80036
rect 165666 79960 165718 79966
rect 165666 79902 165718 79908
rect 165758 79960 165810 79966
rect 165758 79902 165810 79908
rect 165390 79892 165442 79898
rect 165390 79834 165442 79840
rect 165482 79892 165534 79898
rect 165482 79834 165534 79840
rect 165574 79892 165626 79898
rect 165574 79834 165626 79840
rect 165710 79792 165766 79801
rect 165310 79750 165384 79778
rect 165252 79620 165304 79626
rect 165252 79562 165304 79568
rect 165264 77897 165292 79562
rect 165250 77888 165306 77897
rect 165250 77823 165306 77832
rect 165356 77489 165384 79750
rect 165436 79756 165488 79762
rect 165710 79727 165766 79736
rect 165862 79744 165890 80036
rect 165954 79937 165982 80036
rect 165940 79928 165996 79937
rect 165940 79863 165996 79872
rect 166046 79778 166074 80036
rect 166138 79830 166166 80036
rect 166230 79830 166258 80036
rect 166000 79750 166074 79778
rect 166126 79824 166178 79830
rect 166126 79766 166178 79772
rect 166218 79824 166270 79830
rect 166322 79812 166350 80036
rect 166414 79937 166442 80036
rect 166506 79966 166534 80036
rect 166494 79960 166546 79966
rect 166400 79928 166456 79937
rect 166494 79902 166546 79908
rect 166400 79863 166456 79872
rect 166322 79784 166396 79812
rect 166598 79801 166626 80036
rect 166690 79971 166718 80036
rect 166676 79962 166732 79971
rect 166676 79897 166732 79906
rect 166218 79766 166270 79772
rect 165436 79698 165488 79704
rect 165448 79665 165476 79698
rect 165528 79688 165580 79694
rect 165434 79656 165490 79665
rect 165528 79630 165580 79636
rect 165434 79591 165490 79600
rect 165436 79552 165488 79558
rect 165436 79494 165488 79500
rect 165342 77480 165398 77489
rect 165342 77415 165398 77424
rect 165448 75342 165476 79494
rect 165540 78441 165568 79630
rect 165620 79620 165672 79626
rect 165620 79562 165672 79568
rect 165526 78432 165582 78441
rect 165526 78367 165582 78376
rect 165632 77994 165660 79562
rect 165620 77988 165672 77994
rect 165620 77930 165672 77936
rect 165526 77888 165582 77897
rect 165526 77823 165582 77832
rect 165436 75336 165488 75342
rect 165436 75278 165488 75284
rect 165160 75200 165212 75206
rect 165160 75142 165212 75148
rect 165068 71188 165120 71194
rect 165068 71130 165120 71136
rect 165540 71126 165568 77823
rect 165620 77512 165672 77518
rect 165620 77454 165672 77460
rect 165528 71120 165580 71126
rect 165528 71062 165580 71068
rect 165068 71052 165120 71058
rect 165068 70994 165120 71000
rect 164792 69896 164844 69902
rect 164792 69838 164844 69844
rect 164700 32428 164752 32434
rect 164700 32370 164752 32376
rect 164608 31068 164660 31074
rect 164608 31010 164660 31016
rect 164516 19984 164568 19990
rect 164516 19926 164568 19932
rect 164332 18760 164384 18766
rect 164332 18702 164384 18708
rect 163780 3936 163832 3942
rect 163780 3878 163832 3884
rect 163688 3868 163740 3874
rect 163688 3810 163740 3816
rect 162768 3528 162820 3534
rect 162768 3470 162820 3476
rect 163700 480 163728 3810
rect 164884 3800 164936 3806
rect 164884 3742 164936 3748
rect 164896 480 164924 3742
rect 165080 2990 165108 70994
rect 165632 7614 165660 77454
rect 165724 9518 165752 79727
rect 165862 79716 165936 79744
rect 165804 79212 165856 79218
rect 165804 79154 165856 79160
rect 165816 79082 165844 79154
rect 165804 79076 165856 79082
rect 165804 79018 165856 79024
rect 165804 76628 165856 76634
rect 165804 76570 165856 76576
rect 165816 21554 165844 76570
rect 165908 76226 165936 79716
rect 166000 79642 166028 79750
rect 166000 79614 166120 79642
rect 166368 79626 166396 79784
rect 166584 79792 166640 79801
rect 166448 79756 166500 79762
rect 166782 79744 166810 80036
rect 166874 79966 166902 80036
rect 166966 79971 166994 80036
rect 166862 79960 166914 79966
rect 166862 79902 166914 79908
rect 166952 79962 167008 79971
rect 166952 79897 167008 79906
rect 167058 79778 167086 80036
rect 167150 79812 167178 80036
rect 167242 79937 167270 80036
rect 167228 79928 167284 79937
rect 167228 79863 167284 79872
rect 167150 79784 167224 79812
rect 166584 79727 166640 79736
rect 166448 79698 166500 79704
rect 166736 79716 166810 79744
rect 167012 79750 167086 79778
rect 165988 79552 166040 79558
rect 165988 79494 166040 79500
rect 165896 76220 165948 76226
rect 165896 76162 165948 76168
rect 165896 76084 165948 76090
rect 165896 76026 165948 76032
rect 165804 21548 165856 21554
rect 165804 21490 165856 21496
rect 165908 21486 165936 76026
rect 166000 21622 166028 79494
rect 166092 76634 166120 79614
rect 166264 79620 166316 79626
rect 166264 79562 166316 79568
rect 166356 79620 166408 79626
rect 166356 79562 166408 79568
rect 166172 79552 166224 79558
rect 166172 79494 166224 79500
rect 166184 77518 166212 79494
rect 166276 79472 166304 79562
rect 166276 79444 166396 79472
rect 166264 78668 166316 78674
rect 166264 78610 166316 78616
rect 166276 78334 166304 78610
rect 166264 78328 166316 78334
rect 166264 78270 166316 78276
rect 166172 77512 166224 77518
rect 166172 77454 166224 77460
rect 166264 77512 166316 77518
rect 166264 77454 166316 77460
rect 166080 76628 166132 76634
rect 166080 76570 166132 76576
rect 166078 76528 166134 76537
rect 166078 76463 166134 76472
rect 165988 21616 166040 21622
rect 165988 21558 166040 21564
rect 165896 21480 165948 21486
rect 165896 21422 165948 21428
rect 166092 21418 166120 76463
rect 166172 76220 166224 76226
rect 166172 76162 166224 76168
rect 166184 32570 166212 76162
rect 166276 68474 166304 77454
rect 166368 69834 166396 79444
rect 166460 77518 166488 79698
rect 166540 79620 166592 79626
rect 166540 79562 166592 79568
rect 166448 77512 166500 77518
rect 166448 77454 166500 77460
rect 166552 76090 166580 79562
rect 166632 79348 166684 79354
rect 166632 79290 166684 79296
rect 166644 77314 166672 79290
rect 166736 77353 166764 79716
rect 166816 79620 166868 79626
rect 166816 79562 166868 79568
rect 166828 78441 166856 79562
rect 167012 79404 167040 79750
rect 167092 79620 167144 79626
rect 167092 79562 167144 79568
rect 166920 79376 167040 79404
rect 166920 78606 166948 79376
rect 167104 79336 167132 79562
rect 167012 79308 167132 79336
rect 166908 78600 166960 78606
rect 166908 78542 166960 78548
rect 166814 78432 166870 78441
rect 166814 78367 166870 78376
rect 166814 77480 166870 77489
rect 166814 77415 166870 77424
rect 166722 77344 166778 77353
rect 166632 77308 166684 77314
rect 166722 77279 166778 77288
rect 166632 77250 166684 77256
rect 166540 76084 166592 76090
rect 166540 76026 166592 76032
rect 166828 74534 166856 77415
rect 166736 74506 166856 74534
rect 166736 72826 166764 74506
rect 166724 72820 166776 72826
rect 166724 72762 166776 72768
rect 166356 69828 166408 69834
rect 166356 69770 166408 69776
rect 166264 68468 166316 68474
rect 166264 68410 166316 68416
rect 166172 32564 166224 32570
rect 166172 32506 166224 32512
rect 166080 21412 166132 21418
rect 166080 21354 166132 21360
rect 167012 10334 167040 79308
rect 167092 79212 167144 79218
rect 167092 79154 167144 79160
rect 167104 69766 167132 79154
rect 167196 79082 167224 79784
rect 167334 79744 167362 80036
rect 167288 79716 167362 79744
rect 167426 79744 167454 80036
rect 167518 79812 167546 80036
rect 167610 79937 167638 80036
rect 167596 79928 167652 79937
rect 167702 79898 167730 80036
rect 167596 79863 167652 79872
rect 167690 79892 167742 79898
rect 167690 79834 167742 79840
rect 167518 79784 167592 79812
rect 167426 79716 167500 79744
rect 167288 79218 167316 79716
rect 167368 79484 167420 79490
rect 167368 79426 167420 79432
rect 167276 79212 167328 79218
rect 167276 79154 167328 79160
rect 167380 79150 167408 79426
rect 167368 79144 167420 79150
rect 167368 79086 167420 79092
rect 167184 79076 167236 79082
rect 167184 79018 167236 79024
rect 167184 78940 167236 78946
rect 167184 78882 167236 78888
rect 167276 78940 167328 78946
rect 167276 78882 167328 78888
rect 167196 78538 167224 78882
rect 167184 78532 167236 78538
rect 167184 78474 167236 78480
rect 167182 77752 167238 77761
rect 167182 77687 167184 77696
rect 167236 77687 167238 77696
rect 167184 77658 167236 77664
rect 167184 77512 167236 77518
rect 167184 77454 167236 77460
rect 167092 69760 167144 69766
rect 167092 69702 167144 69708
rect 167092 67108 167144 67114
rect 167092 67050 167144 67056
rect 167104 16574 167132 67050
rect 167196 22914 167224 77454
rect 167288 77382 167316 78882
rect 167368 78260 167420 78266
rect 167368 78202 167420 78208
rect 167276 77376 167328 77382
rect 167276 77318 167328 77324
rect 167276 76832 167328 76838
rect 167276 76774 167328 76780
rect 167184 22908 167236 22914
rect 167184 22850 167236 22856
rect 167288 22846 167316 76774
rect 167380 23050 167408 78202
rect 167368 23044 167420 23050
rect 167368 22986 167420 22992
rect 167472 22982 167500 79716
rect 167564 79200 167592 79784
rect 167794 79744 167822 80036
rect 167886 79830 167914 80036
rect 167978 79898 168006 80036
rect 167966 79892 168018 79898
rect 167966 79834 168018 79840
rect 168070 79830 168098 80036
rect 167874 79824 167926 79830
rect 167874 79766 167926 79772
rect 168058 79824 168110 79830
rect 168162 79801 168190 80036
rect 168254 79812 168282 80036
rect 168346 79937 168374 80036
rect 168438 79966 168466 80036
rect 168426 79960 168478 79966
rect 168332 79928 168388 79937
rect 168426 79902 168478 79908
rect 168530 79898 168558 80036
rect 168622 79966 168650 80036
rect 168714 79971 168742 80036
rect 168610 79960 168662 79966
rect 168610 79902 168662 79908
rect 168700 79962 168756 79971
rect 168806 79966 168834 80036
rect 168332 79863 168388 79872
rect 168518 79892 168570 79898
rect 168700 79897 168756 79906
rect 168794 79960 168846 79966
rect 168794 79902 168846 79908
rect 168518 79834 168570 79840
rect 168898 79812 168926 80036
rect 168058 79766 168110 79772
rect 168148 79792 168204 79801
rect 167656 79716 167822 79744
rect 168254 79784 168328 79812
rect 168148 79727 168204 79736
rect 167656 79626 167684 79716
rect 167920 79688 167972 79694
rect 167920 79630 167972 79636
rect 168104 79688 168156 79694
rect 168104 79630 168156 79636
rect 167644 79620 167696 79626
rect 167644 79562 167696 79568
rect 167736 79620 167788 79626
rect 167736 79562 167788 79568
rect 167828 79620 167880 79626
rect 167828 79562 167880 79568
rect 167564 79172 167684 79200
rect 167552 79076 167604 79082
rect 167552 79018 167604 79024
rect 167564 78266 167592 79018
rect 167552 78260 167604 78266
rect 167552 78202 167604 78208
rect 167550 77344 167606 77353
rect 167550 77279 167606 77288
rect 167564 25566 167592 77279
rect 167656 28286 167684 79172
rect 167748 77518 167776 79562
rect 167736 77512 167788 77518
rect 167736 77454 167788 77460
rect 167840 70394 167868 79562
rect 167932 76838 167960 79630
rect 168012 79212 168064 79218
rect 168012 79154 168064 79160
rect 168024 78674 168052 79154
rect 168012 78668 168064 78674
rect 168012 78610 168064 78616
rect 168010 78024 168066 78033
rect 168010 77959 168066 77968
rect 167920 76832 167972 76838
rect 167920 76774 167972 76780
rect 168024 71058 168052 77959
rect 168116 77625 168144 79630
rect 168300 79200 168328 79784
rect 168852 79784 168926 79812
rect 168380 79756 168432 79762
rect 168380 79698 168432 79704
rect 168208 79172 168328 79200
rect 168102 77616 168158 77625
rect 168102 77551 168158 77560
rect 168208 77353 168236 79172
rect 168392 79150 168420 79698
rect 168472 79688 168524 79694
rect 168472 79630 168524 79636
rect 168380 79144 168432 79150
rect 168380 79086 168432 79092
rect 168288 79076 168340 79082
rect 168288 79018 168340 79024
rect 168300 77790 168328 79018
rect 168378 78704 168434 78713
rect 168378 78639 168380 78648
rect 168432 78639 168434 78648
rect 168380 78610 168432 78616
rect 168378 78432 168434 78441
rect 168378 78367 168434 78376
rect 168392 78169 168420 78367
rect 168378 78160 168434 78169
rect 168378 78095 168434 78104
rect 168288 77784 168340 77790
rect 168288 77726 168340 77732
rect 168484 77722 168512 79630
rect 168564 79620 168616 79626
rect 168564 79562 168616 79568
rect 168472 77716 168524 77722
rect 168472 77658 168524 77664
rect 168576 77602 168604 79562
rect 168656 79144 168708 79150
rect 168656 79086 168708 79092
rect 168484 77574 168604 77602
rect 168194 77344 168250 77353
rect 168194 77279 168250 77288
rect 168012 71052 168064 71058
rect 168012 70994 168064 71000
rect 167748 70366 167868 70394
rect 167748 65618 167776 70366
rect 167736 65612 167788 65618
rect 167736 65554 167788 65560
rect 167644 28280 167696 28286
rect 167644 28222 167696 28228
rect 167552 25560 167604 25566
rect 167552 25502 167604 25508
rect 167460 22976 167512 22982
rect 167460 22918 167512 22924
rect 167276 22840 167328 22846
rect 167276 22782 167328 22788
rect 168484 18698 168512 77574
rect 168668 77489 168696 79086
rect 168748 77716 168800 77722
rect 168748 77658 168800 77664
rect 168654 77480 168710 77489
rect 168654 77415 168710 77424
rect 168564 77376 168616 77382
rect 168564 77318 168616 77324
rect 168472 18692 168524 18698
rect 168472 18634 168524 18640
rect 168576 18630 168604 77318
rect 168760 24546 168788 77658
rect 168852 77382 168880 79784
rect 168990 79744 169018 80036
rect 168944 79716 169018 79744
rect 168944 77500 168972 79716
rect 169082 79676 169110 80036
rect 169174 79830 169202 80036
rect 169266 79898 169294 80036
rect 169254 79892 169306 79898
rect 169254 79834 169306 79840
rect 169162 79824 169214 79830
rect 169358 79812 169386 80036
rect 169450 79937 169478 80036
rect 169436 79928 169492 79937
rect 169436 79863 169492 79872
rect 169358 79784 169432 79812
rect 169162 79766 169214 79772
rect 169300 79688 169352 79694
rect 169082 79648 169156 79676
rect 169024 78260 169076 78266
rect 169024 78202 169076 78208
rect 169036 77568 169064 78202
rect 169128 77704 169156 79648
rect 169300 79630 169352 79636
rect 169208 79620 169260 79626
rect 169208 79562 169260 79568
rect 169220 78266 169248 79562
rect 169208 78260 169260 78266
rect 169208 78202 169260 78208
rect 169128 77676 169248 77704
rect 169036 77540 169156 77568
rect 168944 77472 169064 77500
rect 168840 77376 168892 77382
rect 168840 77318 168892 77324
rect 168932 77376 168984 77382
rect 168932 77318 168984 77324
rect 168840 76832 168892 76838
rect 168840 76774 168892 76780
rect 168748 24540 168800 24546
rect 168748 24482 168800 24488
rect 168852 24410 168880 76774
rect 168944 26926 168972 77318
rect 169036 68406 169064 77472
rect 169128 77382 169156 77540
rect 169116 77376 169168 77382
rect 169116 77318 169168 77324
rect 169116 76628 169168 76634
rect 169116 76570 169168 76576
rect 169128 69698 169156 76570
rect 169220 76566 169248 77676
rect 169208 76560 169260 76566
rect 169208 76502 169260 76508
rect 169312 70394 169340 79630
rect 169404 76838 169432 79784
rect 169542 79744 169570 80036
rect 169496 79716 169570 79744
rect 169634 79744 169662 80036
rect 169726 79971 169754 80036
rect 169712 79962 169768 79971
rect 169712 79897 169768 79906
rect 169818 79898 169846 80036
rect 169910 79966 169938 80036
rect 170002 79966 170030 80036
rect 169898 79960 169950 79966
rect 169898 79902 169950 79908
rect 169990 79960 170042 79966
rect 170094 79937 170122 80036
rect 169990 79902 170042 79908
rect 170080 79928 170136 79937
rect 169806 79892 169858 79898
rect 170186 79898 170214 80036
rect 170278 79966 170306 80036
rect 170370 79971 170398 80036
rect 170266 79960 170318 79966
rect 170266 79902 170318 79908
rect 170356 79962 170412 79971
rect 170080 79863 170136 79872
rect 170174 79892 170226 79898
rect 170356 79897 170412 79906
rect 169806 79834 169858 79840
rect 170174 79834 170226 79840
rect 170462 79778 170490 80036
rect 170554 79898 170582 80036
rect 170542 79892 170594 79898
rect 170542 79834 170594 79840
rect 169760 79756 169812 79762
rect 169634 79716 169708 79744
rect 169392 76832 169444 76838
rect 169392 76774 169444 76780
rect 169496 76634 169524 79716
rect 169576 79620 169628 79626
rect 169576 79562 169628 79568
rect 169484 76628 169536 76634
rect 169484 76570 169536 76576
rect 169588 70394 169616 79562
rect 169680 78849 169708 79716
rect 169760 79698 169812 79704
rect 170128 79756 170180 79762
rect 170462 79750 170536 79778
rect 170128 79698 170180 79704
rect 169666 78840 169722 78849
rect 169666 78775 169722 78784
rect 169668 77512 169720 77518
rect 169668 77454 169720 77460
rect 169680 74534 169708 77454
rect 169772 75138 169800 79698
rect 169944 79688 169996 79694
rect 169944 79630 169996 79636
rect 170034 79656 170090 79665
rect 169852 79620 169904 79626
rect 169852 79562 169904 79568
rect 169760 75132 169812 75138
rect 169760 75074 169812 75080
rect 169680 74506 169800 74534
rect 169312 70366 169524 70394
rect 169588 70366 169708 70394
rect 169116 69692 169168 69698
rect 169116 69634 169168 69640
rect 169024 68400 169076 68406
rect 169024 68342 169076 68348
rect 168932 26920 168984 26926
rect 168932 26862 168984 26868
rect 168840 24404 168892 24410
rect 168840 24346 168892 24352
rect 168564 18624 168616 18630
rect 168564 18566 168616 18572
rect 167104 16546 167224 16574
rect 167000 10328 167052 10334
rect 167000 10270 167052 10276
rect 165712 9512 165764 9518
rect 165712 9454 165764 9460
rect 165620 7608 165672 7614
rect 165620 7550 165672 7556
rect 166080 4820 166132 4826
rect 166080 4762 166132 4768
rect 165068 2984 165120 2990
rect 165068 2926 165120 2932
rect 166092 480 166120 4762
rect 167196 480 167224 16546
rect 169496 4826 169524 70366
rect 169680 24478 169708 70366
rect 169668 24472 169720 24478
rect 169668 24414 169720 24420
rect 169772 11762 169800 74506
rect 169864 24206 169892 79562
rect 169956 24274 169984 79630
rect 170034 79591 170090 79600
rect 170048 79121 170076 79591
rect 170034 79112 170090 79121
rect 170034 79047 170090 79056
rect 170140 77294 170168 79698
rect 170220 79688 170272 79694
rect 170220 79630 170272 79636
rect 170404 79688 170456 79694
rect 170404 79630 170456 79636
rect 170232 77518 170260 79630
rect 170312 79620 170364 79626
rect 170312 79562 170364 79568
rect 170220 77512 170272 77518
rect 170220 77454 170272 77460
rect 170048 77266 170168 77294
rect 170218 77344 170274 77353
rect 170218 77279 170274 77288
rect 169944 24268 169996 24274
rect 169944 24210 169996 24216
rect 169852 24200 169904 24206
rect 169852 24142 169904 24148
rect 170048 24138 170076 77266
rect 170128 75132 170180 75138
rect 170128 75074 170180 75080
rect 170140 64190 170168 75074
rect 170232 65550 170260 77279
rect 170324 73817 170352 79562
rect 170416 77518 170444 79630
rect 170404 77512 170456 77518
rect 170404 77454 170456 77460
rect 170508 76401 170536 79750
rect 170646 79744 170674 80036
rect 170738 79830 170766 80036
rect 170726 79824 170778 79830
rect 170726 79766 170778 79772
rect 170600 79716 170674 79744
rect 170600 78112 170628 79716
rect 170830 79540 170858 80036
rect 170922 79801 170950 80036
rect 171014 79937 171042 80036
rect 171000 79928 171056 79937
rect 171000 79863 171056 79872
rect 171106 79830 171134 80036
rect 171094 79824 171146 79830
rect 170908 79792 170964 79801
rect 171094 79766 171146 79772
rect 171198 79778 171226 80036
rect 171290 79937 171318 80036
rect 171276 79928 171332 79937
rect 171276 79863 171332 79872
rect 171382 79778 171410 80036
rect 171474 79830 171502 80036
rect 171198 79750 171272 79778
rect 171336 79762 171410 79778
rect 171462 79824 171514 79830
rect 171462 79766 171514 79772
rect 170908 79727 170964 79736
rect 171244 79694 171272 79750
rect 171324 79756 171410 79762
rect 171376 79750 171410 79756
rect 171324 79698 171376 79704
rect 171140 79688 171192 79694
rect 171140 79630 171192 79636
rect 171232 79688 171284 79694
rect 171566 79676 171594 80036
rect 171232 79630 171284 79636
rect 171520 79648 171594 79676
rect 170784 79512 170858 79540
rect 170784 78305 170812 79512
rect 171048 79348 171100 79354
rect 171048 79290 171100 79296
rect 171060 79218 171088 79290
rect 171048 79212 171100 79218
rect 171048 79154 171100 79160
rect 170954 79112 171010 79121
rect 170954 79047 171010 79056
rect 170862 78976 170918 78985
rect 170862 78911 170918 78920
rect 170876 78538 170904 78911
rect 170864 78532 170916 78538
rect 170864 78474 170916 78480
rect 170770 78296 170826 78305
rect 170770 78231 170826 78240
rect 170600 78084 170720 78112
rect 170692 77994 170720 78084
rect 170770 78024 170826 78033
rect 170588 77988 170640 77994
rect 170588 77930 170640 77936
rect 170680 77988 170732 77994
rect 170770 77959 170826 77968
rect 170680 77930 170732 77936
rect 170494 76392 170550 76401
rect 170494 76327 170550 76336
rect 170310 73808 170366 73817
rect 170310 73743 170366 73752
rect 170404 70576 170456 70582
rect 170404 70518 170456 70524
rect 170220 65544 170272 65550
rect 170220 65486 170272 65492
rect 170128 64184 170180 64190
rect 170128 64126 170180 64132
rect 170036 24132 170088 24138
rect 170036 24074 170088 24080
rect 169760 11756 169812 11762
rect 169760 11698 169812 11704
rect 169576 5160 169628 5166
rect 169576 5102 169628 5108
rect 169484 4820 169536 4826
rect 169484 4762 169536 4768
rect 168380 3460 168432 3466
rect 168380 3402 168432 3408
rect 168392 480 168420 3402
rect 169588 480 169616 5102
rect 170416 3505 170444 70518
rect 170600 70394 170628 77930
rect 170600 70366 170720 70394
rect 170692 62830 170720 70366
rect 170784 68338 170812 77959
rect 170864 73160 170916 73166
rect 170968 73154 170996 79047
rect 171152 78305 171180 79630
rect 171324 79620 171376 79626
rect 171324 79562 171376 79568
rect 171232 79416 171284 79422
rect 171232 79358 171284 79364
rect 171138 78296 171194 78305
rect 171138 78231 171194 78240
rect 171244 76770 171272 79358
rect 171336 77926 171364 79562
rect 171520 79121 171548 79648
rect 171658 79608 171686 80036
rect 171750 79971 171778 80036
rect 171736 79962 171792 79971
rect 171736 79897 171792 79906
rect 171842 79744 171870 80036
rect 171934 79812 171962 80036
rect 172026 79966 172054 80036
rect 172014 79960 172066 79966
rect 172014 79902 172066 79908
rect 171934 79784 172008 79812
rect 171842 79716 171916 79744
rect 171888 79665 171916 79716
rect 171612 79580 171686 79608
rect 171874 79656 171930 79665
rect 171874 79591 171930 79600
rect 171506 79112 171562 79121
rect 171506 79047 171562 79056
rect 171508 78804 171560 78810
rect 171508 78746 171560 78752
rect 171324 77920 171376 77926
rect 171324 77862 171376 77868
rect 171232 76764 171284 76770
rect 171232 76706 171284 76712
rect 171046 76256 171102 76265
rect 171046 76191 171102 76200
rect 170916 73126 170996 73154
rect 170864 73102 170916 73108
rect 170772 68332 170824 68338
rect 170772 68274 170824 68280
rect 170680 62824 170732 62830
rect 170680 62766 170732 62772
rect 171060 6186 171088 76191
rect 171520 75070 171548 78746
rect 171612 77858 171640 79580
rect 171876 79552 171928 79558
rect 171876 79494 171928 79500
rect 171784 79484 171836 79490
rect 171784 79426 171836 79432
rect 171796 78441 171824 79426
rect 171888 79354 171916 79494
rect 171876 79348 171928 79354
rect 171876 79290 171928 79296
rect 171980 78810 172008 79784
rect 172118 79778 172146 80036
rect 172210 79971 172238 80036
rect 172196 79962 172252 79971
rect 172196 79897 172252 79906
rect 172072 79750 172146 79778
rect 171968 78804 172020 78810
rect 171968 78746 172020 78752
rect 171968 78600 172020 78606
rect 171968 78542 172020 78548
rect 171876 78532 171928 78538
rect 171876 78474 171928 78480
rect 171782 78432 171838 78441
rect 171782 78367 171838 78376
rect 171888 78334 171916 78474
rect 171876 78328 171928 78334
rect 171876 78270 171928 78276
rect 171980 78130 172008 78542
rect 172072 78334 172100 79750
rect 172302 79744 172330 80036
rect 172394 79966 172422 80036
rect 172382 79960 172434 79966
rect 172382 79902 172434 79908
rect 172256 79716 172330 79744
rect 172152 79688 172204 79694
rect 172152 79630 172204 79636
rect 172164 78962 172192 79630
rect 172256 79490 172284 79716
rect 172486 79676 172514 80036
rect 172578 79812 172606 80036
rect 172670 79966 172698 80036
rect 172762 79966 172790 80036
rect 172658 79960 172710 79966
rect 172658 79902 172710 79908
rect 172750 79960 172802 79966
rect 172854 79937 172882 80036
rect 172946 79966 172974 80036
rect 172934 79960 172986 79966
rect 172750 79902 172802 79908
rect 172840 79928 172896 79937
rect 172934 79902 172986 79908
rect 172840 79863 172896 79872
rect 173038 79812 173066 80036
rect 173130 79966 173158 80036
rect 173118 79960 173170 79966
rect 173222 79937 173250 80036
rect 173118 79902 173170 79908
rect 173208 79928 173264 79937
rect 173314 79898 173342 80036
rect 173406 79971 173434 80036
rect 173392 79962 173448 79971
rect 173208 79863 173264 79872
rect 173302 79892 173354 79898
rect 173392 79897 173448 79906
rect 173302 79834 173354 79840
rect 173498 79812 173526 80036
rect 173590 79966 173618 80036
rect 173682 79966 173710 80036
rect 173774 79966 173802 80036
rect 173866 79966 173894 80036
rect 173578 79960 173630 79966
rect 173578 79902 173630 79908
rect 173670 79960 173722 79966
rect 173670 79902 173722 79908
rect 173762 79960 173814 79966
rect 173762 79902 173814 79908
rect 173854 79960 173906 79966
rect 173854 79902 173906 79908
rect 173808 79824 173860 79830
rect 172578 79784 172744 79812
rect 173038 79784 173204 79812
rect 172612 79688 172664 79694
rect 172486 79648 172560 79676
rect 172336 79620 172388 79626
rect 172336 79562 172388 79568
rect 172244 79484 172296 79490
rect 172244 79426 172296 79432
rect 172348 79286 172376 79562
rect 172428 79552 172480 79558
rect 172428 79494 172480 79500
rect 172336 79280 172388 79286
rect 172336 79222 172388 79228
rect 172164 78934 172284 78962
rect 172256 78878 172284 78934
rect 172152 78872 172204 78878
rect 172152 78814 172204 78820
rect 172244 78872 172296 78878
rect 172244 78814 172296 78820
rect 172060 78328 172112 78334
rect 172060 78270 172112 78276
rect 171784 78124 171836 78130
rect 171784 78066 171836 78072
rect 171968 78124 172020 78130
rect 171968 78066 172020 78072
rect 171600 77852 171652 77858
rect 171600 77794 171652 77800
rect 171600 77716 171652 77722
rect 171600 77658 171652 77664
rect 171508 75064 171560 75070
rect 171508 75006 171560 75012
rect 171612 70394 171640 77658
rect 171796 77314 171824 78066
rect 172164 78010 172192 78814
rect 172440 78810 172468 79494
rect 172532 78810 172560 79648
rect 172612 79630 172664 79636
rect 172428 78804 172480 78810
rect 172428 78746 172480 78752
rect 172520 78804 172572 78810
rect 172520 78746 172572 78752
rect 172624 78606 172652 79630
rect 172612 78600 172664 78606
rect 172612 78542 172664 78548
rect 171980 77982 172192 78010
rect 171874 77888 171930 77897
rect 171874 77823 171930 77832
rect 171784 77308 171836 77314
rect 171784 77250 171836 77256
rect 171784 76628 171836 76634
rect 171784 76570 171836 76576
rect 171796 76294 171824 76570
rect 171784 76288 171836 76294
rect 171784 76230 171836 76236
rect 171888 76106 171916 77823
rect 171796 76078 171916 76106
rect 171612 70366 171732 70394
rect 171704 26994 171732 70366
rect 171796 28354 171824 76078
rect 171980 75970 172008 77982
rect 172716 77926 172744 79784
rect 172888 79756 172940 79762
rect 172888 79698 172940 79704
rect 172704 77920 172756 77926
rect 172704 77862 172756 77868
rect 172152 77784 172204 77790
rect 172152 77726 172204 77732
rect 172060 77580 172112 77586
rect 172060 77522 172112 77528
rect 171888 75942 172008 75970
rect 171784 28348 171836 28354
rect 171784 28290 171836 28296
rect 171692 26988 171744 26994
rect 171692 26930 171744 26936
rect 171048 6180 171100 6186
rect 171048 6122 171100 6128
rect 170772 3664 170824 3670
rect 170772 3606 170824 3612
rect 170402 3496 170458 3505
rect 170402 3431 170458 3440
rect 170784 480 170812 3606
rect 171888 3194 171916 75942
rect 171966 75168 172022 75177
rect 171966 75103 172022 75112
rect 171980 33114 172008 75103
rect 171968 33108 172020 33114
rect 171968 33050 172020 33056
rect 172072 3466 172100 77522
rect 172164 36582 172192 77726
rect 172242 77616 172298 77625
rect 172242 77551 172298 77560
rect 172152 36576 172204 36582
rect 172152 36518 172204 36524
rect 172256 23186 172284 77551
rect 172336 77512 172388 77518
rect 172336 77454 172388 77460
rect 172244 23180 172296 23186
rect 172244 23122 172296 23128
rect 172348 4146 172376 77454
rect 172900 77217 172928 79698
rect 173176 79529 173204 79784
rect 173346 79792 173402 79801
rect 173256 79756 173308 79762
rect 173498 79784 173572 79812
rect 173346 79727 173402 79736
rect 173256 79698 173308 79704
rect 173162 79520 173218 79529
rect 173162 79455 173218 79464
rect 173268 79257 173296 79698
rect 173360 79393 173388 79727
rect 173440 79688 173492 79694
rect 173440 79630 173492 79636
rect 173346 79384 173402 79393
rect 173346 79319 173402 79328
rect 173254 79248 173310 79257
rect 173254 79183 173310 79192
rect 173452 78849 173480 79630
rect 173544 79422 173572 79784
rect 173808 79766 173860 79772
rect 173624 79756 173676 79762
rect 173624 79698 173676 79704
rect 173716 79756 173768 79762
rect 173716 79698 173768 79704
rect 173532 79416 173584 79422
rect 173532 79358 173584 79364
rect 173438 78840 173494 78849
rect 173438 78775 173494 78784
rect 173636 78713 173664 79698
rect 173728 78985 173756 79698
rect 173714 78976 173770 78985
rect 173714 78911 173770 78920
rect 173622 78704 173678 78713
rect 173820 78674 173848 79766
rect 173958 79744 173986 80036
rect 173912 79716 173986 79744
rect 173622 78639 173678 78648
rect 173808 78668 173860 78674
rect 173808 78610 173860 78616
rect 173912 78577 173940 79716
rect 174050 79676 174078 80036
rect 174142 79778 174170 80036
rect 174234 79880 174262 80036
rect 174326 79948 174354 80036
rect 174326 79920 174400 79948
rect 174234 79852 174308 79880
rect 174142 79750 174216 79778
rect 174004 79648 174078 79676
rect 174004 79354 174032 79648
rect 173992 79348 174044 79354
rect 173992 79290 174044 79296
rect 173898 78568 173954 78577
rect 173898 78503 173954 78512
rect 174188 78441 174216 79750
rect 174174 78432 174230 78441
rect 174174 78367 174230 78376
rect 172886 77208 172942 77217
rect 172886 77143 172942 77152
rect 173162 77072 173218 77081
rect 173162 77007 173218 77016
rect 172520 76356 172572 76362
rect 172520 76298 172572 76304
rect 172532 75886 172560 76298
rect 172520 75880 172572 75886
rect 172520 75822 172572 75828
rect 172428 75064 172480 75070
rect 172428 75006 172480 75012
rect 172336 4140 172388 4146
rect 172336 4082 172388 4088
rect 172440 3806 172468 75006
rect 173176 5250 173204 77007
rect 173346 76936 173402 76945
rect 173346 76871 173402 76880
rect 173256 75948 173308 75954
rect 173256 75890 173308 75896
rect 173268 5386 173296 75890
rect 173360 5522 173388 76871
rect 173992 76832 174044 76838
rect 173992 76774 174044 76780
rect 173898 75848 173954 75857
rect 173898 75783 173954 75792
rect 173532 74928 173584 74934
rect 173532 74870 173584 74876
rect 173544 70242 173572 74870
rect 173440 70236 173492 70242
rect 173440 70178 173492 70184
rect 173532 70236 173584 70242
rect 173532 70178 173584 70184
rect 173452 16574 173480 70178
rect 173452 16546 173756 16574
rect 173360 5494 173664 5522
rect 173268 5358 173480 5386
rect 173176 5222 173296 5250
rect 172428 3800 172480 3806
rect 172428 3742 172480 3748
rect 172060 3460 172112 3466
rect 172060 3402 172112 3408
rect 173268 3398 173296 5222
rect 173256 3392 173308 3398
rect 173256 3334 173308 3340
rect 173452 3330 173480 5358
rect 173636 3874 173664 5494
rect 173624 3868 173676 3874
rect 173624 3810 173676 3816
rect 173164 3324 173216 3330
rect 173164 3266 173216 3272
rect 173440 3324 173492 3330
rect 173440 3266 173492 3272
rect 171876 3188 171928 3194
rect 171876 3130 171928 3136
rect 171968 2984 172020 2990
rect 171968 2926 172020 2932
rect 171980 480 172008 2926
rect 173176 480 173204 3266
rect 173728 3126 173756 16546
rect 173716 3120 173768 3126
rect 173716 3062 173768 3068
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 173912 354 173940 75783
rect 174004 23254 174032 76774
rect 174280 74534 174308 79852
rect 174372 76838 174400 79920
rect 174464 76838 174492 80378
rect 174544 80300 174596 80306
rect 174544 80242 174596 80248
rect 174556 79898 174584 80242
rect 174636 80232 174688 80238
rect 174636 80174 174688 80180
rect 174544 79892 174596 79898
rect 174544 79834 174596 79840
rect 174648 79218 174676 80174
rect 174740 79966 174768 80582
rect 174832 80170 174860 80582
rect 174912 80368 174964 80374
rect 174912 80310 174964 80316
rect 174924 80170 174952 80310
rect 174820 80164 174872 80170
rect 174820 80106 174872 80112
rect 174912 80164 174964 80170
rect 174912 80106 174964 80112
rect 174728 79960 174780 79966
rect 174728 79902 174780 79908
rect 175016 79665 175044 80582
rect 176108 80504 176160 80510
rect 176108 80446 176160 80452
rect 175464 80096 175516 80102
rect 175464 80038 175516 80044
rect 175556 80096 175608 80102
rect 176120 80073 176148 80446
rect 176384 80300 176436 80306
rect 176384 80242 176436 80248
rect 175556 80038 175608 80044
rect 176106 80064 176162 80073
rect 175002 79656 175058 79665
rect 175002 79591 175058 79600
rect 174636 79212 174688 79218
rect 174636 79154 174688 79160
rect 174728 79212 174780 79218
rect 174728 79154 174780 79160
rect 174740 78878 174768 79154
rect 174728 78872 174780 78878
rect 174728 78814 174780 78820
rect 175476 78033 175504 80038
rect 175568 79898 175596 80038
rect 176106 79999 176162 80008
rect 175556 79892 175608 79898
rect 175556 79834 175608 79840
rect 176292 79416 176344 79422
rect 176292 79358 176344 79364
rect 176200 79348 176252 79354
rect 176200 79290 176252 79296
rect 176212 79121 176240 79290
rect 176198 79112 176254 79121
rect 176198 79047 176254 79056
rect 176198 78160 176254 78169
rect 176198 78095 176254 78104
rect 175462 78024 175518 78033
rect 175462 77959 175518 77968
rect 176212 77722 176240 78095
rect 176304 77858 176332 79358
rect 176292 77852 176344 77858
rect 176292 77794 176344 77800
rect 176200 77716 176252 77722
rect 176200 77658 176252 77664
rect 176396 77450 176424 80242
rect 178604 80034 178632 80718
rect 178592 80028 178644 80034
rect 178592 79970 178644 79976
rect 176752 78872 176804 78878
rect 176752 78814 176804 78820
rect 176764 78606 176792 78814
rect 176752 78600 176804 78606
rect 176752 78542 176804 78548
rect 178776 78328 178828 78334
rect 178776 78270 178828 78276
rect 176384 77444 176436 77450
rect 176384 77386 176436 77392
rect 178788 77353 178816 78270
rect 178774 77344 178830 77353
rect 178774 77279 178830 77288
rect 174360 76832 174412 76838
rect 174360 76774 174412 76780
rect 174452 76832 174504 76838
rect 174452 76774 174504 76780
rect 174188 74506 174308 74534
rect 174188 70394 174216 74506
rect 174096 70366 174216 70394
rect 174096 45558 174124 70366
rect 175278 68504 175334 68513
rect 175278 68439 175334 68448
rect 174084 45552 174136 45558
rect 174084 45494 174136 45500
rect 173992 23248 174044 23254
rect 173992 23190 174044 23196
rect 175292 16574 175320 68439
rect 176658 32600 176714 32609
rect 176658 32535 176714 32544
rect 175292 16546 175504 16574
rect 175476 480 175504 16546
rect 176672 3670 176700 32535
rect 176752 26036 176804 26042
rect 176752 25978 176804 25984
rect 176660 3664 176712 3670
rect 176660 3606 176712 3612
rect 176764 3482 176792 25978
rect 179420 25968 179472 25974
rect 179420 25910 179472 25916
rect 179432 16574 179460 25910
rect 179892 24342 179920 130455
rect 180076 79558 180104 536794
rect 180156 111852 180208 111858
rect 180156 111794 180208 111800
rect 180064 79552 180116 79558
rect 180064 79494 180116 79500
rect 180168 78305 180196 111794
rect 180812 110673 180840 700266
rect 184204 683188 184256 683194
rect 184204 683130 184256 683136
rect 180892 670744 180944 670750
rect 180892 670686 180944 670692
rect 180904 113393 180932 670686
rect 182824 643136 182876 643142
rect 182824 643078 182876 643084
rect 180984 618316 181036 618322
rect 180984 618258 181036 618264
rect 180996 114753 181024 618258
rect 181076 514820 181128 514826
rect 181076 514762 181128 514768
rect 181088 117473 181116 514762
rect 181168 357468 181220 357474
rect 181168 357410 181220 357416
rect 181180 121553 181208 357410
rect 182180 305040 182232 305046
rect 182180 304982 182232 304988
rect 181444 142928 181496 142934
rect 181444 142870 181496 142876
rect 181352 141568 181404 141574
rect 181352 141510 181404 141516
rect 181258 129704 181314 129713
rect 181258 129639 181314 129648
rect 181166 121544 181222 121553
rect 181166 121479 181222 121488
rect 181074 117464 181130 117473
rect 181074 117399 181130 117408
rect 180982 114744 181038 114753
rect 180982 114679 181038 114688
rect 180890 113384 180946 113393
rect 180890 113319 180946 113328
rect 180798 110664 180854 110673
rect 180798 110599 180854 110608
rect 180154 78296 180210 78305
rect 180154 78231 180210 78240
rect 181272 59362 181300 129639
rect 181364 80510 181392 141510
rect 181456 109313 181484 142870
rect 181536 139460 181588 139466
rect 181536 139402 181588 139408
rect 181548 128353 181576 139402
rect 181534 128344 181590 128353
rect 181534 128279 181590 128288
rect 182192 122913 182220 304982
rect 182272 139392 182324 139398
rect 182272 139334 182324 139340
rect 182284 124273 182312 139334
rect 182364 139324 182416 139330
rect 182364 139266 182416 139272
rect 182376 125633 182404 139266
rect 182362 125624 182418 125633
rect 182362 125559 182418 125568
rect 182270 124264 182326 124273
rect 182270 124199 182326 124208
rect 182178 122904 182234 122913
rect 182178 122839 182234 122848
rect 181442 109304 181498 109313
rect 181442 109239 181498 109248
rect 182732 104848 182784 104854
rect 182732 104790 182784 104796
rect 182744 103873 182772 104790
rect 182730 103864 182786 103873
rect 182730 103799 182786 103808
rect 182272 101516 182324 101522
rect 182272 101458 182324 101464
rect 182284 101153 182312 101458
rect 182270 101144 182326 101153
rect 182270 101079 182326 101088
rect 182456 100020 182508 100026
rect 182456 99962 182508 99968
rect 182468 99793 182496 99962
rect 182454 99784 182510 99793
rect 182454 99719 182510 99728
rect 182180 98524 182232 98530
rect 182180 98466 182232 98472
rect 182192 98433 182220 98466
rect 182178 98424 182234 98433
rect 182178 98359 182234 98368
rect 182548 97436 182600 97442
rect 182548 97378 182600 97384
rect 182560 97073 182588 97378
rect 182546 97064 182602 97073
rect 182546 96999 182602 97008
rect 182548 93152 182600 93158
rect 182548 93094 182600 93100
rect 182560 91633 182588 93094
rect 182546 91624 182602 91633
rect 182546 91559 182602 91568
rect 181352 80504 181404 80510
rect 181352 80446 181404 80452
rect 182836 77353 182864 643078
rect 182916 484424 182968 484430
rect 182916 484366 182968 484372
rect 182928 77722 182956 484366
rect 183008 418192 183060 418198
rect 183008 418134 183060 418140
rect 183020 92993 183048 418134
rect 183100 271924 183152 271930
rect 183100 271866 183152 271872
rect 183006 92984 183062 92993
rect 183006 92919 183062 92928
rect 183006 80744 183062 80753
rect 183006 80679 183062 80688
rect 182916 77716 182968 77722
rect 182916 77658 182968 77664
rect 182822 77344 182878 77353
rect 182822 77279 182878 77288
rect 181444 72820 181496 72826
rect 181444 72762 181496 72768
rect 181260 59356 181312 59362
rect 181260 59298 181312 59304
rect 179880 24336 179932 24342
rect 179880 24278 179932 24284
rect 181456 16574 181484 72762
rect 183020 24342 183048 80679
rect 183112 79286 183140 271866
rect 183192 151836 183244 151842
rect 183192 151778 183244 151784
rect 183100 79280 183152 79286
rect 183100 79222 183152 79228
rect 183204 79218 183232 151778
rect 183468 108996 183520 109002
rect 183468 108938 183520 108944
rect 183480 107953 183508 108938
rect 183466 107944 183522 107953
rect 183466 107879 183522 107888
rect 183468 107636 183520 107642
rect 183468 107578 183520 107584
rect 183480 106593 183508 107578
rect 183466 106584 183522 106593
rect 183466 106519 183522 106528
rect 183468 106276 183520 106282
rect 183468 106218 183520 106224
rect 183480 105233 183508 106218
rect 183466 105224 183522 105233
rect 183466 105159 183522 105168
rect 183468 102672 183520 102678
rect 183468 102614 183520 102620
rect 183480 102513 183508 102614
rect 183466 102504 183522 102513
rect 183466 102439 183522 102448
rect 184216 100026 184244 683130
rect 184296 630692 184348 630698
rect 184296 630634 184348 630640
rect 184204 100020 184256 100026
rect 184204 99962 184256 99968
rect 184308 98530 184336 630634
rect 184388 576904 184440 576910
rect 184388 576846 184440 576852
rect 184296 98524 184348 98530
rect 184296 98466 184348 98472
rect 184400 97442 184428 576846
rect 185596 101522 185624 700266
rect 188356 102678 188384 700334
rect 189736 104854 189764 700402
rect 192496 106282 192524 700470
rect 193876 107642 193904 700538
rect 196636 109002 196664 700606
rect 196716 138032 196768 138038
rect 196716 137974 196768 137980
rect 196624 108996 196676 109002
rect 196624 108938 196676 108944
rect 193864 107636 193916 107642
rect 193864 107578 193916 107584
rect 192484 106276 192536 106282
rect 192484 106218 192536 106224
rect 189724 104848 189776 104854
rect 189724 104790 189776 104796
rect 188344 102672 188396 102678
rect 188344 102614 188396 102620
rect 185584 101516 185636 101522
rect 185584 101458 185636 101464
rect 193864 99408 193916 99414
rect 193864 99350 193916 99356
rect 184388 97436 184440 97442
rect 184388 97378 184440 97384
rect 183468 96620 183520 96626
rect 183468 96562 183520 96568
rect 183480 95713 183508 96562
rect 183466 95704 183522 95713
rect 183466 95639 183522 95648
rect 183468 95192 183520 95198
rect 183468 95134 183520 95140
rect 183480 94353 183508 95134
rect 183466 94344 183522 94353
rect 183466 94279 183522 94288
rect 183468 91792 183520 91798
rect 183468 91734 183520 91740
rect 183376 90364 183428 90370
rect 183376 90306 183428 90312
rect 183388 88913 183416 90306
rect 183480 90273 183508 91734
rect 183466 90264 183522 90273
rect 183466 90199 183522 90208
rect 183468 89004 183520 89010
rect 183468 88946 183520 88952
rect 183374 88904 183430 88913
rect 183374 88839 183430 88848
rect 183376 87644 183428 87650
rect 183376 87586 183428 87592
rect 183388 86193 183416 87586
rect 183480 87553 183508 88946
rect 183466 87544 183522 87553
rect 183466 87479 183522 87488
rect 183374 86184 183430 86193
rect 183374 86119 183430 86128
rect 183468 85536 183520 85542
rect 183468 85478 183520 85484
rect 183480 84833 183508 85478
rect 183466 84824 183522 84833
rect 183466 84759 183522 84768
rect 193876 84182 193904 99350
rect 196728 85542 196756 137974
rect 196716 85536 196768 85542
rect 196716 85478 196768 85484
rect 183468 84176 183520 84182
rect 183468 84118 183520 84124
rect 193864 84176 193916 84182
rect 193864 84118 193916 84124
rect 183480 83473 183508 84118
rect 183466 83464 183522 83473
rect 183466 83399 183522 83408
rect 183282 82104 183338 82113
rect 183282 82039 183338 82048
rect 183192 79212 183244 79218
rect 183192 79154 183244 79160
rect 183296 60722 183324 82039
rect 200120 80300 200172 80306
rect 200120 80242 200172 80248
rect 195980 79076 196032 79082
rect 195980 79018 196032 79024
rect 193862 75712 193918 75721
rect 193862 75647 193918 75656
rect 189080 74316 189132 74322
rect 189080 74258 189132 74264
rect 189092 71670 189120 74258
rect 193876 73710 193904 75647
rect 194598 74488 194654 74497
rect 194598 74423 194654 74432
rect 193864 73704 193916 73710
rect 193864 73646 193916 73652
rect 189080 71664 189132 71670
rect 189080 71606 189132 71612
rect 190460 70984 190512 70990
rect 190460 70926 190512 70932
rect 189080 67040 189132 67046
rect 189080 66982 189132 66988
rect 184940 63164 184992 63170
rect 184940 63106 184992 63112
rect 183284 60716 183336 60722
rect 183284 60658 183336 60664
rect 183560 25900 183612 25906
rect 183560 25842 183612 25848
rect 183008 24336 183060 24342
rect 183008 24278 183060 24284
rect 183572 16574 183600 25842
rect 179432 16546 180288 16574
rect 181456 16546 181576 16574
rect 183572 16546 183784 16574
rect 177856 3664 177908 3670
rect 177856 3606 177908 3612
rect 177948 3664 178000 3670
rect 177948 3606 178000 3612
rect 176672 3454 176792 3482
rect 176672 480 176700 3454
rect 177868 480 177896 3606
rect 177960 3398 177988 3606
rect 179052 3460 179104 3466
rect 179052 3402 179104 3408
rect 177948 3392 178000 3398
rect 177948 3334 178000 3340
rect 179064 480 179092 3402
rect 180260 480 180288 16546
rect 181548 3466 181576 16546
rect 181444 3460 181496 3466
rect 181444 3402 181496 3408
rect 181536 3460 181588 3466
rect 181536 3402 181588 3408
rect 181456 480 181484 3402
rect 182548 3120 182600 3126
rect 182548 3062 182600 3068
rect 182560 480 182588 3062
rect 183756 480 183784 16546
rect 184952 4214 184980 63106
rect 185032 44872 185084 44878
rect 185032 44814 185084 44820
rect 184940 4208 184992 4214
rect 184940 4150 184992 4156
rect 185044 3482 185072 44814
rect 187700 32768 187752 32774
rect 187700 32710 187752 32716
rect 186320 25832 186372 25838
rect 186320 25774 186372 25780
rect 186332 16574 186360 25774
rect 187712 16574 187740 32710
rect 189092 16574 189120 66982
rect 186332 16546 186912 16574
rect 187712 16546 188568 16574
rect 189092 16546 189304 16574
rect 186136 4208 186188 4214
rect 186136 4150 186188 4156
rect 184952 3454 185072 3482
rect 184952 480 184980 3454
rect 186148 480 186176 4150
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 188540 480 188568 16546
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189276 354 189304 16546
rect 189694 354 189806 480
rect 189276 326 189806 354
rect 190472 354 190500 70926
rect 193218 68368 193274 68377
rect 193218 68303 193274 68312
rect 191838 34096 191894 34105
rect 191838 34031 191894 34040
rect 191852 16574 191880 34031
rect 191852 16546 192064 16574
rect 192036 480 192064 16546
rect 193232 480 193260 68303
rect 193310 25528 193366 25537
rect 193310 25463 193366 25472
rect 193324 16574 193352 25463
rect 194612 16574 194640 74423
rect 195992 16574 196020 79018
rect 197360 76424 197412 76430
rect 197360 76366 197412 76372
rect 197372 16574 197400 76366
rect 198740 33992 198792 33998
rect 198740 33934 198792 33940
rect 193324 16546 194456 16574
rect 194612 16546 195192 16574
rect 195992 16546 196848 16574
rect 197372 16546 197952 16574
rect 194428 480 194456 16546
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 189694 -960 189806 326
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 196820 480 196848 16546
rect 197924 480 197952 16546
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 33934
rect 200132 16574 200160 80242
rect 201512 79626 201540 702986
rect 218992 700670 219020 703520
rect 218980 700664 219032 700670
rect 218980 700606 219032 700612
rect 214564 524476 214616 524482
rect 214564 524418 214616 524424
rect 211804 470620 211856 470626
rect 211804 470562 211856 470568
rect 211816 95198 211844 470562
rect 214576 96626 214604 524418
rect 224224 364404 224276 364410
rect 224224 364346 224276 364352
rect 221464 311908 221516 311914
rect 221464 311850 221516 311856
rect 220084 258120 220136 258126
rect 220084 258062 220136 258068
rect 217324 218068 217376 218074
rect 217324 218010 217376 218016
rect 215944 178084 215996 178090
rect 215944 178026 215996 178032
rect 214564 96620 214616 96626
rect 214564 96562 214616 96568
rect 211804 95192 211856 95198
rect 211804 95134 211856 95140
rect 215956 87650 215984 178026
rect 217336 89010 217364 218010
rect 220096 90370 220124 258062
rect 221476 91798 221504 311850
rect 224236 93158 224264 364346
rect 234632 145654 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 697610 267688 703520
rect 283852 700602 283880 703520
rect 283840 700596 283892 700602
rect 283840 700538 283892 700544
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 234620 145648 234672 145654
rect 234620 145590 234672 145596
rect 224224 93152 224276 93158
rect 224224 93094 224276 93100
rect 221464 91792 221516 91798
rect 221464 91734 221516 91740
rect 220084 90364 220136 90370
rect 220084 90306 220136 90312
rect 217324 89004 217376 89010
rect 217324 88946 217376 88952
rect 215944 87644 215996 87650
rect 215944 87586 215996 87592
rect 231860 80232 231912 80238
rect 231860 80174 231912 80180
rect 201500 79620 201552 79626
rect 201500 79562 201552 79568
rect 213920 78940 213972 78946
rect 213920 78882 213972 78888
rect 208400 76492 208452 76498
rect 208400 76434 208452 76440
rect 208412 74322 208440 76434
rect 208400 74316 208452 74322
rect 208400 74258 208452 74264
rect 209780 73772 209832 73778
rect 209780 73714 209832 73720
rect 207020 60172 207072 60178
rect 207020 60114 207072 60120
rect 205640 33924 205692 33930
rect 205640 33866 205692 33872
rect 201500 32700 201552 32706
rect 201500 32642 201552 32648
rect 200132 16546 200344 16574
rect 200316 480 200344 16546
rect 201512 4214 201540 32642
rect 204260 27396 204312 27402
rect 204260 27338 204312 27344
rect 201592 25764 201644 25770
rect 201592 25706 201644 25712
rect 201500 4208 201552 4214
rect 201500 4150 201552 4156
rect 201604 3482 201632 25706
rect 204272 16574 204300 27338
rect 205652 16574 205680 33866
rect 204272 16546 205128 16574
rect 205652 16546 206232 16574
rect 203892 6860 203944 6866
rect 203892 6802 203944 6808
rect 202696 4208 202748 4214
rect 202696 4150 202748 4156
rect 201512 3454 201632 3482
rect 201512 480 201540 3454
rect 202708 480 202736 4150
rect 203904 480 203932 6802
rect 205100 480 205128 16546
rect 206204 480 206232 16546
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 60114
rect 208400 27328 208452 27334
rect 208400 27270 208452 27276
rect 208412 16574 208440 27270
rect 208412 16546 208624 16574
rect 208596 480 208624 16546
rect 209792 480 209820 73714
rect 209872 69624 209924 69630
rect 209872 69566 209924 69572
rect 209884 16574 209912 69566
rect 212538 17640 212594 17649
rect 212538 17575 212594 17584
rect 212552 16574 212580 17575
rect 213932 16574 213960 78882
rect 226340 77240 226392 77246
rect 226340 77182 226392 77188
rect 223580 74520 223632 74526
rect 223580 74462 223632 74468
rect 214104 73704 214156 73710
rect 214104 73646 214156 73652
rect 214116 70990 214144 73646
rect 215300 71732 215352 71738
rect 215300 71674 215352 71680
rect 214104 70984 214156 70990
rect 214104 70926 214156 70932
rect 215312 69018 215340 71674
rect 215300 69012 215352 69018
rect 215300 68954 215352 68960
rect 218152 69012 218204 69018
rect 218152 68954 218204 68960
rect 218164 65822 218192 68954
rect 220820 66972 220872 66978
rect 220820 66914 220872 66920
rect 218060 65816 218112 65822
rect 218060 65758 218112 65764
rect 218152 65816 218204 65822
rect 218152 65758 218204 65764
rect 215300 27260 215352 27266
rect 215300 27202 215352 27208
rect 209884 16546 211016 16574
rect 212552 16546 213408 16574
rect 213932 16546 214512 16574
rect 210988 480 211016 16546
rect 213092 5092 213144 5098
rect 213092 5034 213144 5040
rect 213104 3874 213132 5034
rect 212172 3868 212224 3874
rect 212172 3810 212224 3816
rect 213092 3868 213144 3874
rect 213092 3810 213144 3816
rect 212184 480 212212 3810
rect 213380 480 213408 16546
rect 214484 480 214512 16546
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 27202
rect 216864 5024 216916 5030
rect 216864 4966 216916 4972
rect 216876 480 216904 4966
rect 218072 480 218100 65758
rect 219440 33856 219492 33862
rect 219440 33798 219492 33804
rect 218152 27192 218204 27198
rect 218152 27134 218204 27140
rect 218164 16574 218192 27134
rect 219452 16574 219480 33798
rect 220832 16574 220860 66914
rect 218164 16546 219296 16574
rect 219452 16546 220032 16574
rect 220832 16546 221136 16574
rect 219268 480 219296 16546
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 16546
rect 222752 7948 222804 7954
rect 222752 7890 222804 7896
rect 222764 480 222792 7890
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 74462
rect 226248 65816 226300 65822
rect 226248 65758 226300 65764
rect 224960 63096 225012 63102
rect 224960 63038 225012 63044
rect 224972 16574 225000 63038
rect 226260 60178 226288 65758
rect 226248 60172 226300 60178
rect 226248 60114 226300 60120
rect 224972 16546 225184 16574
rect 225156 480 225184 16546
rect 226352 480 226380 77182
rect 229192 75812 229244 75818
rect 229192 75754 229244 75760
rect 229204 74186 229232 75754
rect 230478 74352 230534 74361
rect 230478 74287 230534 74296
rect 229100 74180 229152 74186
rect 229100 74122 229152 74128
rect 229192 74180 229244 74186
rect 229192 74122 229244 74128
rect 229112 71738 229140 74122
rect 229100 71732 229152 71738
rect 229100 71674 229152 71680
rect 226430 33960 226486 33969
rect 226430 33895 226486 33904
rect 226444 16574 226472 33895
rect 230492 16574 230520 74287
rect 226444 16546 227576 16574
rect 230492 16546 231072 16574
rect 227548 480 227576 16546
rect 229374 13424 229430 13433
rect 229374 13359 229430 13368
rect 228730 6080 228786 6089
rect 228730 6015 228786 6024
rect 228744 480 228772 6015
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229388 354 229416 13359
rect 231044 480 231072 16546
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 80174
rect 252560 80164 252612 80170
rect 252560 80106 252612 80112
rect 249800 79144 249852 79150
rect 249800 79086 249852 79092
rect 242164 77648 242216 77654
rect 242164 77590 242216 77596
rect 240140 77172 240192 77178
rect 240140 77114 240192 77120
rect 238760 65748 238812 65754
rect 238760 65690 238812 65696
rect 233240 60104 233292 60110
rect 233240 60046 233292 60052
rect 233252 16574 233280 60046
rect 236000 27124 236052 27130
rect 236000 27066 236052 27072
rect 234620 18896 234672 18902
rect 234620 18838 234672 18844
rect 233252 16546 233464 16574
rect 233436 480 233464 16546
rect 234632 480 234660 18838
rect 236012 16574 236040 27066
rect 238772 16574 238800 65690
rect 236012 16546 236592 16574
rect 238772 16546 239352 16574
rect 235816 6792 235868 6798
rect 235816 6734 235868 6740
rect 235828 480 235856 6734
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 237656 16176 237708 16182
rect 237656 16118 237708 16124
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 16118
rect 239324 480 239352 16546
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240152 354 240180 77114
rect 242176 20194 242204 77590
rect 247038 76800 247094 76809
rect 247038 76735 247094 76744
rect 243728 75880 243780 75886
rect 243728 75822 243780 75828
rect 243740 74526 243768 75822
rect 243728 74520 243780 74526
rect 243728 74462 243780 74468
rect 244278 74216 244334 74225
rect 244278 74151 244334 74160
rect 242900 28620 242952 28626
rect 242900 28562 242952 28568
rect 241520 20188 241572 20194
rect 241520 20130 241572 20136
rect 242164 20188 242216 20194
rect 242164 20130 242216 20136
rect 241532 16574 241560 20130
rect 241532 16546 241744 16574
rect 241716 480 241744 16546
rect 242912 4214 242940 28562
rect 244292 16574 244320 74151
rect 245658 58576 245714 58585
rect 245658 58511 245714 58520
rect 245672 16574 245700 58511
rect 247052 16574 247080 76735
rect 247684 60172 247736 60178
rect 247684 60114 247736 60120
rect 247696 50386 247724 60114
rect 247684 50380 247736 50386
rect 247684 50322 247736 50328
rect 248418 20088 248474 20097
rect 248418 20023 248474 20032
rect 244292 16546 245240 16574
rect 245672 16546 245976 16574
rect 247052 16546 247632 16574
rect 242992 7880 243044 7886
rect 242992 7822 243044 7828
rect 242900 4208 242952 4214
rect 242900 4150 242952 4156
rect 243004 3482 243032 7822
rect 244096 4208 244148 4214
rect 244096 4150 244148 4156
rect 242912 3454 243032 3482
rect 242912 480 242940 3454
rect 244108 480 244136 4150
rect 245212 480 245240 16546
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 16546
rect 247604 480 247632 16546
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248432 354 248460 20023
rect 249812 16574 249840 79086
rect 251180 74452 251232 74458
rect 251180 74394 251232 74400
rect 250444 70372 250496 70378
rect 250444 70314 250496 70320
rect 250456 54398 250484 70314
rect 250444 54392 250496 54398
rect 250444 54334 250496 54340
rect 249812 16546 250024 16574
rect 249996 480 250024 16546
rect 251192 4214 251220 74394
rect 251272 28552 251324 28558
rect 251272 28494 251324 28500
rect 251180 4208 251232 4214
rect 251180 4150 251232 4156
rect 251284 3482 251312 28494
rect 252572 16574 252600 80106
rect 266372 78878 266400 697546
rect 299492 144226 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 299480 144220 299532 144226
rect 299480 144162 299532 144168
rect 267832 79008 267884 79014
rect 267832 78950 267884 78956
rect 266360 78872 266412 78878
rect 266360 78814 266412 78820
rect 255964 78532 256016 78538
rect 255964 78474 256016 78480
rect 255320 71596 255372 71602
rect 255320 71538 255372 71544
rect 255332 69018 255360 71538
rect 255320 69012 255372 69018
rect 255320 68954 255372 68960
rect 253020 54392 253072 54398
rect 253020 54334 253072 54340
rect 253032 51066 253060 54334
rect 253020 51060 253072 51066
rect 253020 51002 253072 51008
rect 253940 28484 253992 28490
rect 253940 28426 253992 28432
rect 253952 16574 253980 28426
rect 255976 20262 256004 78474
rect 260840 77104 260892 77110
rect 260840 77046 260892 77052
rect 258080 75744 258132 75750
rect 258080 75686 258132 75692
rect 258092 72894 258120 75686
rect 259460 75676 259512 75682
rect 259460 75618 259512 75624
rect 258080 72888 258132 72894
rect 258080 72830 258132 72836
rect 259472 72826 259500 75618
rect 259460 72820 259512 72826
rect 259460 72762 259512 72768
rect 258724 71732 258776 71738
rect 258724 71674 258776 71680
rect 257344 70984 257396 70990
rect 257344 70926 257396 70932
rect 256700 66904 256752 66910
rect 256700 66846 256752 66852
rect 255320 20256 255372 20262
rect 255320 20198 255372 20204
rect 255964 20256 256016 20262
rect 255964 20198 256016 20204
rect 255332 16574 255360 20198
rect 252572 16546 253520 16574
rect 253952 16546 254256 16574
rect 255332 16546 255912 16574
rect 252376 4208 252428 4214
rect 252376 4150 252428 4156
rect 251192 3454 251312 3482
rect 251192 480 251220 3454
rect 252388 480 252416 4150
rect 253492 480 253520 16546
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 255884 480 255912 16546
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 256712 354 256740 66846
rect 257356 61674 257384 70926
rect 257344 61668 257396 61674
rect 257344 61610 257396 61616
rect 258736 59362 258764 71674
rect 258816 69012 258868 69018
rect 258816 68954 258868 68960
rect 258828 59974 258856 68954
rect 258816 59968 258868 59974
rect 258816 59910 258868 59916
rect 258724 59356 258776 59362
rect 258724 59298 258776 59304
rect 258724 51060 258776 51066
rect 258724 51002 258776 51008
rect 258736 39370 258764 51002
rect 258724 39364 258776 39370
rect 258724 39306 258776 39312
rect 259460 33788 259512 33794
rect 259460 33730 259512 33736
rect 258080 28416 258132 28422
rect 258080 28358 258132 28364
rect 258092 16574 258120 28358
rect 258092 16546 258304 16574
rect 258276 480 258304 16546
rect 259472 480 259500 33730
rect 260852 16574 260880 77046
rect 264244 71528 264296 71534
rect 264244 71470 264296 71476
rect 264256 64462 264284 71470
rect 264244 64456 264296 64462
rect 264244 64398 264296 64404
rect 263598 62792 263654 62801
rect 263598 62727 263654 62736
rect 262864 61668 262916 61674
rect 262864 61610 262916 61616
rect 261484 59356 261536 59362
rect 261484 59298 261536 59304
rect 261496 56574 261524 59298
rect 261484 56568 261536 56574
rect 261484 56510 261536 56516
rect 262876 54466 262904 61610
rect 262864 54460 262916 54466
rect 262864 54402 262916 54408
rect 262220 20324 262272 20330
rect 262220 20266 262272 20272
rect 262232 16574 262260 20266
rect 263612 16574 263640 62727
rect 264336 59968 264388 59974
rect 264336 59910 264388 59916
rect 264244 56568 264296 56574
rect 264244 56510 264296 56516
rect 264256 46850 264284 56510
rect 264348 53106 264376 59910
rect 264336 53100 264388 53106
rect 264336 53042 264388 53048
rect 264244 46844 264296 46850
rect 264244 46786 264296 46792
rect 267004 46844 267056 46850
rect 267004 46786 267056 46792
rect 266358 33824 266414 33833
rect 266358 33759 266414 33768
rect 266372 16574 266400 33759
rect 267016 32706 267044 46786
rect 267004 32700 267056 32706
rect 267004 32642 267056 32648
rect 260852 16546 261800 16574
rect 262232 16546 262536 16574
rect 263612 16546 264192 16574
rect 266372 16546 266584 16574
rect 260656 7812 260708 7818
rect 260656 7754 260708 7760
rect 260668 480 260696 7754
rect 261772 480 261800 16546
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 264164 480 264192 16546
rect 265346 9616 265402 9625
rect 265346 9551 265402 9560
rect 265360 480 265388 9551
rect 266556 480 266584 16546
rect 267844 6914 267872 78950
rect 315304 78464 315356 78470
rect 315304 78406 315356 78412
rect 296720 77036 296772 77042
rect 296720 76978 296772 76984
rect 282918 76664 282974 76673
rect 282918 76599 282974 76608
rect 270040 74384 270092 74390
rect 270040 74326 270092 74332
rect 268200 72888 268252 72894
rect 268200 72830 268252 72836
rect 268212 66230 268240 72830
rect 270052 67590 270080 74326
rect 275376 72820 275428 72826
rect 275376 72762 275428 72768
rect 271880 71460 271932 71466
rect 271880 71402 271932 71408
rect 271788 70304 271840 70310
rect 271788 70246 271840 70252
rect 270040 67584 270092 67590
rect 270040 67526 270092 67532
rect 271800 66502 271828 70246
rect 271892 68202 271920 71402
rect 271880 68196 271932 68202
rect 271880 68138 271932 68144
rect 275284 68196 275336 68202
rect 275284 68138 275336 68144
rect 275192 67584 275244 67590
rect 275192 67526 275244 67532
rect 271788 66496 271840 66502
rect 271788 66438 271840 66444
rect 268200 66224 268252 66230
rect 268200 66166 268252 66172
rect 271144 66224 271196 66230
rect 271144 66166 271196 66172
rect 269764 64456 269816 64462
rect 269764 64398 269816 64404
rect 269776 50998 269804 64398
rect 269856 54460 269908 54466
rect 269856 54402 269908 54408
rect 269764 50992 269816 50998
rect 269764 50934 269816 50940
rect 269868 42974 269896 54402
rect 271156 49706 271184 66166
rect 274640 63028 274692 63034
rect 274640 62970 274692 62976
rect 273168 50992 273220 50998
rect 273168 50934 273220 50940
rect 271144 49700 271196 49706
rect 271144 49642 271196 49648
rect 273180 46306 273208 50934
rect 273168 46300 273220 46306
rect 273168 46242 273220 46248
rect 269856 42968 269908 42974
rect 269856 42910 269908 42916
rect 274652 16574 274680 62970
rect 275204 61674 275232 67526
rect 275192 61668 275244 61674
rect 275192 61610 275244 61616
rect 275296 58682 275324 68138
rect 275388 63782 275416 72762
rect 280068 72752 280120 72758
rect 280068 72694 280120 72700
rect 278780 66496 278832 66502
rect 278780 66438 278832 66444
rect 275376 63776 275428 63782
rect 275376 63718 275428 63724
rect 278412 63776 278464 63782
rect 278412 63718 278464 63724
rect 275284 58676 275336 58682
rect 275284 58618 275336 58624
rect 278424 56574 278452 63718
rect 278792 63646 278820 66438
rect 280080 65754 280108 72694
rect 280068 65748 280120 65754
rect 280068 65690 280120 65696
rect 278780 63640 278832 63646
rect 278780 63582 278832 63588
rect 278412 56568 278464 56574
rect 278412 56510 278464 56516
rect 280804 56568 280856 56574
rect 280804 56510 280856 56516
rect 274732 50380 274784 50386
rect 274732 50322 274784 50328
rect 274744 46578 274772 50322
rect 277492 49700 277544 49706
rect 277492 49642 277544 49648
rect 274732 46572 274784 46578
rect 274732 46514 274784 46520
rect 277504 46238 277532 49642
rect 279424 46572 279476 46578
rect 279424 46514 279476 46520
rect 277492 46232 277544 46238
rect 277492 46174 277544 46180
rect 276020 42968 276072 42974
rect 276020 42910 276072 42916
rect 276032 39438 276060 42910
rect 276020 39432 276072 39438
rect 276020 39374 276072 39380
rect 278044 39364 278096 39370
rect 278044 39306 278096 39312
rect 278056 34610 278084 39306
rect 278044 34604 278096 34610
rect 278044 34546 278096 34552
rect 275284 32700 275336 32706
rect 275284 32642 275336 32648
rect 275296 18902 275324 32642
rect 279436 30326 279464 46514
rect 280816 42294 280844 56510
rect 281356 53100 281408 53106
rect 281356 53042 281408 53048
rect 281368 45626 281396 53042
rect 282184 46300 282236 46306
rect 282184 46242 282236 46248
rect 281356 45620 281408 45626
rect 281356 45562 281408 45568
rect 280804 42288 280856 42294
rect 280804 42230 280856 42236
rect 282196 37942 282224 46242
rect 282184 37936 282236 37942
rect 282184 37878 282236 37884
rect 279424 30320 279476 30326
rect 279424 30262 279476 30268
rect 275284 18896 275336 18902
rect 275284 18838 275336 18844
rect 282932 16574 282960 76599
rect 288532 75608 288584 75614
rect 288532 75550 288584 75556
rect 288440 75540 288492 75546
rect 288440 75482 288492 75488
rect 288452 72214 288480 75482
rect 288440 72208 288492 72214
rect 288440 72150 288492 72156
rect 286324 71664 286376 71670
rect 286324 71606 286376 71612
rect 283012 63640 283064 63646
rect 283012 63582 283064 63588
rect 283024 58750 283052 63582
rect 286336 58818 286364 71606
rect 287612 71392 287664 71398
rect 287612 71334 287664 71340
rect 287624 66230 287652 71334
rect 288544 69018 288572 75550
rect 296074 72584 296130 72593
rect 296074 72519 296130 72528
rect 288532 69012 288584 69018
rect 288532 68954 288584 68960
rect 295340 69012 295392 69018
rect 295340 68954 295392 68960
rect 287612 66224 287664 66230
rect 287612 66166 287664 66172
rect 291108 66224 291160 66230
rect 291108 66166 291160 66172
rect 286324 58812 286376 58818
rect 286324 58754 286376 58760
rect 283012 58744 283064 58750
rect 283012 58686 283064 58692
rect 291120 58682 291148 66166
rect 295352 65754 295380 68954
rect 292856 65748 292908 65754
rect 292856 65690 292908 65696
rect 295340 65748 295392 65754
rect 295340 65690 295392 65696
rect 292580 61600 292632 61606
rect 292580 61542 292632 61548
rect 291844 58744 291896 58750
rect 291844 58686 291896 58692
rect 283656 58676 283708 58682
rect 283656 58618 283708 58624
rect 291108 58676 291160 58682
rect 291108 58618 291160 58624
rect 283668 54534 283696 58618
rect 291856 54670 291884 58686
rect 291844 54664 291896 54670
rect 291844 54606 291896 54612
rect 283656 54528 283708 54534
rect 283656 54470 283708 54476
rect 288440 46232 288492 46238
rect 288440 46174 288492 46180
rect 287704 45620 287756 45626
rect 287704 45562 287756 45568
rect 284300 42288 284352 42294
rect 284300 42230 284352 42236
rect 284312 37534 284340 42230
rect 284944 39432 284996 39438
rect 284944 39374 284996 39380
rect 284300 37528 284352 37534
rect 284300 37470 284352 37476
rect 284956 23254 284984 39374
rect 287428 37528 287480 37534
rect 287428 37470 287480 37476
rect 287440 35358 287468 37470
rect 287060 35352 287112 35358
rect 287060 35294 287112 35300
rect 287428 35352 287480 35358
rect 287428 35294 287480 35300
rect 285680 34604 285732 34610
rect 285680 34546 285732 34552
rect 285692 32706 285720 34546
rect 285680 32700 285732 32706
rect 285680 32642 285732 32648
rect 286324 30320 286376 30326
rect 286324 30262 286376 30268
rect 285680 29912 285732 29918
rect 285680 29854 285732 29860
rect 284944 23248 284996 23254
rect 284944 23190 284996 23196
rect 285692 16574 285720 29854
rect 286336 24750 286364 30262
rect 286324 24744 286376 24750
rect 286324 24686 286376 24692
rect 287072 16574 287100 35294
rect 287716 28966 287744 45562
rect 288452 40050 288480 46174
rect 288440 40044 288492 40050
rect 288440 39986 288492 39992
rect 291844 40044 291896 40050
rect 291844 39986 291896 39992
rect 291200 35284 291252 35290
rect 291200 35226 291252 35232
rect 287704 28960 287756 28966
rect 287704 28902 287756 28908
rect 291108 28960 291160 28966
rect 291108 28902 291160 28908
rect 291120 25770 291148 28902
rect 291108 25764 291160 25770
rect 291108 25706 291160 25712
rect 289820 24676 289872 24682
rect 289820 24618 289872 24624
rect 288440 18896 288492 18902
rect 288440 18838 288492 18844
rect 274652 16546 274864 16574
rect 282932 16546 283144 16574
rect 285692 16546 286640 16574
rect 287072 16546 287376 16574
rect 267752 6886 267872 6914
rect 267752 480 267780 6886
rect 271236 6724 271288 6730
rect 271236 6666 271288 6672
rect 270040 6656 270092 6662
rect 270040 6598 270092 6604
rect 268844 4072 268896 4078
rect 268844 4014 268896 4020
rect 268856 480 268884 4014
rect 270052 480 270080 6598
rect 271248 480 271276 6666
rect 273628 6588 273680 6594
rect 273628 6530 273680 6536
rect 272432 4004 272484 4010
rect 272432 3946 272484 3952
rect 272444 480 272472 3946
rect 273640 480 273668 6530
rect 274836 480 274864 16546
rect 281906 9480 281962 9489
rect 281906 9415 281962 9424
rect 278320 7744 278372 7750
rect 278320 7686 278372 7692
rect 276020 6520 276072 6526
rect 276020 6462 276072 6468
rect 276032 480 276060 6462
rect 277124 6452 277176 6458
rect 277124 6394 277176 6400
rect 277136 480 277164 6394
rect 278332 480 278360 7686
rect 280710 6896 280766 6905
rect 280710 6831 280766 6840
rect 279516 6384 279568 6390
rect 279516 6326 279568 6332
rect 279528 480 279556 6326
rect 280724 480 280752 6831
rect 281920 480 281948 9415
rect 283116 480 283144 16546
rect 284298 6760 284354 6769
rect 284298 6695 284354 6704
rect 284312 480 284340 6695
rect 285404 3392 285456 3398
rect 285404 3334 285456 3340
rect 285416 480 285444 3334
rect 286612 480 286640 16546
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 288452 16182 288480 18838
rect 288440 16176 288492 16182
rect 288440 16118 288492 16124
rect 288992 4140 289044 4146
rect 288992 4082 289044 4088
rect 289004 480 289032 4082
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 289832 354 289860 24618
rect 291212 16574 291240 35226
rect 291856 31210 291884 39986
rect 291844 31204 291896 31210
rect 291844 31146 291896 31152
rect 291212 16546 291424 16574
rect 291396 480 291424 16546
rect 292592 480 292620 61542
rect 292868 60994 292896 65690
rect 292856 60988 292908 60994
rect 292856 60930 292908 60936
rect 295984 60988 296036 60994
rect 295984 60930 296036 60936
rect 295340 54664 295392 54670
rect 295340 54606 295392 54612
rect 292672 54528 292724 54534
rect 292672 54470 292724 54476
rect 292684 46238 292712 54470
rect 295352 51746 295380 54606
rect 295340 51740 295392 51746
rect 295340 51682 295392 51688
rect 292672 46232 292724 46238
rect 292672 46174 292724 46180
rect 293960 32700 294012 32706
rect 293960 32642 294012 32648
rect 293972 29986 294000 32642
rect 293960 29980 294012 29986
rect 293960 29922 294012 29928
rect 295996 27130 296024 60930
rect 296088 57254 296116 72519
rect 296168 72208 296220 72214
rect 296168 72150 296220 72156
rect 296180 58750 296208 72150
rect 296168 58744 296220 58750
rect 296168 58686 296220 58692
rect 296076 57248 296128 57254
rect 296076 57190 296128 57196
rect 295984 27124 296036 27130
rect 295984 27066 296036 27072
rect 292672 25696 292724 25702
rect 292672 25638 292724 25644
rect 292684 16574 292712 25638
rect 292764 24744 292816 24750
rect 292764 24686 292816 24692
rect 292776 18902 292804 24686
rect 292764 18896 292816 18902
rect 292764 18838 292816 18844
rect 296732 16574 296760 76978
rect 301136 74248 301188 74254
rect 301136 74190 301188 74196
rect 298098 72448 298154 72457
rect 298098 72383 298154 72392
rect 297364 61668 297416 61674
rect 297364 61610 297416 61616
rect 297376 54534 297404 61610
rect 297364 54528 297416 54534
rect 297364 54470 297416 54476
rect 292684 16546 293264 16574
rect 296732 16546 297312 16574
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 296076 9648 296128 9654
rect 296076 9590 296128 9596
rect 294880 4956 294932 4962
rect 294880 4898 294932 4904
rect 294892 480 294920 4898
rect 296088 480 296116 9590
rect 297284 480 297312 16546
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 354 298140 72383
rect 301148 71398 301176 74190
rect 307760 72684 307812 72690
rect 307760 72626 307812 72632
rect 301136 71392 301188 71398
rect 301136 71334 301188 71340
rect 306930 71088 306986 71097
rect 306930 71023 306986 71032
rect 306944 67590 306972 71023
rect 306932 67584 306984 67590
rect 306932 67526 306984 67532
rect 303620 65748 303672 65754
rect 303620 65690 303672 65696
rect 303632 59362 303660 65690
rect 306380 61532 306432 61538
rect 306380 61474 306432 61480
rect 305000 60036 305052 60042
rect 305000 59978 305052 59984
rect 303620 59356 303672 59362
rect 303620 59298 303672 59304
rect 298744 58812 298796 58818
rect 298744 58754 298796 58760
rect 298284 37936 298336 37942
rect 298284 37878 298336 37884
rect 298296 30054 298324 37878
rect 298284 30048 298336 30054
rect 298284 29990 298336 29996
rect 298756 29918 298784 58754
rect 301596 57248 301648 57254
rect 301596 57190 301648 57196
rect 301608 46850 301636 57190
rect 301596 46844 301648 46850
rect 301596 46786 301648 46792
rect 304264 46844 304316 46850
rect 304264 46786 304316 46792
rect 301504 46232 301556 46238
rect 301504 46174 301556 46180
rect 299204 35352 299256 35358
rect 299204 35294 299256 35300
rect 299216 31142 299244 35294
rect 299204 31136 299256 31142
rect 299204 31078 299256 31084
rect 298744 29912 298796 29918
rect 298744 29854 298796 29860
rect 301516 24886 301544 46174
rect 301596 31204 301648 31210
rect 301596 31146 301648 31152
rect 301504 24880 301556 24886
rect 301504 24822 301556 24828
rect 299296 23248 299348 23254
rect 299296 23190 299348 23196
rect 299308 20398 299336 23190
rect 301608 21826 301636 31146
rect 304276 28422 304304 46786
rect 304264 28416 304316 28422
rect 304264 28358 304316 28364
rect 302884 27124 302936 27130
rect 302884 27066 302936 27072
rect 302240 25764 302292 25770
rect 302240 25706 302292 25712
rect 302252 23322 302280 25706
rect 302240 23316 302292 23322
rect 302240 23258 302292 23264
rect 301596 21820 301648 21826
rect 301596 21762 301648 21768
rect 299296 20392 299348 20398
rect 299296 20334 299348 20340
rect 302056 18896 302108 18902
rect 302056 18838 302108 18844
rect 300858 17504 300914 17513
rect 300858 17439 300914 17448
rect 300872 16574 300900 17439
rect 300872 16546 301544 16574
rect 298744 16176 298796 16182
rect 298744 16118 298796 16124
rect 298756 6390 298784 16118
rect 299662 9344 299718 9353
rect 299662 9279 299718 9288
rect 298744 6384 298796 6390
rect 298744 6326 298796 6332
rect 299676 480 299704 9279
rect 300766 6624 300822 6633
rect 300766 6559 300822 6568
rect 300780 480 300808 6559
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 16546
rect 302068 15298 302096 18838
rect 302896 16182 302924 27066
rect 303620 27056 303672 27062
rect 303620 26998 303672 27004
rect 303632 16574 303660 26998
rect 304264 21820 304316 21826
rect 304264 21762 304316 21768
rect 304276 16574 304304 21762
rect 305012 16574 305040 59978
rect 305644 24880 305696 24886
rect 305644 24822 305696 24828
rect 303632 16546 303936 16574
rect 304276 16546 304396 16574
rect 305012 16546 305592 16574
rect 302884 16176 302936 16182
rect 302884 16118 302936 16124
rect 302056 15292 302108 15298
rect 302056 15234 302108 15240
rect 303160 3936 303212 3942
rect 303160 3878 303212 3884
rect 303172 480 303200 3878
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 304264 15292 304316 15298
rect 304264 15234 304316 15240
rect 304276 13802 304304 15234
rect 304264 13796 304316 13802
rect 304264 13738 304316 13744
rect 304368 12374 304396 16546
rect 304356 12368 304408 12374
rect 304356 12310 304408 12316
rect 305564 480 305592 16546
rect 305656 14890 305684 24822
rect 305644 14884 305696 14890
rect 305644 14826 305696 14832
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306392 354 306420 61474
rect 307024 59356 307076 59362
rect 307024 59298 307076 59304
rect 307036 49706 307064 59298
rect 307024 49700 307076 49706
rect 307024 49642 307076 49648
rect 307024 13796 307076 13802
rect 307024 13738 307076 13744
rect 307036 6458 307064 13738
rect 307024 6452 307076 6458
rect 307024 6394 307076 6400
rect 307772 3398 307800 72626
rect 311900 72616 311952 72622
rect 311900 72558 311952 72564
rect 311164 71392 311216 71398
rect 311164 71334 311216 71340
rect 309784 67584 309836 67590
rect 309784 67526 309836 67532
rect 309796 57254 309824 67526
rect 311176 65754 311204 71334
rect 311164 65748 311216 65754
rect 311164 65690 311216 65696
rect 311164 58676 311216 58682
rect 311164 58618 311216 58624
rect 309784 57248 309836 57254
rect 309784 57190 309836 57196
rect 311176 53106 311204 58618
rect 311164 53100 311216 53106
rect 311164 53042 311216 53048
rect 311164 30048 311216 30054
rect 311164 29990 311216 29996
rect 311176 23254 311204 29990
rect 311164 23248 311216 23254
rect 311164 23190 311216 23196
rect 311912 16574 311940 72558
rect 313924 58744 313976 58750
rect 313924 58686 313976 58692
rect 313936 53514 313964 58686
rect 313924 53508 313976 53514
rect 313924 53450 313976 53456
rect 311992 49700 312044 49706
rect 311992 49642 312044 49648
rect 312004 46102 312032 49642
rect 311992 46096 312044 46102
rect 311992 46038 312044 46044
rect 313280 31136 313332 31142
rect 313280 31078 313332 31084
rect 313292 27062 313320 31078
rect 313280 27056 313332 27062
rect 313280 26998 313332 27004
rect 313280 23316 313332 23322
rect 313280 23258 313332 23264
rect 313292 20330 313320 23258
rect 313280 20324 313332 20330
rect 313280 20266 313332 20272
rect 311912 16546 312216 16574
rect 309600 14884 309652 14890
rect 309600 14826 309652 14832
rect 309612 9654 309640 14826
rect 311440 14816 311492 14822
rect 311440 14758 311492 14764
rect 309784 10464 309836 10470
rect 309784 10406 309836 10412
rect 309600 9648 309652 9654
rect 309600 9590 309652 9596
rect 307944 7676 307996 7682
rect 307944 7618 307996 7624
rect 307760 3392 307812 3398
rect 307760 3334 307812 3340
rect 307956 480 307984 7618
rect 309048 3392 309100 3398
rect 309048 3334 309100 3340
rect 309060 480 309088 3334
rect 306718 354 306830 480
rect 306392 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 10406
rect 311452 480 311480 14758
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312188 354 312216 16546
rect 313924 16176 313976 16182
rect 313924 16118 313976 16124
rect 312544 12368 312596 12374
rect 312544 12310 312596 12316
rect 312556 3942 312584 12310
rect 313832 10396 313884 10402
rect 313832 10338 313884 10344
rect 313096 9648 313148 9654
rect 313096 9590 313148 9596
rect 313108 5574 313136 9590
rect 313096 5568 313148 5574
rect 313096 5510 313148 5516
rect 312544 3936 312596 3942
rect 312544 3878 312596 3884
rect 313844 480 313872 10338
rect 313936 6526 313964 16118
rect 315316 9654 315344 78406
rect 331232 77926 331260 702986
rect 348804 700534 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 348792 700528 348844 700534
rect 348792 700470 348844 700476
rect 364352 140146 364380 702406
rect 364340 140140 364392 140146
rect 364340 140082 364392 140088
rect 397472 78810 397500 703520
rect 413664 700466 413692 703520
rect 413652 700460 413704 700466
rect 413652 700402 413704 700408
rect 429212 142866 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 429200 142860 429252 142866
rect 429200 142802 429252 142808
rect 430580 80096 430632 80102
rect 430580 80038 430632 80044
rect 397460 78804 397512 78810
rect 397460 78746 397512 78752
rect 426440 78736 426492 78742
rect 426440 78678 426492 78684
rect 331220 77920 331272 77926
rect 331220 77862 331272 77868
rect 331128 76968 331180 76974
rect 331128 76910 331180 76916
rect 322940 74316 322992 74322
rect 322940 74258 322992 74264
rect 318800 74112 318852 74118
rect 318800 74054 318852 74060
rect 316684 71324 316736 71330
rect 316684 71266 316736 71272
rect 316040 65748 316092 65754
rect 316040 65690 316092 65696
rect 316052 62626 316080 65690
rect 316040 62620 316092 62626
rect 316040 62562 316092 62568
rect 316696 41886 316724 71266
rect 316776 53508 316828 53514
rect 316776 53450 316828 53456
rect 316788 42838 316816 53450
rect 318156 53100 318208 53106
rect 318156 53042 318208 53048
rect 318064 51740 318116 51746
rect 318064 51682 318116 51688
rect 317420 46096 317472 46102
rect 317420 46038 317472 46044
rect 317432 43450 317460 46038
rect 317420 43444 317472 43450
rect 317420 43386 317472 43392
rect 316776 42832 316828 42838
rect 316776 42774 316828 42780
rect 316684 41880 316736 41886
rect 316684 41822 316736 41828
rect 318076 31550 318104 51682
rect 318168 44742 318196 53042
rect 318156 44736 318208 44742
rect 318156 44678 318208 44684
rect 318064 31544 318116 31550
rect 318064 31486 318116 31492
rect 317418 29880 317474 29889
rect 317418 29815 317474 29824
rect 317432 16574 317460 29815
rect 318812 16574 318840 74054
rect 322952 71330 322980 74258
rect 324320 74044 324372 74050
rect 324320 73986 324372 73992
rect 324332 71398 324360 73986
rect 324320 71392 324372 71398
rect 324320 71334 324372 71340
rect 330484 71392 330536 71398
rect 330484 71334 330536 71340
rect 322940 71324 322992 71330
rect 322940 71266 322992 71272
rect 327724 70236 327776 70242
rect 327724 70178 327776 70184
rect 326988 70168 327040 70174
rect 326988 70110 327040 70116
rect 327000 67522 327028 70110
rect 326988 67516 327040 67522
rect 326988 67458 327040 67464
rect 318984 62620 319036 62626
rect 318984 62562 319036 62568
rect 318996 60450 319024 62562
rect 318984 60444 319036 60450
rect 318984 60386 319036 60392
rect 323584 57248 323636 57254
rect 323584 57190 323636 57196
rect 319444 42832 319496 42838
rect 319444 42774 319496 42780
rect 319456 23458 319484 42774
rect 319812 41880 319864 41886
rect 319812 41822 319864 41828
rect 319824 37262 319852 41822
rect 323596 40050 323624 57190
rect 326344 54528 326396 54534
rect 326344 54470 326396 54476
rect 324320 44736 324372 44742
rect 324320 44678 324372 44684
rect 324332 40730 324360 44678
rect 324320 40724 324372 40730
rect 324320 40666 324372 40672
rect 323584 40044 323636 40050
rect 323584 39986 323636 39992
rect 326356 39370 326384 54470
rect 327736 45150 327764 70178
rect 327816 70100 327868 70106
rect 327816 70042 327868 70048
rect 327828 60654 327856 70042
rect 329104 67516 329156 67522
rect 329104 67458 329156 67464
rect 327816 60648 327868 60654
rect 327816 60590 327868 60596
rect 327908 60444 327960 60450
rect 327908 60386 327960 60392
rect 327920 52426 327948 60386
rect 329116 56574 329144 67458
rect 330496 65754 330524 71334
rect 331140 69018 331168 76910
rect 346400 76900 346452 76906
rect 346400 76842 346452 76848
rect 339130 75576 339186 75585
rect 339130 75511 339186 75520
rect 331864 73976 331916 73982
rect 331864 73918 331916 73924
rect 331128 69012 331180 69018
rect 331128 68954 331180 68960
rect 330484 65748 330536 65754
rect 330484 65690 330536 65696
rect 329104 56568 329156 56574
rect 329104 56510 329156 56516
rect 327908 52420 327960 52426
rect 327908 52362 327960 52368
rect 331876 50386 331904 73918
rect 339144 73302 339172 75511
rect 340144 75472 340196 75478
rect 340144 75414 340196 75420
rect 339132 73296 339184 73302
rect 339132 73238 339184 73244
rect 332600 71324 332652 71330
rect 332600 71266 332652 71272
rect 332612 68610 332640 71266
rect 339408 71256 339460 71262
rect 339408 71198 339460 71204
rect 338764 70032 338816 70038
rect 338764 69974 338816 69980
rect 336004 69012 336056 69018
rect 336004 68954 336056 68960
rect 332600 68604 332652 68610
rect 332600 68546 332652 68552
rect 332600 60648 332652 60654
rect 332600 60590 332652 60596
rect 332612 56642 332640 60590
rect 336016 58682 336044 68954
rect 338120 64320 338172 64326
rect 338120 64262 338172 64268
rect 336004 58676 336056 58682
rect 336004 58618 336056 58624
rect 332600 56636 332652 56642
rect 332600 56578 332652 56584
rect 336004 56636 336056 56642
rect 336004 56578 336056 56584
rect 333980 56568 334032 56574
rect 333980 56510 334032 56516
rect 333992 53106 334020 56510
rect 333980 53100 334032 53106
rect 333980 53042 334032 53048
rect 332600 52420 332652 52426
rect 332600 52362 332652 52368
rect 331864 50380 331916 50386
rect 331864 50322 331916 50328
rect 332612 49706 332640 52362
rect 332600 49700 332652 49706
rect 332600 49642 332652 49648
rect 327724 45144 327776 45150
rect 327724 45086 327776 45092
rect 332600 45144 332652 45150
rect 332600 45086 332652 45092
rect 330484 40724 330536 40730
rect 330484 40666 330536 40672
rect 326436 40044 326488 40050
rect 326436 39986 326488 39992
rect 326344 39364 326396 39370
rect 326344 39306 326396 39312
rect 319812 37256 319864 37262
rect 319812 37198 319864 37204
rect 322848 37256 322900 37262
rect 322848 37198 322900 37204
rect 322860 33794 322888 37198
rect 322848 33788 322900 33794
rect 322848 33730 322900 33736
rect 322940 31544 322992 31550
rect 322940 31486 322992 31492
rect 320824 29980 320876 29986
rect 320824 29922 320876 29928
rect 320836 24070 320864 29922
rect 321744 27056 321796 27062
rect 321744 26998 321796 27004
rect 320824 24064 320876 24070
rect 320824 24006 320876 24012
rect 319444 23452 319496 23458
rect 319444 23394 319496 23400
rect 321756 22166 321784 26998
rect 321744 22160 321796 22166
rect 321744 22102 321796 22108
rect 322204 20324 322256 20330
rect 322204 20266 322256 20272
rect 317432 16546 318104 16574
rect 318812 16546 319760 16574
rect 316038 10432 316094 10441
rect 316038 10367 316094 10376
rect 315304 9648 315356 9654
rect 315304 9590 315356 9596
rect 315026 9208 315082 9217
rect 315026 9143 315082 9152
rect 313924 6520 313976 6526
rect 313924 6462 313976 6468
rect 314660 5568 314712 5574
rect 314660 5510 314712 5516
rect 314672 4010 314700 5510
rect 314660 4004 314712 4010
rect 314660 3946 314712 3952
rect 315040 480 315068 9143
rect 316052 3398 316080 10367
rect 316222 7576 316278 7585
rect 316222 7511 316278 7520
rect 316040 3392 316092 3398
rect 316040 3334 316092 3340
rect 316236 480 316264 7511
rect 317328 3392 317380 3398
rect 317328 3334 317380 3340
rect 317340 480 317368 3334
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 319732 480 319760 16546
rect 322216 8362 322244 20266
rect 322204 8356 322256 8362
rect 322204 8298 322256 8304
rect 322756 6520 322808 6526
rect 322756 6462 322808 6468
rect 320916 6384 320968 6390
rect 320916 6326 320968 6332
rect 320928 480 320956 6326
rect 322112 3936 322164 3942
rect 322112 3878 322164 3884
rect 322124 480 322152 3878
rect 322768 3330 322796 6462
rect 322756 3324 322808 3330
rect 322756 3266 322808 3272
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 322952 354 322980 31486
rect 326448 31278 326476 39986
rect 329104 33788 329156 33794
rect 329104 33730 329156 33736
rect 326436 31272 326488 31278
rect 326436 31214 326488 31220
rect 326436 29912 326488 29918
rect 326436 29854 326488 29860
rect 323492 28416 323544 28422
rect 323492 28358 323544 28364
rect 323504 20330 323532 28358
rect 326344 23452 326396 23458
rect 326344 23394 326396 23400
rect 323584 23248 323636 23254
rect 323584 23190 323636 23196
rect 323492 20324 323544 20330
rect 323492 20266 323544 20272
rect 323596 12442 323624 23190
rect 324320 22160 324372 22166
rect 324320 22102 324372 22108
rect 324332 17066 324360 22102
rect 324320 17060 324372 17066
rect 324320 17002 324372 17008
rect 323584 12436 323636 12442
rect 323584 12378 323636 12384
rect 326252 12436 326304 12442
rect 326252 12378 326304 12384
rect 326264 6914 326292 12378
rect 326356 11778 326384 23394
rect 326448 12374 326476 29854
rect 327724 24064 327776 24070
rect 327724 24006 327776 24012
rect 326528 20392 326580 20398
rect 326528 20334 326580 20340
rect 326540 16182 326568 20334
rect 327080 17060 327132 17066
rect 327080 17002 327132 17008
rect 327092 16574 327120 17002
rect 327092 16546 327396 16574
rect 326528 16176 326580 16182
rect 326528 16118 326580 16124
rect 326436 12368 326488 12374
rect 326436 12310 326488 12316
rect 326356 11750 326476 11778
rect 326264 6886 326384 6914
rect 324412 4004 324464 4010
rect 324412 3946 324464 3952
rect 324424 480 324452 3946
rect 325608 3324 325660 3330
rect 325608 3266 325660 3272
rect 325620 480 325648 3266
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 6886
rect 326448 3126 326476 11750
rect 327080 8356 327132 8362
rect 327080 8298 327132 8304
rect 326436 3120 326488 3126
rect 326436 3062 326488 3068
rect 327092 2990 327120 8298
rect 327368 6914 327396 16546
rect 327736 8906 327764 24006
rect 329116 21826 329144 33730
rect 330496 27606 330524 40666
rect 332612 39438 332640 45086
rect 336016 44198 336044 56578
rect 337384 49700 337436 49706
rect 337384 49642 337436 49648
rect 336004 44192 336056 44198
rect 336004 44134 336056 44140
rect 332600 39432 332652 39438
rect 332600 39374 332652 39380
rect 331220 31272 331272 31278
rect 331220 31214 331272 31220
rect 330484 27600 330536 27606
rect 330484 27542 330536 27548
rect 331232 26518 331260 31214
rect 337396 31210 337424 49642
rect 337936 39364 337988 39370
rect 337936 39306 337988 39312
rect 337948 37262 337976 39306
rect 337936 37256 337988 37262
rect 337936 37198 337988 37204
rect 337384 31204 337436 31210
rect 337384 31146 337436 31152
rect 332600 29844 332652 29850
rect 332600 29786 332652 29792
rect 331220 26512 331272 26518
rect 331220 26454 331272 26460
rect 329104 21820 329156 21826
rect 329104 21762 329156 21768
rect 327724 8900 327776 8906
rect 327724 8842 327776 8848
rect 330392 8900 330444 8906
rect 330392 8842 330444 8848
rect 327368 6886 328040 6914
rect 327080 2984 327132 2990
rect 327080 2926 327132 2932
rect 328012 480 328040 6886
rect 329196 6452 329248 6458
rect 329196 6394 329248 6400
rect 329208 480 329236 6394
rect 330404 480 330432 8842
rect 332612 3210 332640 29786
rect 334256 27600 334308 27606
rect 334256 27542 334308 27548
rect 334268 24682 334296 27542
rect 335360 26512 335412 26518
rect 335360 26454 335412 26460
rect 334256 24676 334308 24682
rect 334256 24618 334308 24624
rect 335372 16574 335400 26454
rect 338132 16574 338160 64262
rect 338776 60790 338804 69974
rect 339420 66774 339448 71198
rect 339408 66768 339460 66774
rect 339408 66710 339460 66716
rect 338764 60784 338816 60790
rect 338764 60726 338816 60732
rect 340156 54534 340184 75414
rect 341064 73296 341116 73302
rect 341064 73238 341116 73244
rect 340880 72548 340932 72554
rect 340880 72490 340932 72496
rect 340788 65748 340840 65754
rect 340788 65690 340840 65696
rect 340800 61606 340828 65690
rect 340788 61600 340840 61606
rect 340788 61542 340840 61548
rect 340144 54528 340196 54534
rect 340144 54470 340196 54476
rect 340144 53100 340196 53106
rect 340144 53042 340196 53048
rect 339960 50380 340012 50386
rect 339960 50322 340012 50328
rect 339972 46238 340000 50322
rect 339960 46232 340012 46238
rect 339960 46174 340012 46180
rect 340156 44878 340184 53042
rect 340144 44872 340196 44878
rect 340144 44814 340196 44820
rect 339408 44192 339460 44198
rect 339408 44134 339460 44140
rect 339420 40730 339448 44134
rect 339408 40724 339460 40730
rect 339408 40666 339460 40672
rect 340144 39432 340196 39438
rect 340144 39374 340196 39380
rect 340156 36650 340184 39374
rect 340144 36644 340196 36650
rect 340144 36586 340196 36592
rect 339500 29776 339552 29782
rect 339500 29718 339552 29724
rect 335372 16546 336320 16574
rect 338132 16546 338712 16574
rect 332692 12368 332744 12374
rect 332692 12310 332744 12316
rect 332704 3398 332732 12310
rect 332692 3392 332744 3398
rect 332692 3334 332744 3340
rect 333888 3392 333940 3398
rect 333888 3334 333940 3340
rect 332612 3182 332732 3210
rect 331588 3120 331640 3126
rect 331588 3062 331640 3068
rect 331600 480 331628 3062
rect 332704 480 332732 3182
rect 333900 480 333928 3334
rect 335084 2984 335136 2990
rect 335084 2926 335136 2932
rect 335096 480 335124 2926
rect 336292 480 336320 16546
rect 337016 16176 337068 16182
rect 337016 16118 337068 16124
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337028 354 337056 16118
rect 338684 480 338712 16546
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339512 354 339540 29718
rect 340892 3210 340920 72490
rect 341076 68678 341104 73238
rect 346412 69018 346440 76842
rect 374000 76832 374052 76838
rect 374000 76774 374052 76780
rect 369122 75440 369178 75449
rect 359372 75404 359424 75410
rect 369122 75375 369178 75384
rect 359372 75346 359424 75352
rect 347504 74520 347556 74526
rect 347504 74462 347556 74468
rect 346400 69012 346452 69018
rect 346400 68954 346452 68960
rect 341064 68672 341116 68678
rect 341064 68614 341116 68620
rect 347228 68604 347280 68610
rect 347228 68546 347280 68552
rect 345664 66768 345716 66774
rect 345664 66710 345716 66716
rect 340972 62960 341024 62966
rect 340972 62902 341024 62908
rect 340984 3398 341012 62902
rect 344284 60784 344336 60790
rect 344284 60726 344336 60732
rect 343640 54528 343692 54534
rect 343640 54470 343692 54476
rect 343652 50386 343680 54470
rect 343640 50380 343692 50386
rect 343640 50322 343692 50328
rect 344296 47326 344324 60726
rect 344284 47320 344336 47326
rect 344284 47262 344336 47268
rect 344284 43444 344336 43450
rect 344284 43386 344336 43392
rect 341064 40724 341116 40730
rect 341064 40666 341116 40672
rect 341076 37194 341104 40666
rect 342904 37256 342956 37262
rect 342904 37198 342956 37204
rect 341064 37188 341116 37194
rect 341064 37130 341116 37136
rect 342916 31142 342944 37198
rect 344296 33998 344324 43386
rect 345676 39370 345704 66710
rect 347240 61538 347268 68546
rect 347516 66230 347544 74462
rect 349802 74080 349858 74089
rect 349802 74015 349858 74024
rect 349816 71738 349844 74015
rect 354680 72480 354732 72486
rect 354680 72422 354732 72428
rect 349804 71732 349856 71738
rect 349804 71674 349856 71680
rect 349804 69012 349856 69018
rect 349804 68954 349856 68960
rect 347504 66224 347556 66230
rect 347504 66166 347556 66172
rect 347228 61532 347280 61538
rect 347228 61474 347280 61480
rect 349816 48278 349844 68954
rect 352564 68672 352616 68678
rect 352564 68614 352616 68620
rect 349988 66224 350040 66230
rect 349988 66166 350040 66172
rect 350000 62014 350028 66166
rect 352576 64054 352604 68614
rect 353298 68232 353354 68241
rect 353298 68167 353354 68176
rect 352564 64048 352616 64054
rect 352564 63990 352616 63996
rect 349988 62008 350040 62014
rect 349988 61950 350040 61956
rect 351918 51776 351974 51785
rect 351918 51711 351974 51720
rect 349804 48272 349856 48278
rect 349804 48214 349856 48220
rect 346400 47320 346452 47326
rect 346400 47262 346452 47268
rect 346412 44946 346440 47262
rect 349804 46232 349856 46238
rect 349804 46174 349856 46180
rect 346400 44940 346452 44946
rect 346400 44882 346452 44888
rect 345664 39364 345716 39370
rect 345664 39306 345716 39312
rect 344376 37188 344428 37194
rect 344376 37130 344428 37136
rect 344284 33992 344336 33998
rect 344284 33934 344336 33940
rect 342904 31136 342956 31142
rect 342904 31078 342956 31084
rect 344388 28490 344416 37130
rect 347596 33992 347648 33998
rect 347596 33934 347648 33940
rect 347044 31204 347096 31210
rect 347044 31146 347096 31152
rect 346400 29708 346452 29714
rect 346400 29650 346452 29656
rect 344376 28484 344428 28490
rect 344376 28426 344428 28432
rect 342260 24676 342312 24682
rect 342260 24618 342312 24624
rect 342272 17270 342300 24618
rect 344284 21820 344336 21826
rect 344284 21762 344336 21768
rect 343640 21752 343692 21758
rect 343640 21694 343692 21700
rect 342260 17264 342312 17270
rect 342260 17206 342312 17212
rect 342904 16108 342956 16114
rect 342904 16050 342956 16056
rect 340972 3392 341024 3398
rect 340972 3334 341024 3340
rect 342168 3392 342220 3398
rect 342168 3334 342220 3340
rect 340892 3182 341012 3210
rect 340984 480 341012 3182
rect 342180 480 342208 3334
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 16050
rect 343652 6914 343680 21694
rect 344296 16114 344324 21762
rect 346412 16574 346440 29650
rect 347056 18902 347084 31146
rect 347608 28422 347636 33934
rect 349816 31754 349844 46174
rect 349804 31748 349856 31754
rect 349804 31690 349856 31696
rect 349158 29744 349214 29753
rect 349158 29679 349214 29688
rect 348884 28484 348936 28490
rect 348884 28426 348936 28432
rect 347596 28416 347648 28422
rect 347596 28358 347648 28364
rect 348896 25294 348924 28426
rect 348884 25288 348936 25294
rect 348884 25230 348936 25236
rect 347044 18896 347096 18902
rect 347044 18838 347096 18844
rect 348700 17264 348752 17270
rect 348700 17206 348752 17212
rect 346412 16546 346992 16574
rect 344284 16108 344336 16114
rect 344284 16050 344336 16056
rect 345296 12300 345348 12306
rect 345296 12242 345348 12248
rect 343652 6886 344600 6914
rect 344572 480 344600 6886
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 12242
rect 346964 480 346992 16546
rect 348712 12442 348740 17206
rect 348700 12436 348752 12442
rect 348700 12378 348752 12384
rect 348056 6316 348108 6322
rect 348056 6258 348108 6264
rect 348068 480 348096 6258
rect 349172 1290 349200 29679
rect 351828 25288 351880 25294
rect 351828 25230 351880 25236
rect 351840 18086 351868 25230
rect 351828 18080 351880 18086
rect 351828 18022 351880 18028
rect 351932 16574 351960 51711
rect 352012 48272 352064 48278
rect 352012 48214 352064 48220
rect 352024 42770 352052 48214
rect 352104 44872 352156 44878
rect 352104 44814 352156 44820
rect 352012 42764 352064 42770
rect 352012 42706 352064 42712
rect 352116 40730 352144 44814
rect 352104 40724 352156 40730
rect 352104 40666 352156 40672
rect 353312 16574 353340 68167
rect 353944 62008 353996 62014
rect 353944 61950 353996 61956
rect 353956 51066 353984 61950
rect 354036 61600 354088 61606
rect 354036 61542 354088 61548
rect 354048 53174 354076 61542
rect 354036 53168 354088 53174
rect 354036 53110 354088 53116
rect 353944 51060 353996 51066
rect 353944 51002 353996 51008
rect 353392 31748 353444 31754
rect 353392 31690 353444 31696
rect 353404 27742 353432 31690
rect 353484 31136 353536 31142
rect 353484 31078 353536 31084
rect 353392 27736 353444 27742
rect 353392 27678 353444 27684
rect 353496 26314 353524 31078
rect 353484 26308 353536 26314
rect 353484 26250 353536 26256
rect 351932 16546 352880 16574
rect 353312 16546 353616 16574
rect 349252 12232 349304 12238
rect 349252 12174 349304 12180
rect 349160 1284 349212 1290
rect 349160 1226 349212 1232
rect 349264 480 349292 12174
rect 351642 6488 351698 6497
rect 351642 6423 351698 6432
rect 350448 1284 350500 1290
rect 350448 1226 350500 1232
rect 350460 480 350488 1226
rect 351656 480 351684 6423
rect 352852 480 352880 16546
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 353588 354 353616 16546
rect 354692 6914 354720 72422
rect 359384 71738 359412 75346
rect 362960 73908 363012 73914
rect 362960 73850 363012 73856
rect 355508 71732 355560 71738
rect 355508 71674 355560 71680
rect 359372 71732 359424 71738
rect 359372 71674 359424 71680
rect 355520 68678 355548 71674
rect 362972 71262 363000 73850
rect 368480 73840 368532 73846
rect 368480 73782 368532 73788
rect 365076 71732 365128 71738
rect 365076 71674 365128 71680
rect 362960 71256 363012 71262
rect 362960 71198 363012 71204
rect 361580 69964 361632 69970
rect 361580 69906 361632 69912
rect 355508 68672 355560 68678
rect 355508 68614 355560 68620
rect 359280 68672 359332 68678
rect 359280 68614 359332 68620
rect 358820 68536 358872 68542
rect 358820 68478 358872 68484
rect 357348 64048 357400 64054
rect 357348 63990 357400 63996
rect 357360 59362 357388 63990
rect 357348 59356 357400 59362
rect 357348 59298 357400 59304
rect 356244 53168 356296 53174
rect 356244 53110 356296 53116
rect 356256 47666 356284 53110
rect 356704 51060 356756 51066
rect 356704 51002 356756 51008
rect 356244 47660 356296 47666
rect 356244 47602 356296 47608
rect 355324 42764 355376 42770
rect 355324 42706 355376 42712
rect 355336 37262 355364 42706
rect 355324 37256 355376 37262
rect 355324 37198 355376 37204
rect 356716 35358 356744 51002
rect 356704 35352 356756 35358
rect 356704 35294 356756 35300
rect 357440 35216 357492 35222
rect 357440 35158 357492 35164
rect 356704 28416 356756 28422
rect 356704 28358 356756 28364
rect 356060 27736 356112 27742
rect 356060 27678 356112 27684
rect 356072 24682 356100 27678
rect 356152 26308 356204 26314
rect 356152 26250 356204 26256
rect 356060 24676 356112 24682
rect 356060 24618 356112 24624
rect 356164 23254 356192 26250
rect 356152 23248 356204 23254
rect 356152 23190 356204 23196
rect 356716 19310 356744 28358
rect 356704 19304 356756 19310
rect 356704 19246 356756 19252
rect 354772 18080 354824 18086
rect 354772 18022 354824 18028
rect 354784 12238 354812 18022
rect 357348 16108 357400 16114
rect 357348 16050 357400 16056
rect 357072 12436 357124 12442
rect 357072 12378 357124 12384
rect 354772 12232 354824 12238
rect 354772 12174 354824 12180
rect 357084 8906 357112 12378
rect 357360 12306 357388 16050
rect 357348 12300 357400 12306
rect 357348 12242 357400 12248
rect 357072 8900 357124 8906
rect 357072 8842 357124 8848
rect 354692 6886 355272 6914
rect 355244 480 355272 6886
rect 356336 3800 356388 3806
rect 356336 3742 356388 3748
rect 356348 480 356376 3742
rect 357452 2514 357480 35158
rect 358084 20324 358136 20330
rect 358084 20266 358136 20272
rect 358096 16114 358124 20266
rect 358832 16574 358860 68478
rect 359292 65754 359320 68614
rect 359280 65748 359332 65754
rect 359280 65690 359332 65696
rect 361592 64938 361620 69906
rect 365088 68270 365116 71674
rect 365076 68264 365128 68270
rect 365076 68206 365128 68212
rect 361580 64932 361632 64938
rect 361580 64874 361632 64880
rect 364984 64932 365036 64938
rect 364984 64874 365036 64880
rect 363604 61532 363656 61538
rect 363604 61474 363656 61480
rect 362960 61464 363012 61470
rect 362960 61406 363012 61412
rect 362224 58676 362276 58682
rect 362224 58618 362276 58624
rect 362236 52426 362264 58618
rect 362224 52420 362276 52426
rect 362224 52362 362276 52368
rect 359464 50380 359516 50386
rect 359464 50322 359516 50328
rect 359476 18970 359504 50322
rect 359556 44940 359608 44946
rect 359556 44882 359608 44888
rect 359568 27606 359596 44882
rect 362224 39364 362276 39370
rect 362224 39306 362276 39312
rect 360844 37256 360896 37262
rect 360844 37198 360896 37204
rect 360856 28830 360884 37198
rect 362132 36644 362184 36650
rect 362132 36586 362184 36592
rect 361580 35352 361632 35358
rect 361580 35294 361632 35300
rect 361592 33046 361620 35294
rect 361580 33040 361632 33046
rect 361580 32982 361632 32988
rect 362144 32706 362172 36586
rect 362132 32700 362184 32706
rect 362132 32642 362184 32648
rect 360844 28824 360896 28830
rect 360844 28766 360896 28772
rect 359556 27600 359608 27606
rect 359556 27542 359608 27548
rect 362236 20670 362264 39306
rect 362224 20664 362276 20670
rect 362224 20606 362276 20612
rect 359556 19304 359608 19310
rect 359556 19246 359608 19252
rect 359464 18964 359516 18970
rect 359464 18906 359516 18912
rect 358832 16546 359504 16574
rect 358084 16108 358136 16114
rect 358084 16050 358136 16056
rect 357532 13184 357584 13190
rect 357532 13126 357584 13132
rect 357440 2508 357492 2514
rect 357440 2450 357492 2456
rect 357544 480 357572 13126
rect 358728 2508 358780 2514
rect 358728 2450 358780 2456
rect 358740 480 358768 2450
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 16546
rect 359568 3806 359596 19246
rect 362972 16574 363000 61406
rect 363616 53786 363644 61474
rect 363696 59356 363748 59362
rect 363696 59298 363748 59304
rect 363604 53780 363656 53786
rect 363604 53722 363656 53728
rect 363708 53310 363736 59298
rect 364996 54534 365024 64874
rect 364984 54528 365036 54534
rect 364984 54470 365036 54476
rect 366548 53780 366600 53786
rect 366548 53722 366600 53728
rect 363696 53304 363748 53310
rect 363696 53246 363748 53252
rect 365628 52420 365680 52426
rect 365628 52362 365680 52368
rect 365640 48278 365668 52362
rect 366560 49842 366588 53722
rect 367008 53304 367060 53310
rect 367008 53246 367060 53252
rect 366548 49836 366600 49842
rect 366548 49778 366600 49784
rect 365628 48272 365680 48278
rect 365628 48214 365680 48220
rect 367020 48210 367048 53246
rect 367008 48204 367060 48210
rect 367008 48146 367060 48152
rect 364984 33040 365036 33046
rect 364984 32982 365036 32988
rect 363328 27600 363380 27606
rect 363328 27542 363380 27548
rect 363340 24750 363368 27542
rect 363328 24744 363380 24750
rect 363328 24686 363380 24692
rect 362972 16546 363552 16574
rect 361120 16040 361172 16046
rect 361120 15982 361172 15988
rect 359556 3800 359608 3806
rect 359556 3742 359608 3748
rect 361132 480 361160 15982
rect 362316 8900 362368 8906
rect 362316 8842 362368 8848
rect 362328 480 362356 8842
rect 363524 480 363552 16546
rect 364996 11694 365024 32982
rect 365168 28824 365220 28830
rect 365168 28766 365220 28772
rect 365076 20664 365128 20670
rect 365076 20606 365128 20612
rect 364984 11688 365036 11694
rect 364984 11630 365036 11636
rect 365088 7682 365116 20606
rect 365180 17950 365208 28766
rect 365168 17944 365220 17950
rect 365168 17886 365220 17892
rect 368492 16574 368520 73782
rect 369136 73710 369164 75375
rect 369124 73704 369176 73710
rect 369124 73646 369176 73652
rect 370504 71256 370556 71262
rect 370504 71198 370556 71204
rect 369124 68264 369176 68270
rect 369124 68206 369176 68212
rect 369136 56574 369164 68206
rect 369124 56568 369176 56574
rect 369124 56510 369176 56516
rect 370516 55894 370544 71198
rect 370964 65748 371016 65754
rect 370964 65690 371016 65696
rect 370976 61810 371004 65690
rect 370964 61804 371016 61810
rect 370964 61746 371016 61752
rect 371884 56568 371936 56574
rect 371884 56510 371936 56516
rect 370504 55888 370556 55894
rect 370504 55830 370556 55836
rect 370504 48272 370556 48278
rect 370504 48214 370556 48220
rect 370516 32774 370544 48214
rect 371240 48204 371292 48210
rect 371240 48146 371292 48152
rect 371252 43178 371280 48146
rect 371240 43172 371292 43178
rect 371240 43114 371292 43120
rect 370504 32768 370556 32774
rect 370504 32710 370556 32716
rect 371896 31142 371924 56510
rect 373264 49836 373316 49842
rect 373264 49778 373316 49784
rect 372618 35184 372674 35193
rect 372618 35119 372674 35128
rect 371884 31136 371936 31142
rect 371884 31078 371936 31084
rect 369124 24744 369176 24750
rect 369124 24686 369176 24692
rect 369136 19038 369164 24686
rect 369860 24676 369912 24682
rect 369860 24618 369912 24624
rect 369872 20330 369900 24618
rect 369952 23248 370004 23254
rect 369952 23190 370004 23196
rect 369860 20324 369912 20330
rect 369860 20266 369912 20272
rect 369124 19032 369176 19038
rect 369124 18974 369176 18980
rect 369964 17406 369992 23190
rect 369952 17400 370004 17406
rect 369952 17342 370004 17348
rect 372632 16574 372660 35119
rect 368492 16546 369440 16574
rect 372632 16546 372936 16574
rect 365718 15872 365774 15881
rect 365718 15807 365774 15816
rect 365076 7676 365128 7682
rect 365076 7618 365128 7624
rect 364616 3868 364668 3874
rect 364616 3810 364668 3816
rect 364628 480 364656 3810
rect 365732 3210 365760 15807
rect 365812 13116 365864 13122
rect 365812 13058 365864 13064
rect 365824 3398 365852 13058
rect 367744 11688 367796 11694
rect 367744 11630 367796 11636
rect 367756 3874 367784 11630
rect 367744 3868 367796 3874
rect 367744 3810 367796 3816
rect 368204 3800 368256 3806
rect 368204 3742 368256 3748
rect 365812 3392 365864 3398
rect 365812 3334 365864 3340
rect 367008 3392 367060 3398
rect 367008 3334 367060 3340
rect 365732 3182 365852 3210
rect 365824 480 365852 3182
rect 367020 480 367048 3334
rect 368216 480 368244 3742
rect 369412 480 369440 16546
rect 370134 13288 370190 13297
rect 370134 13223 370190 13232
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370148 354 370176 13223
rect 371238 13152 371294 13161
rect 371238 13087 371294 13096
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 371252 354 371280 13087
rect 372908 480 372936 16546
rect 373276 7750 373304 49778
rect 373448 17944 373500 17950
rect 373448 17886 373500 17892
rect 373460 12306 373488 17886
rect 373356 12300 373408 12306
rect 373356 12242 373408 12248
rect 373448 12300 373500 12306
rect 373448 12242 373500 12248
rect 373264 7744 373316 7750
rect 373264 7686 373316 7692
rect 373368 6322 373396 12242
rect 373356 6316 373408 6322
rect 373356 6258 373408 6264
rect 374012 1170 374040 76774
rect 408500 76764 408552 76770
rect 408500 76706 408552 76712
rect 382924 74180 382976 74186
rect 382924 74122 382976 74128
rect 378414 73944 378470 73953
rect 378414 73879 378470 73888
rect 374736 73704 374788 73710
rect 374736 73646 374788 73652
rect 374092 64252 374144 64258
rect 374092 64194 374144 64200
rect 374104 3398 374132 64194
rect 374644 54528 374696 54534
rect 374644 54470 374696 54476
rect 374184 47660 374236 47666
rect 374184 47602 374236 47608
rect 374196 44674 374224 47602
rect 374184 44668 374236 44674
rect 374184 44610 374236 44616
rect 374656 31822 374684 54470
rect 374748 54398 374776 73646
rect 378428 71806 378456 73879
rect 378416 71800 378468 71806
rect 378416 71742 378468 71748
rect 376668 61804 376720 61810
rect 376668 61746 376720 61752
rect 376680 57254 376708 61746
rect 376668 57248 376720 57254
rect 376668 57190 376720 57196
rect 374736 54392 374788 54398
rect 374736 54334 374788 54340
rect 380164 54392 380216 54398
rect 380164 54334 380216 54340
rect 376024 43172 376076 43178
rect 376024 43114 376076 43120
rect 375288 40724 375340 40730
rect 375288 40666 375340 40672
rect 375300 37942 375328 40666
rect 375288 37936 375340 37942
rect 375288 37878 375340 37884
rect 376036 33862 376064 43114
rect 380176 37330 380204 54334
rect 380164 37324 380216 37330
rect 380164 37266 380216 37272
rect 382936 35970 382964 74122
rect 384764 71800 384816 71806
rect 384764 71742 384816 71748
rect 384776 67590 384804 71742
rect 384764 67584 384816 67590
rect 384764 67526 384816 67532
rect 387064 67584 387116 67590
rect 387064 67526 387116 67532
rect 384396 57248 384448 57254
rect 384396 57190 384448 57196
rect 383016 44668 383068 44674
rect 383016 44610 383068 44616
rect 382924 35964 382976 35970
rect 382924 35906 382976 35912
rect 376024 33856 376076 33862
rect 376024 33798 376076 33804
rect 383028 33794 383056 44610
rect 384304 37324 384356 37330
rect 384304 37266 384356 37272
rect 383016 33788 383068 33794
rect 383016 33730 383068 33736
rect 378140 32768 378192 32774
rect 378140 32710 378192 32716
rect 374736 32700 374788 32706
rect 374736 32642 374788 32648
rect 374644 31816 374696 31822
rect 374644 31758 374696 31764
rect 374748 25702 374776 32642
rect 377404 31816 377456 31822
rect 377404 31758 377456 31764
rect 374736 25696 374788 25702
rect 374736 25638 374788 25644
rect 377416 24886 377444 31758
rect 378152 28966 378180 32710
rect 378784 31136 378836 31142
rect 378784 31078 378836 31084
rect 378140 28960 378192 28966
rect 378140 28902 378192 28908
rect 378796 27742 378824 31078
rect 381544 28960 381596 28966
rect 381544 28902 381596 28908
rect 378784 27736 378836 27742
rect 378784 27678 378836 27684
rect 377404 24880 377456 24886
rect 377404 24822 377456 24828
rect 380164 24880 380216 24886
rect 380164 24822 380216 24828
rect 379520 20324 379572 20330
rect 379520 20266 379572 20272
rect 378692 19032 378744 19038
rect 378692 18974 378744 18980
rect 377404 18964 377456 18970
rect 377404 18906 377456 18912
rect 375380 17400 375432 17406
rect 375380 17342 375432 17348
rect 375392 13122 375420 17342
rect 377416 13870 377444 18906
rect 377404 13864 377456 13870
rect 377404 13806 377456 13812
rect 375380 13116 375432 13122
rect 375380 13058 375432 13064
rect 376024 12232 376076 12238
rect 376024 12174 376076 12180
rect 376036 5574 376064 12174
rect 378704 11694 378732 18974
rect 379532 17950 379560 20266
rect 379520 17944 379572 17950
rect 379520 17886 379572 17892
rect 380176 15230 380204 24822
rect 380164 15224 380216 15230
rect 380164 15166 380216 15172
rect 380900 13864 380952 13870
rect 380900 13806 380952 13812
rect 379520 12300 379572 12306
rect 379520 12242 379572 12248
rect 378692 11688 378744 11694
rect 378692 11630 378744 11636
rect 376484 7676 376536 7682
rect 376484 7618 376536 7624
rect 376024 5568 376076 5574
rect 376024 5510 376076 5516
rect 374092 3392 374144 3398
rect 374092 3334 374144 3340
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 374012 1142 374132 1170
rect 374104 480 374132 1142
rect 375300 480 375328 3334
rect 376496 480 376524 7618
rect 378048 6316 378100 6322
rect 378048 6258 378100 6264
rect 377680 3868 377732 3874
rect 377680 3810 377732 3816
rect 377692 480 377720 3810
rect 378060 3058 378088 6258
rect 378876 5568 378928 5574
rect 378876 5510 378928 5516
rect 378048 3052 378100 3058
rect 378048 2994 378100 3000
rect 378888 480 378916 5510
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 370566 -960 370678 326
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379532 354 379560 12242
rect 380912 7682 380940 13806
rect 381268 11688 381320 11694
rect 381268 11630 381320 11636
rect 381176 7744 381228 7750
rect 381176 7686 381228 7692
rect 380900 7676 380952 7682
rect 380900 7618 380952 7624
rect 381188 480 381216 7686
rect 381280 6934 381308 11630
rect 381556 7750 381584 28902
rect 381636 25696 381688 25702
rect 381636 25638 381688 25644
rect 381648 12442 381676 25638
rect 382280 17944 382332 17950
rect 382280 17886 382332 17892
rect 382292 14754 382320 17886
rect 382924 15224 382976 15230
rect 382924 15166 382976 15172
rect 382372 14816 382424 14822
rect 382372 14758 382424 14764
rect 382280 14748 382332 14754
rect 382280 14690 382332 14696
rect 381728 13116 381780 13122
rect 381728 13058 381780 13064
rect 381636 12436 381688 12442
rect 381636 12378 381688 12384
rect 381544 7744 381596 7750
rect 381544 7686 381596 7692
rect 381268 6928 381320 6934
rect 381268 6870 381320 6876
rect 381740 6322 381768 13058
rect 381728 6316 381780 6322
rect 381728 6258 381780 6264
rect 382384 3398 382412 14758
rect 382936 3806 382964 15166
rect 384316 5574 384344 37266
rect 384408 32842 384436 57190
rect 385684 35964 385736 35970
rect 385684 35906 385736 35912
rect 384488 33856 384540 33862
rect 384488 33798 384540 33804
rect 384396 32836 384448 32842
rect 384396 32778 384448 32784
rect 384500 24682 384528 33798
rect 385040 27736 385092 27742
rect 385040 27678 385092 27684
rect 384488 24676 384540 24682
rect 384488 24618 384540 24624
rect 384396 12436 384448 12442
rect 384396 12378 384448 12384
rect 384304 5568 384356 5574
rect 384304 5510 384356 5516
rect 382924 3800 382976 3806
rect 382924 3742 382976 3748
rect 382372 3392 382424 3398
rect 382372 3334 382424 3340
rect 383568 3392 383620 3398
rect 383568 3334 383620 3340
rect 382372 3052 382424 3058
rect 382372 2994 382424 3000
rect 382384 480 382412 2994
rect 383580 480 383608 3334
rect 384408 3194 384436 12378
rect 384764 6928 384816 6934
rect 385052 6914 385080 27678
rect 385696 16046 385724 35906
rect 387076 30326 387104 67526
rect 387708 55888 387760 55894
rect 387708 55830 387760 55836
rect 387720 51270 387748 55830
rect 387708 51264 387760 51270
rect 387708 51206 387760 51212
rect 391204 51264 391256 51270
rect 391204 51206 391256 51212
rect 388444 37936 388496 37942
rect 388444 37878 388496 37884
rect 387064 30320 387116 30326
rect 387064 30262 387116 30268
rect 385868 16108 385920 16114
rect 385868 16050 385920 16056
rect 385684 16040 385736 16046
rect 385684 15982 385736 15988
rect 385880 13802 385908 16050
rect 385868 13796 385920 13802
rect 385868 13738 385920 13744
rect 385052 6886 386000 6914
rect 384764 6870 384816 6876
rect 384396 3188 384448 3194
rect 384396 3130 384448 3136
rect 384776 480 384804 6870
rect 385972 480 386000 6886
rect 387156 5568 387208 5574
rect 387156 5510 387208 5516
rect 387168 480 387196 5510
rect 388456 3874 388484 37878
rect 391216 23458 391244 51206
rect 396724 33788 396776 33794
rect 396724 33730 396776 33736
rect 391940 32836 391992 32842
rect 391940 32778 391992 32784
rect 391952 29714 391980 32778
rect 392584 30320 392636 30326
rect 392584 30262 392636 30268
rect 391940 29708 391992 29714
rect 391940 29650 391992 29656
rect 391204 23452 391256 23458
rect 391204 23394 391256 23400
rect 388536 18896 388588 18902
rect 388536 18838 388588 18844
rect 388444 3868 388496 3874
rect 388444 3810 388496 3816
rect 388548 3806 388576 18838
rect 392596 17270 392624 30262
rect 393320 23452 393372 23458
rect 393320 23394 393372 23400
rect 392584 17264 392636 17270
rect 392584 17206 392636 17212
rect 393332 16574 393360 23394
rect 396736 20670 396764 33730
rect 397552 29708 397604 29714
rect 397552 29650 397604 29656
rect 397460 28348 397512 28354
rect 397460 28290 397512 28296
rect 396724 20664 396776 20670
rect 396724 20606 396776 20612
rect 397184 17264 397236 17270
rect 397184 17206 397236 17212
rect 393332 16546 394280 16574
rect 390560 16040 390612 16046
rect 390560 15982 390612 15988
rect 390572 12442 390600 15982
rect 392584 13796 392636 13802
rect 392584 13738 392636 13744
rect 390560 12436 390612 12442
rect 390560 12378 390612 12384
rect 390652 12164 390704 12170
rect 390652 12106 390704 12112
rect 388260 3800 388312 3806
rect 388260 3742 388312 3748
rect 388536 3800 388588 3806
rect 388536 3742 388588 3748
rect 388272 480 388300 3742
rect 389456 3188 389508 3194
rect 389456 3130 389508 3136
rect 389468 480 389496 3130
rect 390664 480 390692 12106
rect 391848 7744 391900 7750
rect 391848 7686 391900 7692
rect 391860 480 391888 7686
rect 392596 6390 392624 13738
rect 393044 7676 393096 7682
rect 393044 7618 393096 7624
rect 392584 6384 392636 6390
rect 392584 6326 392636 6332
rect 393056 480 393084 7618
rect 394252 480 394280 16546
rect 397196 12442 397224 17206
rect 397472 16574 397500 28290
rect 397564 27606 397592 29650
rect 397552 27600 397604 27606
rect 397552 27542 397604 27548
rect 400864 27600 400916 27606
rect 400864 27542 400916 27548
rect 398932 20664 398984 20670
rect 398932 20606 398984 20612
rect 397472 16546 397776 16574
rect 395344 12436 395396 12442
rect 395344 12378 395396 12384
rect 397184 12436 397236 12442
rect 397184 12378 397236 12384
rect 395252 6316 395304 6322
rect 395252 6258 395304 6264
rect 395264 3074 395292 6258
rect 395356 3262 395384 12378
rect 396540 3868 396592 3874
rect 396540 3810 396592 3816
rect 395344 3256 395396 3262
rect 395344 3198 395396 3204
rect 395264 3046 395384 3074
rect 395356 480 395384 3046
rect 396552 480 396580 3810
rect 397748 480 397776 16546
rect 398104 6384 398156 6390
rect 398104 6326 398156 6332
rect 398116 3874 398144 6326
rect 398104 3868 398156 3874
rect 398104 3810 398156 3816
rect 398840 3800 398892 3806
rect 398840 3742 398892 3748
rect 398852 1986 398880 3742
rect 398944 3398 398972 20606
rect 400876 18018 400904 27542
rect 407212 24676 407264 24682
rect 407212 24618 407264 24624
rect 404360 23180 404412 23186
rect 404360 23122 404412 23128
rect 400864 18012 400916 18018
rect 400864 17954 400916 17960
rect 402980 18012 403032 18018
rect 402980 17954 403032 17960
rect 402992 16574 403020 17954
rect 402992 16546 403664 16574
rect 402520 14748 402572 14754
rect 402520 14690 402572 14696
rect 398932 3392 398984 3398
rect 398932 3334 398984 3340
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 398852 1958 398972 1986
rect 398944 480 398972 1958
rect 400140 480 400168 3334
rect 401324 3256 401376 3262
rect 401324 3198 401376 3204
rect 401336 480 401364 3198
rect 402532 480 402560 14690
rect 403636 480 403664 16546
rect 403716 12436 403768 12442
rect 403716 12378 403768 12384
rect 403728 3330 403756 12378
rect 403716 3324 403768 3330
rect 403716 3266 403768 3272
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 23122
rect 406016 3324 406068 3330
rect 406016 3266 406068 3272
rect 406028 480 406056 3266
rect 407224 480 407252 24618
rect 408512 16574 408540 76706
rect 412640 61396 412692 61402
rect 412640 61338 412692 61344
rect 409880 29640 409932 29646
rect 409880 29582 409932 29588
rect 409892 16574 409920 29582
rect 411260 26988 411312 26994
rect 411260 26930 411312 26936
rect 411272 16574 411300 26930
rect 408512 16546 409184 16574
rect 409892 16546 410840 16574
rect 411272 16546 411944 16574
rect 408408 3868 408460 3874
rect 408408 3810 408460 3816
rect 408420 480 408448 3810
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410812 480 410840 16546
rect 411916 480 411944 16546
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 61338
rect 425058 48920 425114 48929
rect 425058 48855 425114 48864
rect 418160 36576 418212 36582
rect 418160 36518 418212 36524
rect 414020 25628 414072 25634
rect 414020 25570 414072 25576
rect 414032 16574 414060 25570
rect 416780 24608 416832 24614
rect 416780 24550 416832 24556
rect 415400 20120 415452 20126
rect 415400 20062 415452 20068
rect 414032 16546 414336 16574
rect 414308 480 414336 16546
rect 415412 3210 415440 20062
rect 416792 16574 416820 24550
rect 418172 16574 418200 36518
rect 422298 22672 422354 22681
rect 422298 22607 422354 22616
rect 422312 16574 422340 22607
rect 423678 17368 423734 17377
rect 423678 17303 423734 17312
rect 416792 16546 417464 16574
rect 418172 16546 418568 16574
rect 422312 16546 422616 16574
rect 415492 15972 415544 15978
rect 415492 15914 415544 15920
rect 415504 3398 415532 15914
rect 415492 3392 415544 3398
rect 415492 3334 415544 3340
rect 416688 3392 416740 3398
rect 416688 3334 416740 3340
rect 415412 3182 415532 3210
rect 415504 480 415532 3182
rect 416700 480 416728 3334
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 420184 15904 420236 15910
rect 420184 15846 420236 15852
rect 420196 480 420224 15846
rect 420918 10296 420974 10305
rect 420918 10231 420974 10240
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 10231
rect 422588 480 422616 16546
rect 423692 3210 423720 17303
rect 425072 16574 425100 48855
rect 426452 16574 426480 78678
rect 430592 16574 430620 80038
rect 436744 78396 436796 78402
rect 436744 78338 436796 78344
rect 433340 76696 433392 76702
rect 433340 76638 433392 76644
rect 431958 61432 432014 61441
rect 431958 61367 432014 61376
rect 425072 16546 425744 16574
rect 426452 16546 426848 16574
rect 430592 16546 430896 16574
rect 423770 11928 423826 11937
rect 423770 11863 423826 11872
rect 423784 3398 423812 11863
rect 423772 3392 423824 3398
rect 423772 3334 423824 3340
rect 424968 3392 425020 3398
rect 424968 3334 425020 3340
rect 423692 3182 423812 3210
rect 423784 480 423812 3182
rect 424980 480 425008 3334
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 16546
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426820 354 426848 16546
rect 429200 14680 429252 14686
rect 429200 14622 429252 14628
rect 428464 12096 428516 12102
rect 428464 12038 428516 12044
rect 428476 480 428504 12038
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 426134 -960 426246 326
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429212 354 429240 14622
rect 430868 480 430896 16546
rect 431972 3398 432000 61367
rect 433352 16574 433380 76638
rect 436756 16574 436784 78338
rect 462332 78033 462360 703520
rect 478524 700398 478552 703520
rect 478512 700392 478564 700398
rect 478512 700334 478564 700340
rect 494072 141438 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 494060 141432 494112 141438
rect 494060 141374 494112 141380
rect 527192 79490 527220 703520
rect 543476 700330 543504 703520
rect 559668 702434 559696 703520
rect 558932 702406 559696 702434
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 558932 140078 558960 702406
rect 580262 697232 580318 697241
rect 580262 697167 580318 697176
rect 579618 683904 579674 683913
rect 579618 683839 579674 683848
rect 579632 683194 579660 683839
rect 579620 683188 579672 683194
rect 579620 683130 579672 683136
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 579710 630864 579766 630873
rect 579710 630799 579766 630808
rect 579724 630698 579752 630799
rect 579712 630692 579764 630698
rect 579712 630634 579764 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 579802 524512 579858 524521
rect 579802 524447 579804 524456
rect 579856 524447 579858 524456
rect 579804 524418 579856 524424
rect 579986 511320 580042 511329
rect 579986 511255 580042 511264
rect 580000 510678 580028 511255
rect 579988 510672 580040 510678
rect 579988 510614 580040 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579618 471472 579674 471481
rect 579618 471407 579674 471416
rect 579632 470626 579660 471407
rect 579620 470620 579672 470626
rect 579620 470562 579672 470568
rect 579618 458144 579674 458153
rect 579618 458079 579674 458088
rect 579632 456822 579660 458079
rect 579620 456816 579672 456822
rect 579620 456758 579672 456764
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580184 364410 580212 365055
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580184 311914 580212 312015
rect 580172 311908 580224 311914
rect 580172 311850 580224 311856
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580184 298178 580212 298687
rect 580172 298172 580224 298178
rect 580172 298114 580224 298120
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580184 271930 580212 272167
rect 580172 271924 580224 271930
rect 580172 271866 580224 271872
rect 579618 258904 579674 258913
rect 579618 258839 579674 258848
rect 579632 258126 579660 258839
rect 579620 258120 579672 258126
rect 579620 258062 579672 258068
rect 580170 245576 580226 245585
rect 580170 245511 580226 245520
rect 580184 244322 580212 245511
rect 580172 244316 580224 244322
rect 580172 244258 580224 244264
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 580184 218074 580212 218991
rect 580172 218068 580224 218074
rect 580172 218010 580224 218016
rect 580170 205728 580226 205737
rect 580170 205663 580172 205672
rect 580224 205663 580226 205672
rect 580172 205634 580224 205640
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580184 178090 580212 179143
rect 580172 178084 580224 178090
rect 580172 178026 580224 178032
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580184 165646 580212 165815
rect 580172 165640 580224 165646
rect 580172 165582 580224 165588
rect 579986 152688 580042 152697
rect 579986 152623 580042 152632
rect 580000 151842 580028 152623
rect 579988 151836 580040 151842
rect 579988 151778 580040 151784
rect 558920 140072 558972 140078
rect 558920 140014 558972 140020
rect 580170 139360 580226 139369
rect 580170 139295 580226 139304
rect 580184 138038 580212 139295
rect 580172 138032 580224 138038
rect 580172 137974 580224 137980
rect 579986 112840 580042 112849
rect 579986 112775 580042 112784
rect 580000 111858 580028 112775
rect 579988 111852 580040 111858
rect 579988 111794 580040 111800
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580184 99414 580212 99447
rect 580172 99408 580224 99414
rect 580172 99350 580224 99356
rect 580172 89140 580224 89146
rect 580172 89082 580224 89088
rect 554778 80336 554834 80345
rect 554778 80271 554834 80280
rect 527180 79484 527232 79490
rect 527180 79426 527232 79432
rect 483020 78260 483072 78266
rect 483020 78202 483072 78208
rect 462318 78024 462374 78033
rect 462318 77959 462374 77968
rect 480260 77308 480312 77314
rect 480260 77250 480312 77256
rect 471980 76628 472032 76634
rect 471980 76570 472032 76576
rect 440238 42120 440294 42129
rect 440238 42055 440294 42064
rect 433352 16546 434024 16574
rect 436756 16546 436876 16574
rect 432052 12028 432104 12034
rect 432052 11970 432104 11976
rect 431960 3392 432012 3398
rect 431960 3334 432012 3340
rect 432064 480 432092 11970
rect 433248 3392 433300 3398
rect 433248 3334 433300 3340
rect 433260 480 433288 3334
rect 429630 354 429742 480
rect 429212 326 429742 354
rect 429630 -960 429742 326
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 436744 14612 436796 14618
rect 436744 14554 436796 14560
rect 435088 11960 435140 11966
rect 435088 11902 435140 11908
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 11902
rect 436756 480 436784 14554
rect 436848 5030 436876 16546
rect 439136 14544 439188 14550
rect 439136 14486 439188 14492
rect 436836 5024 436888 5030
rect 436836 4966 436888 4972
rect 437940 3732 437992 3738
rect 437940 3674 437992 3680
rect 437952 480 437980 3674
rect 439148 480 439176 14486
rect 440252 3210 440280 42055
rect 447140 32632 447192 32638
rect 447140 32574 447192 32580
rect 447152 16574 447180 32574
rect 454040 21684 454092 21690
rect 454040 21626 454092 21632
rect 449900 20188 449952 20194
rect 449900 20130 449952 20136
rect 449912 16574 449940 20130
rect 447152 16546 447456 16574
rect 449912 16546 450952 16574
rect 442630 14784 442686 14793
rect 442630 14719 442686 14728
rect 440332 11892 440384 11898
rect 440332 11834 440384 11840
rect 440344 3398 440372 11834
rect 440332 3392 440384 3398
rect 440332 3334 440384 3340
rect 441528 3392 441580 3398
rect 441528 3334 441580 3340
rect 440252 3182 440372 3210
rect 440344 480 440372 3182
rect 441540 480 441568 3334
rect 442644 480 442672 14719
rect 443366 14648 443422 14657
rect 443366 14583 443422 14592
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 354 443408 14583
rect 445024 9580 445076 9586
rect 445024 9522 445076 9528
rect 445036 480 445064 9522
rect 446220 9444 446272 9450
rect 446220 9386 446272 9392
rect 446232 480 446260 9386
rect 447428 480 447456 16546
rect 449900 9512 449952 9518
rect 449900 9454 449952 9460
rect 448612 9376 448664 9382
rect 448612 9318 448664 9324
rect 448624 480 448652 9318
rect 449808 9308 449860 9314
rect 449808 9250 449860 9256
rect 449164 7608 449216 7614
rect 449164 7550 449216 7556
rect 449176 3806 449204 7550
rect 449164 3800 449216 3806
rect 449164 3742 449216 3748
rect 449820 480 449848 9250
rect 449912 3738 449940 9454
rect 449900 3732 449952 3738
rect 449900 3674 449952 3680
rect 450924 480 450952 16546
rect 452108 9240 452160 9246
rect 452108 9182 452160 9188
rect 452120 480 452148 9182
rect 453304 9172 453356 9178
rect 453304 9114 453356 9120
rect 453316 480 453344 9114
rect 443798 354 443910 480
rect 443380 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454052 354 454080 21626
rect 456800 20256 456852 20262
rect 456800 20198 456852 20204
rect 455696 9104 455748 9110
rect 455696 9046 455748 9052
rect 455708 480 455736 9046
rect 456812 3398 456840 20198
rect 471992 16574 472020 76570
rect 474004 32564 474056 32570
rect 474004 32506 474056 32512
rect 471992 16546 472296 16574
rect 468208 11824 468260 11830
rect 468208 11766 468260 11772
rect 465172 9648 465224 9654
rect 465172 9590 465224 9596
rect 456890 9072 456946 9081
rect 456890 9007 456946 9016
rect 463976 9036 464028 9042
rect 456800 3392 456852 3398
rect 456800 3334 456852 3340
rect 456904 480 456932 9007
rect 463976 8978 464028 8984
rect 459190 8936 459246 8945
rect 459190 8871 459246 8880
rect 458088 3392 458140 3398
rect 458088 3334 458140 3340
rect 458100 480 458128 3334
rect 459204 480 459232 8871
rect 460386 6352 460442 6361
rect 460386 6287 460442 6296
rect 460400 480 460428 6287
rect 461584 3664 461636 3670
rect 461584 3606 461636 3612
rect 461596 480 461624 3606
rect 462780 3596 462832 3602
rect 462780 3538 462832 3544
rect 462792 480 462820 3538
rect 463988 480 464016 8978
rect 465184 480 465212 9590
rect 467472 8968 467524 8974
rect 467472 8910 467524 8916
rect 466276 3528 466328 3534
rect 466276 3470 466328 3476
rect 466288 480 466316 3470
rect 467484 480 467512 8910
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468220 354 468248 11766
rect 471060 6248 471112 6254
rect 471060 6190 471112 6196
rect 469862 3904 469918 3913
rect 469862 3839 469918 3848
rect 469876 480 469904 3839
rect 471072 480 471100 6190
rect 472268 480 472296 16546
rect 473910 11792 473966 11801
rect 473910 11727 473966 11736
rect 473450 3768 473506 3777
rect 473450 3703 473506 3712
rect 473464 480 473492 3703
rect 473924 490 473952 11727
rect 474016 3534 474044 32506
rect 480272 16574 480300 77250
rect 481640 75336 481692 75342
rect 481640 75278 481692 75284
rect 480272 16546 480576 16574
rect 478142 11656 478198 11665
rect 478142 11591 478198 11600
rect 476946 3632 477002 3641
rect 476946 3567 477002 3576
rect 474004 3528 474056 3534
rect 474004 3470 474056 3476
rect 475750 3360 475806 3369
rect 475750 3295 475806 3304
rect 468638 354 468750 480
rect 468220 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 473924 462 474136 490
rect 475764 480 475792 3295
rect 476960 480 476988 3567
rect 478156 480 478184 11591
rect 479340 4956 479392 4962
rect 479340 4898 479392 4904
rect 479352 480 479380 4898
rect 480548 480 480576 16546
rect 481652 3602 481680 75278
rect 481732 62892 481784 62898
rect 481732 62834 481784 62840
rect 481640 3596 481692 3602
rect 481640 3538 481692 3544
rect 481744 480 481772 62834
rect 483032 16574 483060 78202
rect 498200 78192 498252 78198
rect 498200 78134 498252 78140
rect 496818 75304 496874 75313
rect 489920 75268 489972 75274
rect 496818 75239 496874 75248
rect 489920 75210 489972 75216
rect 484400 65680 484452 65686
rect 484400 65622 484452 65628
rect 484412 16574 484440 65622
rect 488540 47592 488592 47598
rect 488540 47534 488592 47540
rect 485780 32496 485832 32502
rect 485780 32438 485832 32444
rect 485792 16574 485820 32438
rect 488552 16574 488580 47534
rect 483032 16546 484072 16574
rect 484412 16546 484808 16574
rect 485792 16546 486464 16574
rect 488552 16546 488856 16574
rect 482468 3596 482520 3602
rect 482468 3538 482520 3544
rect 474108 354 474136 462
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482480 354 482508 3538
rect 484044 480 484072 16546
rect 482806 354 482918 480
rect 482480 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 486436 480 486464 16546
rect 487620 4888 487672 4894
rect 487620 4830 487672 4836
rect 487632 480 487660 4830
rect 488828 480 488856 16546
rect 489932 480 489960 75210
rect 494058 65512 494114 65521
rect 494058 65447 494114 65456
rect 492680 23112 492732 23118
rect 492680 23054 492732 23060
rect 492692 16574 492720 23054
rect 494072 16574 494100 65447
rect 495438 17232 495494 17241
rect 495438 17167 495494 17176
rect 492692 16546 493088 16574
rect 494072 16546 494744 16574
rect 492312 14476 492364 14482
rect 492312 14418 492364 14424
rect 491114 3496 491170 3505
rect 491114 3431 491170 3440
rect 491128 480 491156 3431
rect 492324 480 492352 14418
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494716 480 494744 16546
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 17167
rect 496832 16574 496860 75239
rect 496832 16546 497136 16574
rect 497108 480 497136 16546
rect 498212 480 498240 78134
rect 532700 78124 532752 78130
rect 532700 78066 532752 78072
rect 506480 75200 506532 75206
rect 506480 75142 506532 75148
rect 500960 71188 501012 71194
rect 500960 71130 501012 71136
rect 499580 31068 499632 31074
rect 499580 31010 499632 31016
rect 498292 18828 498344 18834
rect 498292 18770 498344 18776
rect 498304 16574 498332 18770
rect 499592 16574 499620 31010
rect 500972 16574 501000 71130
rect 505100 69896 505152 69902
rect 505100 69838 505152 69844
rect 503720 32428 503772 32434
rect 503720 32370 503772 32376
rect 502340 18760 502392 18766
rect 502340 18702 502392 18708
rect 502352 16574 502380 18702
rect 498304 16546 498976 16574
rect 499592 16546 500632 16574
rect 500972 16546 501368 16574
rect 502352 16546 503024 16574
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498948 354 498976 16546
rect 500604 480 500632 16546
rect 499366 354 499478 480
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501340 354 501368 16546
rect 502996 480 503024 16546
rect 501758 354 501870 480
rect 501340 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503732 354 503760 32370
rect 505112 16574 505140 69838
rect 505112 16546 505416 16574
rect 505388 480 505416 16546
rect 506492 3602 506520 75142
rect 507860 71120 507912 71126
rect 507860 71062 507912 71068
rect 506572 20052 506624 20058
rect 506572 19994 506624 20000
rect 506480 3596 506532 3602
rect 506480 3538 506532 3544
rect 506584 3482 506612 19994
rect 507872 16574 507900 71062
rect 523040 69828 523092 69834
rect 523040 69770 523092 69776
rect 511998 64152 512054 64161
rect 511998 64087 512054 64096
rect 509240 19984 509292 19990
rect 509240 19926 509292 19932
rect 509252 16574 509280 19926
rect 507872 16546 508912 16574
rect 509252 16546 509648 16574
rect 507308 3596 507360 3602
rect 507308 3538 507360 3544
rect 506492 3454 506612 3482
rect 506492 480 506520 3454
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507320 354 507348 3538
rect 508884 480 508912 16546
rect 507646 354 507758 480
rect 507320 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 511262 14512 511318 14521
rect 511262 14447 511318 14456
rect 511276 480 511304 14447
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 64087
rect 514760 62824 514812 62830
rect 514760 62766 514812 62772
rect 513378 19952 513434 19961
rect 513378 19887 513434 19896
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 19887
rect 514772 3534 514800 62766
rect 514850 32464 514906 32473
rect 514850 32399 514906 32408
rect 514760 3528 514812 3534
rect 514760 3470 514812 3476
rect 514864 3346 514892 32399
rect 516140 21616 516192 21622
rect 516140 21558 516192 21564
rect 516152 16574 516180 21558
rect 520280 21548 520332 21554
rect 520280 21490 520332 21496
rect 516152 16546 517192 16574
rect 515588 3528 515640 3534
rect 515588 3470 515640 3476
rect 514772 3318 514892 3346
rect 514772 480 514800 3318
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515600 354 515628 3470
rect 517164 480 517192 16546
rect 518348 3596 518400 3602
rect 518348 3538 518400 3544
rect 518360 480 518388 3538
rect 519544 3460 519596 3466
rect 519544 3402 519596 3408
rect 519556 480 519584 3402
rect 515926 354 516038 480
rect 515600 326 516038 354
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520292 354 520320 21490
rect 521844 3800 521896 3806
rect 521844 3742 521896 3748
rect 521856 480 521884 3742
rect 523052 480 523080 69770
rect 525800 68468 525852 68474
rect 525800 68410 525852 68416
rect 523132 21480 523184 21486
rect 523132 21422 523184 21428
rect 523144 16574 523172 21422
rect 525812 16574 525840 68410
rect 529938 67008 529994 67017
rect 529938 66943 529994 66952
rect 527180 21412 527232 21418
rect 527180 21354 527232 21360
rect 527192 16574 527220 21354
rect 523144 16546 523816 16574
rect 525812 16546 526208 16574
rect 527192 16546 527864 16574
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 520710 -960 520822 326
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 523788 354 523816 16546
rect 525432 3732 525484 3738
rect 525432 3674 525484 3680
rect 525444 480 525472 3674
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527836 480 527864 16546
rect 529018 5128 529074 5137
rect 529018 5063 529074 5072
rect 529032 480 529060 5063
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 529952 354 529980 66943
rect 531318 21312 531374 21321
rect 531318 21247 531374 21256
rect 531332 480 531360 21247
rect 532712 16574 532740 78066
rect 549258 75168 549314 75177
rect 549258 75103 549314 75112
rect 539600 71052 539652 71058
rect 539600 70994 539652 71000
rect 536840 69760 536892 69766
rect 536840 69702 536892 69708
rect 535460 25560 535512 25566
rect 535460 25502 535512 25508
rect 534080 23044 534132 23050
rect 534080 22986 534132 22992
rect 534092 16574 534120 22986
rect 535472 16574 535500 25502
rect 536852 16574 536880 69702
rect 538220 22976 538272 22982
rect 538220 22918 538272 22924
rect 532712 16546 533752 16574
rect 534092 16546 534488 16574
rect 535472 16546 536144 16574
rect 536852 16546 537248 16574
rect 532054 13016 532110 13025
rect 532054 12951 532110 12960
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532068 354 532096 12951
rect 533724 480 533752 16546
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536116 480 536144 16546
rect 537220 480 537248 16546
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 22918
rect 539612 3534 539640 70994
rect 547878 66872 547934 66881
rect 547878 66807 547934 66816
rect 543740 65612 543792 65618
rect 543740 65554 543792 65560
rect 539692 28280 539744 28286
rect 539692 28222 539744 28228
rect 539600 3528 539652 3534
rect 539600 3470 539652 3476
rect 539704 3346 539732 28222
rect 540980 22908 541032 22914
rect 540980 22850 541032 22856
rect 540992 16574 541020 22850
rect 543752 16574 543780 65554
rect 545120 22840 545172 22846
rect 545120 22782 545172 22788
rect 545132 16574 545160 22782
rect 546498 18592 546554 18601
rect 546498 18527 546554 18536
rect 540992 16546 542032 16574
rect 543752 16546 544424 16574
rect 545132 16546 545528 16574
rect 540428 3528 540480 3534
rect 540428 3470 540480 3476
rect 539612 3318 539732 3346
rect 539612 480 539640 3318
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540440 354 540468 3470
rect 542004 480 542032 16546
rect 542728 10328 542780 10334
rect 542728 10270 542780 10276
rect 540766 354 540878 480
rect 540440 326 540878 354
rect 540766 -960 540878 326
rect 541962 -960 542074 480
rect 542740 354 542768 10270
rect 544396 480 544424 16546
rect 545500 480 545528 16546
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 18527
rect 547892 480 547920 66807
rect 549272 16574 549300 75103
rect 550638 47560 550694 47569
rect 550638 47495 550694 47504
rect 550652 16574 550680 47495
rect 552020 24540 552072 24546
rect 552020 24482 552072 24488
rect 552032 16574 552060 24482
rect 553400 18692 553452 18698
rect 553400 18634 553452 18640
rect 553412 16574 553440 18634
rect 549272 16546 550312 16574
rect 550652 16546 551048 16574
rect 552032 16546 552704 16574
rect 553412 16546 553808 16574
rect 549074 6216 549130 6225
rect 549074 6151 549130 6160
rect 549088 480 549116 6151
rect 550284 480 550312 16546
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 552676 480 552704 16546
rect 553780 480 553808 16546
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 80271
rect 580184 79354 580212 89082
rect 580276 79393 580304 697167
rect 580538 670712 580594 670721
rect 580538 670647 580594 670656
rect 580354 591016 580410 591025
rect 580354 590951 580410 590960
rect 580368 80850 580396 590951
rect 580446 431624 580502 431633
rect 580446 431559 580502 431568
rect 580356 80844 580408 80850
rect 580356 80786 580408 80792
rect 580460 79801 580488 431559
rect 580552 431254 580580 670647
rect 580540 431248 580592 431254
rect 580540 431190 580592 431196
rect 580538 378448 580594 378457
rect 580538 378383 580594 378392
rect 580446 79792 580502 79801
rect 580446 79727 580502 79736
rect 580552 79422 580580 378383
rect 580630 325272 580686 325281
rect 580630 325207 580686 325216
rect 580644 89146 580672 325207
rect 580722 232384 580778 232393
rect 580722 232319 580778 232328
rect 580632 89140 580684 89146
rect 580632 89082 580684 89088
rect 580632 89004 580684 89010
rect 580632 88946 580684 88952
rect 580644 80617 580672 88946
rect 580736 80782 580764 232319
rect 580814 192536 580870 192545
rect 580814 192471 580870 192480
rect 580724 80776 580776 80782
rect 580724 80718 580776 80724
rect 580828 80714 580856 192471
rect 580906 126032 580962 126041
rect 580906 125967 580962 125976
rect 580920 89010 580948 125967
rect 580908 89004 580960 89010
rect 580908 88946 580960 88952
rect 580906 86184 580962 86193
rect 580906 86119 580962 86128
rect 580816 80708 580868 80714
rect 580816 80650 580868 80656
rect 580630 80608 580686 80617
rect 580630 80543 580686 80552
rect 580920 80481 580948 86119
rect 580906 80472 580962 80481
rect 580906 80407 580962 80416
rect 580540 79416 580592 79422
rect 580262 79384 580318 79393
rect 580172 79348 580224 79354
rect 580540 79358 580592 79364
rect 580262 79319 580318 79328
rect 580172 79290 580224 79296
rect 574744 78056 574796 78062
rect 574744 77998 574796 78004
rect 558920 76560 558972 76566
rect 558920 76502 558972 76508
rect 565818 76528 565874 76537
rect 557540 68400 557592 68406
rect 557540 68342 557592 68348
rect 556160 24472 556212 24478
rect 556160 24414 556212 24420
rect 556172 480 556200 24414
rect 556252 18624 556304 18630
rect 556252 18566 556304 18572
rect 556264 16574 556292 18566
rect 557552 16574 557580 68342
rect 558932 16574 558960 76502
rect 565818 76463 565874 76472
rect 564440 69692 564492 69698
rect 564440 69634 564492 69640
rect 560300 26920 560352 26926
rect 560300 26862 560352 26868
rect 560312 16574 560340 26862
rect 563060 24404 563112 24410
rect 563060 24346 563112 24352
rect 556264 16546 556936 16574
rect 557552 16546 558592 16574
rect 558932 16546 559328 16574
rect 560312 16546 560432 16574
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 558564 480 558592 16546
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16546
rect 562048 4820 562100 4826
rect 562048 4762 562100 4768
rect 562060 480 562088 4762
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563072 354 563100 24346
rect 564452 3534 564480 69634
rect 564532 68332 564584 68338
rect 564532 68274 564584 68280
rect 564440 3528 564492 3534
rect 564440 3470 564492 3476
rect 564544 3346 564572 68274
rect 565832 16574 565860 76463
rect 572720 65544 572772 65550
rect 572720 65486 572772 65492
rect 568580 64184 568632 64190
rect 568580 64126 568632 64132
rect 567198 29608 567254 29617
rect 567198 29543 567254 29552
rect 567212 16574 567240 29543
rect 568592 16574 568620 64126
rect 569960 24268 570012 24274
rect 569960 24210 570012 24216
rect 569972 16574 570000 24210
rect 571340 24200 571392 24206
rect 571340 24142 571392 24148
rect 565832 16546 566872 16574
rect 567212 16546 567608 16574
rect 568592 16546 568712 16574
rect 569972 16546 570368 16574
rect 565268 3528 565320 3534
rect 565268 3470 565320 3476
rect 564452 3318 564572 3346
rect 564452 480 564480 3318
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565280 354 565308 3470
rect 566844 480 566872 16546
rect 565606 354 565718 480
rect 565280 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 568684 354 568712 16546
rect 570340 480 570368 16546
rect 569102 354 569214 480
rect 568684 326 569214 354
rect 567998 -960 568110 326
rect 569102 -960 569214 326
rect 570298 -960 570410 480
rect 571352 354 571380 24142
rect 572732 480 572760 65486
rect 572812 24132 572864 24138
rect 572812 24074 572864 24080
rect 572824 16574 572852 24074
rect 572824 16546 573496 16574
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573468 354 573496 16546
rect 574652 11756 574704 11762
rect 574652 11698 574704 11704
rect 574664 3482 574692 11698
rect 574756 3602 574784 77998
rect 581092 77988 581144 77994
rect 581092 77930 581144 77936
rect 578238 73808 578294 73817
rect 578238 73743 578294 73752
rect 578252 16574 578280 73743
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 579620 24336 579672 24342
rect 579620 24278 579672 24284
rect 579632 19825 579660 24278
rect 580264 22772 580316 22778
rect 580264 22714 580316 22720
rect 579618 19816 579674 19825
rect 579618 19751 579674 19760
rect 578252 16546 578648 16574
rect 576308 6180 576360 6186
rect 576308 6122 576360 6128
rect 574744 3596 574796 3602
rect 574744 3538 574796 3544
rect 574664 3454 575152 3482
rect 575124 480 575152 3454
rect 576320 480 576348 6122
rect 577410 4992 577466 5001
rect 577410 4927 577466 4936
rect 577424 480 577452 4927
rect 578620 480 578648 16546
rect 580276 6633 580304 22714
rect 581104 16574 581132 77930
rect 581104 16546 581776 16574
rect 580262 6624 580318 6633
rect 580262 6559 580318 6568
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 581012 480 581040 3402
rect 573886 354 573998 480
rect 573468 326 573998 354
rect 573886 -960 573998 326
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581748 354 581776 16546
rect 583390 4856 583446 4865
rect 583390 4791 583446 4800
rect 583404 480 583432 4791
rect 582166 354 582278 480
rect 581748 326 582278 354
rect 582166 -960 582278 326
rect 583362 -960 583474 480
<< via2 >>
rect 2778 684256 2834 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3054 566888 3110 566944
rect 3238 449520 3294 449576
rect 2962 423544 3018 423600
rect 3054 410488 3110 410544
rect 3054 397432 3110 397488
rect 3330 371320 3386 371376
rect 3330 358400 3386 358456
rect 3330 319232 3386 319288
rect 3330 306176 3386 306232
rect 3330 267144 3386 267200
rect 3330 254088 3386 254144
rect 3330 241032 3386 241088
rect 3330 214920 3386 214976
rect 3330 201864 3386 201920
rect 3330 188808 3386 188864
rect 3514 632068 3516 632088
rect 3516 632068 3568 632088
rect 3568 632068 3570 632088
rect 3514 632032 3570 632068
rect 3514 619112 3570 619168
rect 3606 606056 3662 606112
rect 3514 579944 3570 580000
rect 3514 527876 3570 527912
rect 3514 527856 3516 527876
rect 3516 527856 3568 527876
rect 3568 527856 3570 527876
rect 3514 514820 3570 514856
rect 3514 514800 3516 514820
rect 3516 514800 3568 514820
rect 3568 514800 3570 514820
rect 3514 475632 3570 475688
rect 3514 462576 3570 462632
rect 3514 162868 3516 162888
rect 3516 162868 3568 162888
rect 3568 162868 3570 162888
rect 3514 162832 3570 162868
rect 3514 149776 3570 149832
rect 3514 136720 3570 136776
rect 3330 110608 3386 110664
rect 3514 97552 3570 97608
rect 3514 84632 3570 84688
rect 3790 553832 3846 553888
rect 3698 345344 3754 345400
rect 3974 501744 4030 501800
rect 3882 293120 3938 293176
rect 3790 79328 3846 79384
rect 3974 79464 4030 79520
rect 3606 79192 3662 79248
rect 3422 79056 3478 79112
rect 3238 78920 3294 78976
rect 3054 78784 3110 78840
rect 2778 75248 2834 75304
rect 1398 75112 1454 75168
rect 3422 71612 3424 71632
rect 3424 71612 3476 71632
rect 3476 71612 3478 71632
rect 3422 71576 3478 71612
rect 3054 58520 3110 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3422 32408 3478 32464
rect 3330 19352 3386 19408
rect 3422 6432 3478 6488
rect 4066 4800 4122 4856
rect 117318 137536 117374 137592
rect 117318 136040 117374 136096
rect 117318 134544 117374 134600
rect 117410 133048 117466 133104
rect 117318 131552 117374 131608
rect 117318 130056 117374 130112
rect 117318 128560 117374 128616
rect 117318 127064 117374 127120
rect 117318 125568 117374 125624
rect 117318 124108 117320 124128
rect 117320 124108 117372 124128
rect 117372 124108 117374 124128
rect 117318 124072 117374 124108
rect 117318 122576 117374 122632
rect 117318 121080 117374 121136
rect 117318 119584 117374 119640
rect 117318 118088 117374 118144
rect 117318 116592 117374 116648
rect 117318 115096 117374 115152
rect 118054 113600 118110 113656
rect 118238 92656 118294 92712
rect 118146 91160 118202 91216
rect 118330 89664 118386 89720
rect 119066 112104 119122 112160
rect 119158 110608 119214 110664
rect 119250 109112 119306 109168
rect 118974 107616 119030 107672
rect 118882 106120 118938 106176
rect 118790 104624 118846 104680
rect 118698 103128 118754 103184
rect 118606 95648 118662 95704
rect 118514 94152 118570 94208
rect 118422 88168 118478 88224
rect 118422 86672 118478 86728
rect 118330 82184 118386 82240
rect 71778 77152 71834 77208
rect 37278 76608 37334 76664
rect 20718 76472 20774 76528
rect 20626 4936 20682 4992
rect 42798 19896 42854 19952
rect 41878 8880 41934 8936
rect 40682 6160 40738 6216
rect 57978 73888 58034 73944
rect 53838 73752 53894 73808
rect 57242 9152 57298 9208
rect 56046 9016 56102 9072
rect 89718 75520 89774 75576
rect 75918 75384 75974 75440
rect 71778 74024 71834 74080
rect 74998 10240 75054 10296
rect 73802 6296 73858 6352
rect 91098 44784 91154 44840
rect 92478 10376 92534 10432
rect 111798 76744 111854 76800
rect 110510 10512 110566 10568
rect 109314 7520 109370 7576
rect 111614 7656 111670 7712
rect 118606 85176 118662 85232
rect 118514 83680 118570 83736
rect 118422 80552 118478 80608
rect 118606 80416 118662 80472
rect 120722 102040 120778 102096
rect 120814 100680 120870 100736
rect 120906 98640 120962 98696
rect 120998 97144 121054 97200
rect 179602 126792 179658 126848
rect 179510 120672 179566 120728
rect 179694 119312 179750 119368
rect 179418 116592 179474 116648
rect 179878 130464 179934 130520
rect 179786 112512 179842 112568
rect 124678 80144 124734 80200
rect 119342 78512 119398 78568
rect 124954 79600 125010 79656
rect 125506 79736 125562 79792
rect 125736 79906 125792 79962
rect 125920 79906 125976 79962
rect 125690 78648 125746 78704
rect 125874 78648 125930 78704
rect 126380 79906 126436 79962
rect 126288 79736 126344 79792
rect 126840 79872 126896 79928
rect 127116 79906 127172 79962
rect 126150 78648 126206 78704
rect 126426 78648 126482 78704
rect 127070 79736 127126 79792
rect 127300 79872 127356 79928
rect 127576 79872 127632 79928
rect 127944 79906 128000 79962
rect 126978 79600 127034 79656
rect 127714 79736 127770 79792
rect 128128 79906 128184 79962
rect 127530 79600 127586 79656
rect 127254 76472 127310 76528
rect 127622 22616 127678 22672
rect 127990 79600 128046 79656
rect 127990 78376 128046 78432
rect 128680 79872 128736 79928
rect 128956 79906 129012 79962
rect 128864 79736 128920 79792
rect 129186 79736 129242 79792
rect 129508 79906 129564 79962
rect 129692 79872 129748 79928
rect 129876 79872 129932 79928
rect 130336 79906 130392 79962
rect 128726 78376 128782 78432
rect 128450 76608 128506 76664
rect 129186 77696 129242 77752
rect 129370 79620 129426 79656
rect 129370 79600 129372 79620
rect 129372 79600 129424 79620
rect 129424 79600 129426 79620
rect 129370 78376 129426 78432
rect 129830 79600 129886 79656
rect 129738 78376 129794 78432
rect 130014 78240 130070 78296
rect 129646 77016 129702 77072
rect 130198 78376 130254 78432
rect 130382 75112 130438 75168
rect 131624 79872 131680 79928
rect 131440 79772 131442 79792
rect 131442 79772 131494 79792
rect 131494 79772 131496 79792
rect 131440 79736 131496 79772
rect 132360 79872 132416 79928
rect 131210 79600 131266 79656
rect 131118 78376 131174 78432
rect 130934 78240 130990 78296
rect 132544 79906 132600 79962
rect 131302 77968 131358 78024
rect 132682 77968 132738 78024
rect 133142 77832 133198 77888
rect 133878 79736 133934 79792
rect 134292 79872 134348 79928
rect 134660 79872 134716 79928
rect 134936 79906 134992 79962
rect 135488 79906 135544 79962
rect 135856 79906 135912 79962
rect 133878 76744 133934 76800
rect 134154 77968 134210 78024
rect 134062 77832 134118 77888
rect 134338 79600 134394 79656
rect 133970 75248 134026 75304
rect 134798 79600 134854 79656
rect 135350 79772 135352 79792
rect 135352 79772 135404 79792
rect 135404 79772 135406 79792
rect 135350 79736 135406 79772
rect 135534 79736 135590 79792
rect 136408 79872 136464 79928
rect 135350 79600 135406 79656
rect 135534 78376 135590 78432
rect 135442 78240 135498 78296
rect 135442 75248 135498 75304
rect 136592 79906 136648 79962
rect 136960 79906 137016 79962
rect 136270 79600 136326 79656
rect 136546 78376 136602 78432
rect 137972 79906 138028 79962
rect 138156 79906 138212 79962
rect 138616 79872 138672 79928
rect 138064 79736 138120 79792
rect 137926 78376 137982 78432
rect 138294 79736 138350 79792
rect 139168 79872 139224 79928
rect 139444 79906 139500 79962
rect 138846 79600 138902 79656
rect 139122 79636 139124 79656
rect 139124 79636 139176 79656
rect 139176 79636 139178 79656
rect 139122 79600 139178 79636
rect 139030 78240 139086 78296
rect 139398 78376 139454 78432
rect 139582 79736 139638 79792
rect 139674 79600 139730 79656
rect 140548 79872 140604 79928
rect 140732 79906 140788 79962
rect 140916 79906 140972 79962
rect 139950 77832 140006 77888
rect 140410 78240 140466 78296
rect 140502 78104 140558 78160
rect 140686 78104 140742 78160
rect 140594 77968 140650 78024
rect 141376 79906 141432 79962
rect 142020 79906 142076 79962
rect 142112 79736 142168 79792
rect 142296 79872 142352 79928
rect 142066 79600 142122 79656
rect 142848 79872 142904 79928
rect 142434 77968 142490 78024
rect 143216 79872 143272 79928
rect 143400 79906 143456 79962
rect 143768 79906 143824 79962
rect 142894 79600 142950 79656
rect 143170 79600 143226 79656
rect 143630 79600 143686 79656
rect 143354 78376 143410 78432
rect 144504 79772 144506 79792
rect 144506 79772 144558 79792
rect 144558 79772 144560 79792
rect 144504 79736 144560 79772
rect 144872 79906 144928 79962
rect 144826 79736 144882 79792
rect 145608 79906 145664 79962
rect 144458 79620 144514 79656
rect 144458 79600 144460 79620
rect 144460 79600 144512 79620
rect 144512 79600 144514 79620
rect 144642 78376 144698 78432
rect 145838 79736 145894 79792
rect 145470 79600 145526 79656
rect 146252 79906 146308 79962
rect 146206 79600 146262 79656
rect 146022 77560 146078 77616
rect 146390 76744 146446 76800
rect 147448 79906 147504 79962
rect 147310 79736 147366 79792
rect 147632 79872 147688 79928
rect 148184 79906 148240 79962
rect 147816 79736 147872 79792
rect 147586 78376 147642 78432
rect 147954 79600 148010 79656
rect 147678 76608 147734 76664
rect 148138 79600 148194 79656
rect 147954 78376 148010 78432
rect 148644 79906 148700 79962
rect 148828 79872 148884 79928
rect 149288 79872 149344 79928
rect 149564 79872 149620 79928
rect 149748 79906 149804 79962
rect 150116 79906 150172 79962
rect 150484 79906 150540 79962
rect 150208 79770 150264 79826
rect 148874 78240 148930 78296
rect 149058 78104 149114 78160
rect 148782 77968 148838 78024
rect 149426 79600 149482 79656
rect 150070 79600 150126 79656
rect 149610 78376 149666 78432
rect 149978 78376 150034 78432
rect 151128 79872 151184 79928
rect 151680 79906 151736 79962
rect 152048 79872 152104 79928
rect 150254 78240 150310 78296
rect 150714 79600 150770 79656
rect 151174 79600 151230 79656
rect 151772 79736 151828 79792
rect 152416 79872 152472 79928
rect 152784 79906 152840 79962
rect 153060 79906 153116 79962
rect 151818 79600 151874 79656
rect 151634 78104 151690 78160
rect 152738 78376 152794 78432
rect 153198 78376 153254 78432
rect 153014 78240 153070 78296
rect 153198 78104 153254 78160
rect 153704 79906 153760 79962
rect 153888 79906 153944 79962
rect 154164 79872 154220 79928
rect 154348 79872 154404 79928
rect 153934 79600 153990 79656
rect 154210 79636 154212 79656
rect 154212 79636 154264 79656
rect 154264 79636 154266 79656
rect 154210 79600 154266 79636
rect 154808 79906 154864 79962
rect 154992 79906 155048 79962
rect 154946 79736 155002 79792
rect 154118 77968 154174 78024
rect 154026 77832 154082 77888
rect 154394 78240 154450 78296
rect 154578 78104 154634 78160
rect 154762 79600 154818 79656
rect 154670 75520 154726 75576
rect 155636 79906 155692 79962
rect 155682 79736 155738 79792
rect 156096 79872 156152 79928
rect 156464 79906 156520 79962
rect 156648 79872 156704 79928
rect 156924 79872 156980 79928
rect 157108 79906 157164 79962
rect 156142 77968 156198 78024
rect 156786 79636 156788 79656
rect 156788 79636 156840 79656
rect 156840 79636 156842 79656
rect 156786 79600 156842 79636
rect 156694 78648 156750 78704
rect 156878 74024 156934 74080
rect 157430 79736 157486 79792
rect 157752 79872 157808 79928
rect 158212 79872 158268 79928
rect 157154 78648 157210 78704
rect 157062 77560 157118 77616
rect 157798 79736 157854 79792
rect 157936 79736 157992 79792
rect 157430 78376 157486 78432
rect 157338 78240 157394 78296
rect 157706 78376 157762 78432
rect 158488 79838 158544 79894
rect 158948 79872 159004 79928
rect 158166 78376 158222 78432
rect 158442 77968 158498 78024
rect 158350 77016 158406 77072
rect 158810 78240 158866 78296
rect 158442 75248 158498 75304
rect 159270 79736 159326 79792
rect 159408 79770 159464 79826
rect 159776 79872 159832 79928
rect 159960 79872 160016 79928
rect 159868 79736 159924 79792
rect 160696 79906 160752 79962
rect 159730 77968 159786 78024
rect 160006 79600 160062 79656
rect 160006 75112 160062 75168
rect 154486 4936 154542 4992
rect 158902 4800 158958 4856
rect 160098 19896 160154 19952
rect 160880 79772 160882 79792
rect 160882 79772 160934 79792
rect 160934 79772 160936 79792
rect 160880 79736 160936 79772
rect 161064 79906 161120 79962
rect 161432 79906 161488 79962
rect 161616 79906 161672 79962
rect 161800 79872 161856 79928
rect 162168 79906 162224 79962
rect 162536 79906 162592 79962
rect 160650 79600 160706 79656
rect 160742 78104 160798 78160
rect 161202 77424 161258 77480
rect 161110 75248 161166 75304
rect 161478 78920 161534 78976
rect 161570 78648 161626 78704
rect 161570 3848 161626 3904
rect 161846 79600 161902 79656
rect 161754 75248 161810 75304
rect 162720 79906 162776 79962
rect 162306 79620 162362 79656
rect 162306 79600 162308 79620
rect 162308 79600 162360 79620
rect 162360 79600 162362 79620
rect 162398 77832 162454 77888
rect 162582 79600 162638 79656
rect 162674 79464 162730 79520
rect 163272 79872 163328 79928
rect 162766 78104 162822 78160
rect 162582 77424 162638 77480
rect 162582 75248 162638 75304
rect 161294 3440 161350 3496
rect 163640 79872 163696 79928
rect 163824 79872 163880 79928
rect 163594 79736 163650 79792
rect 163318 79600 163374 79656
rect 163778 79600 163834 79656
rect 164560 79838 164616 79894
rect 163962 75248 164018 75304
rect 164146 75248 164202 75304
rect 165112 79872 165168 79928
rect 164422 75928 164478 75984
rect 165066 79600 165122 79656
rect 165250 77832 165306 77888
rect 165710 79736 165766 79792
rect 165940 79872 165996 79928
rect 166400 79872 166456 79928
rect 166676 79906 166732 79962
rect 165434 79600 165490 79656
rect 165342 77424 165398 77480
rect 165526 78376 165582 78432
rect 165526 77832 165582 77888
rect 166584 79736 166640 79792
rect 166952 79906 167008 79962
rect 167228 79872 167284 79928
rect 166078 76472 166134 76528
rect 166814 78376 166870 78432
rect 166814 77424 166870 77480
rect 166722 77288 166778 77344
rect 167596 79872 167652 79928
rect 167182 77716 167238 77752
rect 167182 77696 167184 77716
rect 167184 77696 167236 77716
rect 167236 77696 167238 77716
rect 168332 79872 168388 79928
rect 168700 79906 168756 79962
rect 168148 79736 168204 79792
rect 167550 77288 167606 77344
rect 168010 77968 168066 78024
rect 168102 77560 168158 77616
rect 168378 78668 168434 78704
rect 168378 78648 168380 78668
rect 168380 78648 168432 78668
rect 168432 78648 168434 78668
rect 168378 78376 168434 78432
rect 168378 78104 168434 78160
rect 168194 77288 168250 77344
rect 168654 77424 168710 77480
rect 169436 79872 169492 79928
rect 169712 79906 169768 79962
rect 170080 79872 170136 79928
rect 170356 79906 170412 79962
rect 169666 78784 169722 78840
rect 170034 79600 170090 79656
rect 170034 79056 170090 79112
rect 170218 77288 170274 77344
rect 171000 79872 171056 79928
rect 170908 79736 170964 79792
rect 171276 79872 171332 79928
rect 170954 79056 171010 79112
rect 170862 78920 170918 78976
rect 170770 78240 170826 78296
rect 170770 77968 170826 78024
rect 170494 76336 170550 76392
rect 170310 73752 170366 73808
rect 171138 78240 171194 78296
rect 171736 79906 171792 79962
rect 171874 79600 171930 79656
rect 171506 79056 171562 79112
rect 171046 76200 171102 76256
rect 172196 79906 172252 79962
rect 171782 78376 171838 78432
rect 172840 79872 172896 79928
rect 173208 79872 173264 79928
rect 173392 79906 173448 79962
rect 171874 77832 171930 77888
rect 170402 3440 170458 3496
rect 171966 75112 172022 75168
rect 172242 77560 172298 77616
rect 173346 79736 173402 79792
rect 173162 79464 173218 79520
rect 173346 79328 173402 79384
rect 173254 79192 173310 79248
rect 173438 78784 173494 78840
rect 173714 78920 173770 78976
rect 173622 78648 173678 78704
rect 173898 78512 173954 78568
rect 174174 78376 174230 78432
rect 172886 77152 172942 77208
rect 173162 77016 173218 77072
rect 173346 76880 173402 76936
rect 173898 75792 173954 75848
rect 175002 79600 175058 79656
rect 176106 80008 176162 80064
rect 176198 79056 176254 79112
rect 176198 78104 176254 78160
rect 175462 77968 175518 78024
rect 178774 77288 178830 77344
rect 175278 68448 175334 68504
rect 176658 32544 176714 32600
rect 181258 129648 181314 129704
rect 181166 121488 181222 121544
rect 181074 117408 181130 117464
rect 180982 114688 181038 114744
rect 180890 113328 180946 113384
rect 180798 110608 180854 110664
rect 180154 78240 180210 78296
rect 181534 128288 181590 128344
rect 182362 125568 182418 125624
rect 182270 124208 182326 124264
rect 182178 122848 182234 122904
rect 181442 109248 181498 109304
rect 182730 103808 182786 103864
rect 182270 101088 182326 101144
rect 182454 99728 182510 99784
rect 182178 98368 182234 98424
rect 182546 97008 182602 97064
rect 182546 91568 182602 91624
rect 183006 92928 183062 92984
rect 183006 80688 183062 80744
rect 182822 77288 182878 77344
rect 183466 107888 183522 107944
rect 183466 106528 183522 106584
rect 183466 105168 183522 105224
rect 183466 102448 183522 102504
rect 183466 95648 183522 95704
rect 183466 94288 183522 94344
rect 183466 90208 183522 90264
rect 183374 88848 183430 88904
rect 183466 87488 183522 87544
rect 183374 86128 183430 86184
rect 183466 84768 183522 84824
rect 183466 83408 183522 83464
rect 183282 82048 183338 82104
rect 193862 75656 193918 75712
rect 194598 74432 194654 74488
rect 193218 68312 193274 68368
rect 191838 34040 191894 34096
rect 193310 25472 193366 25528
rect 212538 17584 212594 17640
rect 230478 74296 230534 74352
rect 226430 33904 226486 33960
rect 229374 13368 229430 13424
rect 228730 6024 228786 6080
rect 247038 76744 247094 76800
rect 244278 74160 244334 74216
rect 245658 58520 245714 58576
rect 248418 20032 248474 20088
rect 263598 62736 263654 62792
rect 266358 33768 266414 33824
rect 265346 9560 265402 9616
rect 282918 76608 282974 76664
rect 296074 72528 296130 72584
rect 281906 9424 281962 9480
rect 280710 6840 280766 6896
rect 284298 6704 284354 6760
rect 298098 72392 298154 72448
rect 306930 71032 306986 71088
rect 300858 17448 300914 17504
rect 299662 9288 299718 9344
rect 300766 6568 300822 6624
rect 317418 29824 317474 29880
rect 339130 75520 339186 75576
rect 316038 10376 316094 10432
rect 315026 9152 315082 9208
rect 316222 7520 316278 7576
rect 369122 75384 369178 75440
rect 349802 74024 349858 74080
rect 353298 68176 353354 68232
rect 351918 51720 351974 51776
rect 349158 29688 349214 29744
rect 351642 6432 351698 6488
rect 372618 35128 372674 35184
rect 365718 15816 365774 15872
rect 370134 13232 370190 13288
rect 371238 13096 371294 13152
rect 378414 73888 378470 73944
rect 425058 48864 425114 48920
rect 422298 22616 422354 22672
rect 423678 17312 423734 17368
rect 420918 10240 420974 10296
rect 431958 61376 432014 61432
rect 423770 11872 423826 11928
rect 580262 697176 580318 697232
rect 579618 683848 579674 683904
rect 580170 644000 580226 644056
rect 579710 630808 579766 630864
rect 580170 617480 580226 617536
rect 580170 577632 580226 577688
rect 580170 564304 580226 564360
rect 580170 537784 580226 537840
rect 579802 524476 579858 524512
rect 579802 524456 579804 524476
rect 579804 524456 579856 524476
rect 579856 524456 579858 524476
rect 579986 511264 580042 511320
rect 580170 484608 580226 484664
rect 579618 471416 579674 471472
rect 579618 458088 579674 458144
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 580170 365064 580226 365120
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 579618 258848 579674 258904
rect 580170 245520 580226 245576
rect 580170 219000 580226 219056
rect 580170 205692 580226 205728
rect 580170 205672 580172 205692
rect 580172 205672 580224 205692
rect 580224 205672 580226 205692
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 579986 152632 580042 152688
rect 580170 139304 580226 139360
rect 579986 112784 580042 112840
rect 580170 99456 580226 99512
rect 554778 80280 554834 80336
rect 462318 77968 462374 78024
rect 440238 42064 440294 42120
rect 442630 14728 442686 14784
rect 443366 14592 443422 14648
rect 456890 9016 456946 9072
rect 459190 8880 459246 8936
rect 460386 6296 460442 6352
rect 469862 3848 469918 3904
rect 473910 11736 473966 11792
rect 473450 3712 473506 3768
rect 478142 11600 478198 11656
rect 476946 3576 477002 3632
rect 475750 3304 475806 3360
rect 496818 75248 496874 75304
rect 494058 65456 494114 65512
rect 495438 17176 495494 17232
rect 491114 3440 491170 3496
rect 511998 64096 512054 64152
rect 511262 14456 511318 14512
rect 513378 19896 513434 19952
rect 514850 32408 514906 32464
rect 529938 66952 529994 67008
rect 529018 5072 529074 5128
rect 531318 21256 531374 21312
rect 549258 75112 549314 75168
rect 532054 12960 532110 13016
rect 547878 66816 547934 66872
rect 546498 18536 546554 18592
rect 550638 47504 550694 47560
rect 549074 6160 549130 6216
rect 580538 670656 580594 670712
rect 580354 590960 580410 591016
rect 580446 431568 580502 431624
rect 580538 378392 580594 378448
rect 580446 79736 580502 79792
rect 580630 325216 580686 325272
rect 580722 232328 580778 232384
rect 580814 192480 580870 192536
rect 580906 125976 580962 126032
rect 580906 86128 580962 86184
rect 580630 80552 580686 80608
rect 580906 80416 580962 80472
rect 580262 79328 580318 79384
rect 565818 76472 565874 76528
rect 567198 29552 567254 29608
rect 578238 73752 578294 73808
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579618 19760 579674 19816
rect 577410 4936 577466 4992
rect 580262 6568 580318 6624
rect 583390 4800 583446 4856
<< metal3 >>
rect -960 697220 480 697460
rect 580257 697234 580323 697237
rect 583520 697234 584960 697324
rect 580257 697232 584960 697234
rect 580257 697176 580262 697232
rect 580318 697176 584960 697232
rect 580257 697174 584960 697176
rect 580257 697171 580323 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 2773 684314 2839 684317
rect -960 684312 2839 684314
rect -960 684256 2778 684312
rect 2834 684256 2839 684312
rect -960 684254 2839 684256
rect -960 684164 480 684254
rect 2773 684251 2839 684254
rect 579613 683906 579679 683909
rect 583520 683906 584960 683996
rect 579613 683904 584960 683906
rect 579613 683848 579618 683904
rect 579674 683848 584960 683904
rect 579613 683846 584960 683848
rect 579613 683843 579679 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580533 670714 580599 670717
rect 583520 670714 584960 670804
rect 580533 670712 584960 670714
rect 580533 670656 580538 670712
rect 580594 670656 584960 670712
rect 580533 670654 584960 670656
rect 580533 670651 580599 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3509 632090 3575 632093
rect -960 632088 3575 632090
rect -960 632032 3514 632088
rect 3570 632032 3575 632088
rect -960 632030 3575 632032
rect -960 631940 480 632030
rect 3509 632027 3575 632030
rect 579705 630866 579771 630869
rect 583520 630866 584960 630956
rect 579705 630864 584960 630866
rect 579705 630808 579710 630864
rect 579766 630808 584960 630864
rect 579705 630806 584960 630808
rect 579705 630803 579771 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3601 606114 3667 606117
rect -960 606112 3667 606114
rect -960 606056 3606 606112
rect 3662 606056 3667 606112
rect -960 606054 3667 606056
rect -960 605964 480 606054
rect 3601 606051 3667 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580349 591018 580415 591021
rect 583520 591018 584960 591108
rect 580349 591016 584960 591018
rect 580349 590960 580354 591016
rect 580410 590960 584960 591016
rect 580349 590958 584960 590960
rect 580349 590955 580415 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3509 580002 3575 580005
rect -960 580000 3575 580002
rect -960 579944 3514 580000
rect 3570 579944 3575 580000
rect -960 579942 3575 579944
rect -960 579852 480 579942
rect 3509 579939 3575 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3049 566946 3115 566949
rect -960 566944 3115 566946
rect -960 566888 3054 566944
rect 3110 566888 3115 566944
rect -960 566886 3115 566888
rect -960 566796 480 566886
rect 3049 566883 3115 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3785 553890 3851 553893
rect -960 553888 3851 553890
rect -960 553832 3790 553888
rect 3846 553832 3851 553888
rect -960 553830 3851 553832
rect -960 553740 480 553830
rect 3785 553827 3851 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3509 527914 3575 527917
rect -960 527912 3575 527914
rect -960 527856 3514 527912
rect 3570 527856 3575 527912
rect -960 527854 3575 527856
rect -960 527764 480 527854
rect 3509 527851 3575 527854
rect 579797 524514 579863 524517
rect 583520 524514 584960 524604
rect 579797 524512 584960 524514
rect 579797 524456 579802 524512
rect 579858 524456 584960 524512
rect 579797 524454 584960 524456
rect 579797 524451 579863 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 579981 511322 580047 511325
rect 583520 511322 584960 511412
rect 579981 511320 584960 511322
rect 579981 511264 579986 511320
rect 580042 511264 584960 511320
rect 579981 511262 584960 511264
rect 579981 511259 580047 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3969 501802 4035 501805
rect -960 501800 4035 501802
rect -960 501744 3974 501800
rect 4030 501744 4035 501800
rect -960 501742 4035 501744
rect -960 501652 480 501742
rect 3969 501739 4035 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3509 475690 3575 475693
rect -960 475688 3575 475690
rect -960 475632 3514 475688
rect 3570 475632 3575 475688
rect -960 475630 3575 475632
rect -960 475540 480 475630
rect 3509 475627 3575 475630
rect 579613 471474 579679 471477
rect 583520 471474 584960 471564
rect 579613 471472 584960 471474
rect 579613 471416 579618 471472
rect 579674 471416 584960 471472
rect 579613 471414 584960 471416
rect 579613 471411 579679 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 579613 458146 579679 458149
rect 583520 458146 584960 458236
rect 579613 458144 584960 458146
rect 579613 458088 579618 458144
rect 579674 458088 584960 458144
rect 579613 458086 584960 458088
rect 579613 458083 579679 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3233 449578 3299 449581
rect -960 449576 3299 449578
rect -960 449520 3238 449576
rect 3294 449520 3299 449576
rect -960 449518 3299 449520
rect -960 449428 480 449518
rect 3233 449515 3299 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580441 431626 580507 431629
rect 583520 431626 584960 431716
rect 580441 431624 584960 431626
rect 580441 431568 580446 431624
rect 580502 431568 584960 431624
rect 580441 431566 584960 431568
rect 580441 431563 580507 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 2957 423602 3023 423605
rect -960 423600 3023 423602
rect -960 423544 2962 423600
rect 3018 423544 3023 423600
rect -960 423542 3023 423544
rect -960 423452 480 423542
rect 2957 423539 3023 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3049 410546 3115 410549
rect -960 410544 3115 410546
rect -960 410488 3054 410544
rect 3110 410488 3115 410544
rect -960 410486 3115 410488
rect -960 410396 480 410486
rect 3049 410483 3115 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3049 397490 3115 397493
rect -960 397488 3115 397490
rect -960 397432 3054 397488
rect 3110 397432 3115 397488
rect -960 397430 3115 397432
rect -960 397340 480 397430
rect 3049 397427 3115 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580533 378450 580599 378453
rect 583520 378450 584960 378540
rect 580533 378448 584960 378450
rect 580533 378392 580538 378448
rect 580594 378392 584960 378448
rect 580533 378390 584960 378392
rect 580533 378387 580599 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3693 345402 3759 345405
rect -960 345400 3759 345402
rect -960 345344 3698 345400
rect 3754 345344 3759 345400
rect -960 345342 3759 345344
rect -960 345252 480 345342
rect 3693 345339 3759 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580625 325274 580691 325277
rect 583520 325274 584960 325364
rect 580625 325272 584960 325274
rect 580625 325216 580630 325272
rect 580686 325216 584960 325272
rect 580625 325214 584960 325216
rect 580625 325211 580691 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3325 306234 3391 306237
rect -960 306232 3391 306234
rect -960 306176 3330 306232
rect 3386 306176 3391 306232
rect -960 306174 3391 306176
rect -960 306084 480 306174
rect 3325 306171 3391 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3877 293178 3943 293181
rect -960 293176 3943 293178
rect -960 293120 3882 293176
rect 3938 293120 3943 293176
rect -960 293118 3943 293120
rect -960 293028 480 293118
rect 3877 293115 3943 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3325 267202 3391 267205
rect -960 267200 3391 267202
rect -960 267144 3330 267200
rect 3386 267144 3391 267200
rect -960 267142 3391 267144
rect -960 267052 480 267142
rect 3325 267139 3391 267142
rect 579613 258906 579679 258909
rect 583520 258906 584960 258996
rect 579613 258904 584960 258906
rect 579613 258848 579618 258904
rect 579674 258848 584960 258904
rect 579613 258846 584960 258848
rect 579613 258843 579679 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3325 254146 3391 254149
rect -960 254144 3391 254146
rect -960 254088 3330 254144
rect 3386 254088 3391 254144
rect -960 254086 3391 254088
rect -960 253996 480 254086
rect 3325 254083 3391 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3325 241090 3391 241093
rect -960 241088 3391 241090
rect -960 241032 3330 241088
rect 3386 241032 3391 241088
rect -960 241030 3391 241032
rect -960 240940 480 241030
rect 3325 241027 3391 241030
rect 580717 232386 580783 232389
rect 583520 232386 584960 232476
rect 580717 232384 584960 232386
rect 580717 232328 580722 232384
rect 580778 232328 584960 232384
rect 580717 232326 584960 232328
rect 580717 232323 580783 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3325 201922 3391 201925
rect -960 201920 3391 201922
rect -960 201864 3330 201920
rect 3386 201864 3391 201920
rect -960 201862 3391 201864
rect -960 201772 480 201862
rect 3325 201859 3391 201862
rect 580809 192538 580875 192541
rect 583520 192538 584960 192628
rect 580809 192536 584960 192538
rect 580809 192480 580814 192536
rect 580870 192480 584960 192536
rect 580809 192478 584960 192480
rect 580809 192475 580875 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3325 188866 3391 188869
rect -960 188864 3391 188866
rect -960 188808 3330 188864
rect 3386 188808 3391 188864
rect -960 188806 3391 188808
rect -960 188716 480 188806
rect 3325 188803 3391 188806
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3509 162890 3575 162893
rect -960 162888 3575 162890
rect -960 162832 3514 162888
rect 3570 162832 3575 162888
rect -960 162830 3575 162832
rect -960 162740 480 162830
rect 3509 162827 3575 162830
rect 579981 152690 580047 152693
rect 583520 152690 584960 152780
rect 579981 152688 584960 152690
rect 579981 152632 579986 152688
rect 580042 152632 584960 152688
rect 579981 152630 584960 152632
rect 579981 152627 580047 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3509 149834 3575 149837
rect -960 149832 3575 149834
rect -960 149776 3514 149832
rect 3570 149776 3575 149832
rect -960 149774 3575 149776
rect -960 149684 480 149774
rect 3509 149771 3575 149774
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect 117313 137594 117379 137597
rect 117313 137592 120060 137594
rect 117313 137536 117318 137592
rect 117374 137536 120060 137592
rect 117313 137534 120060 137536
rect 117313 137531 117379 137534
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 117313 136098 117379 136101
rect 117313 136096 120060 136098
rect 117313 136040 117318 136096
rect 117374 136040 120060 136096
rect 117313 136038 120060 136040
rect 117313 136035 117379 136038
rect 117313 134602 117379 134605
rect 117313 134600 120060 134602
rect 117313 134544 117318 134600
rect 117374 134544 120060 134600
rect 117313 134542 120060 134544
rect 117313 134539 117379 134542
rect 117405 133106 117471 133109
rect 117405 133104 120060 133106
rect 117405 133048 117410 133104
rect 117466 133048 120060 133104
rect 117405 133046 120060 133048
rect 117405 133043 117471 133046
rect 117313 131610 117379 131613
rect 117313 131608 120060 131610
rect 117313 131552 117318 131608
rect 117374 131552 120060 131608
rect 117313 131550 120060 131552
rect 117313 131547 117379 131550
rect 179830 130525 179890 131036
rect 179830 130520 179939 130525
rect 179830 130464 179878 130520
rect 179934 130464 179939 130520
rect 179830 130462 179939 130464
rect 179873 130459 179939 130462
rect 117313 130114 117379 130117
rect 117313 130112 120060 130114
rect 117313 130056 117318 130112
rect 117374 130056 120060 130112
rect 117313 130054 120060 130056
rect 117313 130051 117379 130054
rect 181253 129706 181319 129709
rect 179860 129704 181319 129706
rect 179860 129648 181258 129704
rect 181314 129648 181319 129704
rect 179860 129646 181319 129648
rect 181253 129643 181319 129646
rect 117313 128618 117379 128621
rect 117313 128616 120060 128618
rect 117313 128560 117318 128616
rect 117374 128560 120060 128616
rect 117313 128558 120060 128560
rect 117313 128555 117379 128558
rect 181529 128346 181595 128349
rect 179860 128344 181595 128346
rect 179860 128288 181534 128344
rect 181590 128288 181595 128344
rect 179860 128286 181595 128288
rect 181529 128283 181595 128286
rect 117313 127122 117379 127125
rect 117313 127120 120060 127122
rect 117313 127064 117318 127120
rect 117374 127064 120060 127120
rect 117313 127062 120060 127064
rect 117313 127059 117379 127062
rect 179646 126853 179706 126956
rect 179597 126848 179706 126853
rect 179597 126792 179602 126848
rect 179658 126792 179706 126848
rect 179597 126790 179706 126792
rect 179597 126787 179663 126790
rect 580901 126034 580967 126037
rect 583520 126034 584960 126124
rect 580901 126032 584960 126034
rect 580901 125976 580906 126032
rect 580962 125976 584960 126032
rect 580901 125974 584960 125976
rect 580901 125971 580967 125974
rect 583520 125884 584960 125974
rect 117313 125626 117379 125629
rect 182357 125626 182423 125629
rect 117313 125624 120060 125626
rect 117313 125568 117318 125624
rect 117374 125568 120060 125624
rect 117313 125566 120060 125568
rect 179860 125624 182423 125626
rect 179860 125568 182362 125624
rect 182418 125568 182423 125624
rect 179860 125566 182423 125568
rect 117313 125563 117379 125566
rect 182357 125563 182423 125566
rect 182265 124266 182331 124269
rect 179860 124264 182331 124266
rect 179860 124208 182270 124264
rect 182326 124208 182331 124264
rect 179860 124206 182331 124208
rect 182265 124203 182331 124206
rect 117313 124130 117379 124133
rect 117313 124128 120060 124130
rect 117313 124072 117318 124128
rect 117374 124072 120060 124128
rect 117313 124070 120060 124072
rect 117313 124067 117379 124070
rect -960 123572 480 123812
rect 182173 122906 182239 122909
rect 179860 122904 182239 122906
rect 179860 122848 182178 122904
rect 182234 122848 182239 122904
rect 179860 122846 182239 122848
rect 182173 122843 182239 122846
rect 117313 122634 117379 122637
rect 117313 122632 120060 122634
rect 117313 122576 117318 122632
rect 117374 122576 120060 122632
rect 117313 122574 120060 122576
rect 117313 122571 117379 122574
rect 181161 121546 181227 121549
rect 179860 121544 181227 121546
rect 179860 121488 181166 121544
rect 181222 121488 181227 121544
rect 179860 121486 181227 121488
rect 181161 121483 181227 121486
rect 117313 121138 117379 121141
rect 117313 121136 120060 121138
rect 117313 121080 117318 121136
rect 117374 121080 120060 121136
rect 117313 121078 120060 121080
rect 117313 121075 117379 121078
rect 179505 120730 179571 120733
rect 179462 120728 179571 120730
rect 179462 120672 179510 120728
rect 179566 120672 179571 120728
rect 179462 120667 179571 120672
rect 179462 120156 179522 120667
rect 117313 119642 117379 119645
rect 117313 119640 120060 119642
rect 117313 119584 117318 119640
rect 117374 119584 120060 119640
rect 117313 119582 120060 119584
rect 117313 119579 117379 119582
rect 179689 119370 179755 119373
rect 179646 119368 179755 119370
rect 179646 119312 179694 119368
rect 179750 119312 179755 119368
rect 179646 119307 179755 119312
rect 179646 118796 179706 119307
rect 117313 118146 117379 118149
rect 117313 118144 120060 118146
rect 117313 118088 117318 118144
rect 117374 118088 120060 118144
rect 117313 118086 120060 118088
rect 117313 118083 117379 118086
rect 181069 117466 181135 117469
rect 179860 117464 181135 117466
rect 179860 117408 181074 117464
rect 181130 117408 181135 117464
rect 179860 117406 181135 117408
rect 181069 117403 181135 117406
rect 117313 116650 117379 116653
rect 179413 116650 179479 116653
rect 117313 116648 120060 116650
rect 117313 116592 117318 116648
rect 117374 116592 120060 116648
rect 117313 116590 120060 116592
rect 179413 116648 179522 116650
rect 179413 116592 179418 116648
rect 179474 116592 179522 116648
rect 117313 116587 117379 116590
rect 179413 116587 179522 116592
rect 179462 116076 179522 116587
rect 117313 115154 117379 115157
rect 117313 115152 120060 115154
rect 117313 115096 117318 115152
rect 117374 115096 120060 115152
rect 117313 115094 120060 115096
rect 117313 115091 117379 115094
rect 180977 114746 181043 114749
rect 179860 114744 181043 114746
rect 179860 114688 180982 114744
rect 181038 114688 181043 114744
rect 179860 114686 181043 114688
rect 180977 114683 181043 114686
rect 118049 113658 118115 113661
rect 118049 113656 120060 113658
rect 118049 113600 118054 113656
rect 118110 113600 120060 113656
rect 118049 113598 120060 113600
rect 118049 113595 118115 113598
rect 180885 113386 180951 113389
rect 179860 113384 180951 113386
rect 179860 113328 180890 113384
rect 180946 113328 180951 113384
rect 179860 113326 180951 113328
rect 180885 113323 180951 113326
rect 579981 112842 580047 112845
rect 583520 112842 584960 112932
rect 579981 112840 584960 112842
rect 579981 112784 579986 112840
rect 580042 112784 584960 112840
rect 579981 112782 584960 112784
rect 579981 112779 580047 112782
rect 583520 112692 584960 112782
rect 179781 112570 179847 112573
rect 179781 112568 179890 112570
rect 179781 112512 179786 112568
rect 179842 112512 179890 112568
rect 179781 112507 179890 112512
rect 119061 112162 119127 112165
rect 119061 112160 120060 112162
rect 119061 112104 119066 112160
rect 119122 112104 120060 112160
rect 119061 112102 120060 112104
rect 119061 112099 119127 112102
rect 179830 111996 179890 112507
rect -960 110666 480 110756
rect 3325 110666 3391 110669
rect -960 110664 3391 110666
rect -960 110608 3330 110664
rect 3386 110608 3391 110664
rect -960 110606 3391 110608
rect -960 110516 480 110606
rect 3325 110603 3391 110606
rect 119153 110666 119219 110669
rect 180793 110666 180859 110669
rect 119153 110664 120060 110666
rect 119153 110608 119158 110664
rect 119214 110608 120060 110664
rect 119153 110606 120060 110608
rect 179860 110664 180859 110666
rect 179860 110608 180798 110664
rect 180854 110608 180859 110664
rect 179860 110606 180859 110608
rect 119153 110603 119219 110606
rect 180793 110603 180859 110606
rect 181437 109306 181503 109309
rect 179860 109304 181503 109306
rect 179860 109248 181442 109304
rect 181498 109248 181503 109304
rect 179860 109246 181503 109248
rect 181437 109243 181503 109246
rect 119245 109170 119311 109173
rect 119245 109168 120060 109170
rect 119245 109112 119250 109168
rect 119306 109112 120060 109168
rect 119245 109110 120060 109112
rect 119245 109107 119311 109110
rect 183461 107946 183527 107949
rect 179860 107944 183527 107946
rect 179860 107888 183466 107944
rect 183522 107888 183527 107944
rect 179860 107886 183527 107888
rect 183461 107883 183527 107886
rect 118969 107674 119035 107677
rect 118969 107672 120060 107674
rect 118969 107616 118974 107672
rect 119030 107616 120060 107672
rect 118969 107614 120060 107616
rect 118969 107611 119035 107614
rect 183461 106586 183527 106589
rect 179860 106584 183527 106586
rect 179860 106528 183466 106584
rect 183522 106528 183527 106584
rect 179860 106526 183527 106528
rect 183461 106523 183527 106526
rect 118877 106178 118943 106181
rect 118877 106176 120060 106178
rect 118877 106120 118882 106176
rect 118938 106120 120060 106176
rect 118877 106118 120060 106120
rect 118877 106115 118943 106118
rect 183461 105226 183527 105229
rect 179860 105224 183527 105226
rect 179860 105168 183466 105224
rect 183522 105168 183527 105224
rect 179860 105166 183527 105168
rect 183461 105163 183527 105166
rect 118785 104682 118851 104685
rect 118785 104680 120060 104682
rect 118785 104624 118790 104680
rect 118846 104624 120060 104680
rect 118785 104622 120060 104624
rect 118785 104619 118851 104622
rect 182725 103866 182791 103869
rect 179860 103864 182791 103866
rect 179860 103808 182730 103864
rect 182786 103808 182791 103864
rect 179860 103806 182791 103808
rect 182725 103803 182791 103806
rect 118693 103186 118759 103189
rect 118693 103184 120060 103186
rect 118693 103128 118698 103184
rect 118754 103128 120060 103184
rect 118693 103126 120060 103128
rect 118693 103123 118759 103126
rect 183461 102506 183527 102509
rect 179860 102504 183527 102506
rect 179860 102448 183466 102504
rect 183522 102448 183527 102504
rect 179860 102446 183527 102448
rect 183461 102443 183527 102446
rect 120717 102098 120783 102101
rect 120582 102096 120783 102098
rect 120582 102040 120722 102096
rect 120778 102040 120783 102096
rect 120582 102038 120783 102040
rect 120582 101660 120642 102038
rect 120717 102035 120783 102038
rect 182265 101146 182331 101149
rect 179860 101144 182331 101146
rect 179860 101088 182270 101144
rect 182326 101088 182331 101144
rect 179860 101086 182331 101088
rect 182265 101083 182331 101086
rect 120809 100738 120875 100741
rect 120582 100736 120875 100738
rect 120582 100680 120814 100736
rect 120870 100680 120875 100736
rect 120582 100678 120875 100680
rect 120582 100164 120642 100678
rect 120809 100675 120875 100678
rect 182449 99786 182515 99789
rect 179860 99784 182515 99786
rect 179860 99728 182454 99784
rect 182510 99728 182515 99784
rect 179860 99726 182515 99728
rect 182449 99723 182515 99726
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect 120901 98698 120967 98701
rect 120612 98696 120967 98698
rect 120612 98640 120906 98696
rect 120962 98640 120967 98696
rect 120612 98638 120967 98640
rect 120901 98635 120967 98638
rect 182173 98426 182239 98429
rect 179860 98424 182239 98426
rect 179860 98368 182178 98424
rect 182234 98368 182239 98424
rect 179860 98366 182239 98368
rect 182173 98363 182239 98366
rect -960 97610 480 97700
rect 3509 97610 3575 97613
rect -960 97608 3575 97610
rect -960 97552 3514 97608
rect 3570 97552 3575 97608
rect -960 97550 3575 97552
rect -960 97460 480 97550
rect 3509 97547 3575 97550
rect 120993 97202 121059 97205
rect 120612 97200 121059 97202
rect 120612 97144 120998 97200
rect 121054 97144 121059 97200
rect 120612 97142 121059 97144
rect 120993 97139 121059 97142
rect 182541 97066 182607 97069
rect 179860 97064 182607 97066
rect 179860 97008 182546 97064
rect 182602 97008 182607 97064
rect 179860 97006 182607 97008
rect 182541 97003 182607 97006
rect 118601 95706 118667 95709
rect 183461 95706 183527 95709
rect 118601 95704 120060 95706
rect 118601 95648 118606 95704
rect 118662 95648 120060 95704
rect 118601 95646 120060 95648
rect 179860 95704 183527 95706
rect 179860 95648 183466 95704
rect 183522 95648 183527 95704
rect 179860 95646 183527 95648
rect 118601 95643 118667 95646
rect 183461 95643 183527 95646
rect 183461 94346 183527 94349
rect 179860 94344 183527 94346
rect 179860 94288 183466 94344
rect 183522 94288 183527 94344
rect 179860 94286 183527 94288
rect 183461 94283 183527 94286
rect 118509 94210 118575 94213
rect 118509 94208 120060 94210
rect 118509 94152 118514 94208
rect 118570 94152 120060 94208
rect 118509 94150 120060 94152
rect 118509 94147 118575 94150
rect 183001 92986 183067 92989
rect 179860 92984 183067 92986
rect 179860 92928 183006 92984
rect 183062 92928 183067 92984
rect 179860 92926 183067 92928
rect 183001 92923 183067 92926
rect 118233 92714 118299 92717
rect 118233 92712 120060 92714
rect 118233 92656 118238 92712
rect 118294 92656 120060 92712
rect 118233 92654 120060 92656
rect 118233 92651 118299 92654
rect 182541 91626 182607 91629
rect 179860 91624 182607 91626
rect 179860 91568 182546 91624
rect 182602 91568 182607 91624
rect 179860 91566 182607 91568
rect 182541 91563 182607 91566
rect 118141 91218 118207 91221
rect 118141 91216 120060 91218
rect 118141 91160 118146 91216
rect 118202 91160 120060 91216
rect 118141 91158 120060 91160
rect 118141 91155 118207 91158
rect 183461 90266 183527 90269
rect 179860 90264 183527 90266
rect 179860 90208 183466 90264
rect 183522 90208 183527 90264
rect 179860 90206 183527 90208
rect 183461 90203 183527 90206
rect 118325 89722 118391 89725
rect 118325 89720 120060 89722
rect 118325 89664 118330 89720
rect 118386 89664 120060 89720
rect 118325 89662 120060 89664
rect 118325 89659 118391 89662
rect 183369 88906 183435 88909
rect 179860 88904 183435 88906
rect 179860 88848 183374 88904
rect 183430 88848 183435 88904
rect 179860 88846 183435 88848
rect 183369 88843 183435 88846
rect 118417 88226 118483 88229
rect 118417 88224 120060 88226
rect 118417 88168 118422 88224
rect 118478 88168 120060 88224
rect 118417 88166 120060 88168
rect 118417 88163 118483 88166
rect 183461 87546 183527 87549
rect 179860 87544 183527 87546
rect 179860 87488 183466 87544
rect 183522 87488 183527 87544
rect 179860 87486 183527 87488
rect 183461 87483 183527 87486
rect 118417 86730 118483 86733
rect 118417 86728 120060 86730
rect 118417 86672 118422 86728
rect 118478 86672 120060 86728
rect 118417 86670 120060 86672
rect 118417 86667 118483 86670
rect 183369 86186 183435 86189
rect 179860 86184 183435 86186
rect 179860 86128 183374 86184
rect 183430 86128 183435 86184
rect 179860 86126 183435 86128
rect 183369 86123 183435 86126
rect 580901 86186 580967 86189
rect 583520 86186 584960 86276
rect 580901 86184 584960 86186
rect 580901 86128 580906 86184
rect 580962 86128 584960 86184
rect 580901 86126 584960 86128
rect 580901 86123 580967 86126
rect 583520 86036 584960 86126
rect 118601 85234 118667 85237
rect 118601 85232 120060 85234
rect 118601 85176 118606 85232
rect 118662 85176 120060 85232
rect 118601 85174 120060 85176
rect 118601 85171 118667 85174
rect 183461 84826 183527 84829
rect 179860 84824 183527 84826
rect -960 84690 480 84780
rect 179860 84768 183466 84824
rect 183522 84768 183527 84824
rect 179860 84766 183527 84768
rect 183461 84763 183527 84766
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 118509 83738 118575 83741
rect 118509 83736 120060 83738
rect 118509 83680 118514 83736
rect 118570 83680 120060 83736
rect 118509 83678 120060 83680
rect 118509 83675 118575 83678
rect 183461 83466 183527 83469
rect 179860 83464 183527 83466
rect 179860 83408 183466 83464
rect 183522 83408 183527 83464
rect 179860 83406 183527 83408
rect 183461 83403 183527 83406
rect 118325 82242 118391 82245
rect 118325 82240 120060 82242
rect 118325 82184 118330 82240
rect 118386 82184 120060 82240
rect 118325 82182 120060 82184
rect 118325 82179 118391 82182
rect 183277 82106 183343 82109
rect 179860 82104 183343 82106
rect 179860 82048 183282 82104
rect 183338 82048 183343 82104
rect 179860 82046 183343 82048
rect 183277 82043 183343 82046
rect 183001 80746 183067 80749
rect 179860 80744 183067 80746
rect 179860 80688 183006 80744
rect 183062 80688 183067 80744
rect 179860 80686 183067 80688
rect 183001 80683 183067 80686
rect 118417 80610 118483 80613
rect 580625 80610 580691 80613
rect 118417 80608 580691 80610
rect 118417 80552 118422 80608
rect 118478 80552 580630 80608
rect 580686 80552 580691 80608
rect 118417 80550 580691 80552
rect 118417 80547 118483 80550
rect 580625 80547 580691 80550
rect 118601 80474 118667 80477
rect 580901 80474 580967 80477
rect 118601 80472 580967 80474
rect 118601 80416 118606 80472
rect 118662 80416 580906 80472
rect 580962 80416 580967 80472
rect 118601 80414 580967 80416
rect 118601 80411 118667 80414
rect 580901 80411 580967 80414
rect 554773 80338 554839 80341
rect 168698 80336 554839 80338
rect 168698 80280 554778 80336
rect 554834 80280 554839 80336
rect 168698 80278 554839 80280
rect 124673 80202 124739 80205
rect 124673 80200 128370 80202
rect 124673 80144 124678 80200
rect 124734 80144 128370 80200
rect 124673 80142 128370 80144
rect 124673 80139 124739 80142
rect 125731 79962 125797 79967
rect 125731 79932 125736 79962
rect 125792 79932 125797 79962
rect 125915 79962 125981 79967
rect 125726 79868 125732 79932
rect 125796 79930 125802 79932
rect 125796 79870 125854 79930
rect 125915 79906 125920 79962
rect 125976 79906 125981 79962
rect 125915 79901 125981 79906
rect 126375 79964 126441 79967
rect 127111 79964 127177 79967
rect 126375 79962 126714 79964
rect 126375 79906 126380 79962
rect 126436 79932 126714 79962
rect 127068 79962 127177 79964
rect 126436 79906 126652 79932
rect 126375 79904 126652 79906
rect 126375 79901 126441 79904
rect 125796 79868 125802 79870
rect 125501 79794 125567 79797
rect 125918 79794 125978 79901
rect 126646 79868 126652 79904
rect 126716 79868 126722 79932
rect 126835 79928 126901 79933
rect 127068 79932 127116 79962
rect 126835 79872 126840 79928
rect 126896 79872 126901 79928
rect 126835 79867 126901 79872
rect 127014 79868 127020 79932
rect 127084 79906 127116 79932
rect 127172 79906 127177 79962
rect 127939 79962 128005 79967
rect 127084 79901 127177 79906
rect 127295 79930 127361 79933
rect 127295 79928 127404 79930
rect 127084 79870 127128 79901
rect 127295 79872 127300 79928
rect 127356 79872 127404 79928
rect 127084 79868 127090 79870
rect 127295 79867 127404 79872
rect 127571 79928 127637 79933
rect 127939 79932 127944 79962
rect 128000 79932 128005 79962
rect 128123 79962 128189 79967
rect 127571 79872 127576 79928
rect 127632 79872 127637 79928
rect 127571 79867 127637 79872
rect 127934 79868 127940 79932
rect 128004 79930 128010 79932
rect 128004 79870 128062 79930
rect 128123 79906 128128 79962
rect 128184 79906 128189 79962
rect 128123 79901 128189 79906
rect 128004 79868 128010 79870
rect 126283 79796 126349 79797
rect 126278 79794 126284 79796
rect 125501 79792 125978 79794
rect 125501 79736 125506 79792
rect 125562 79736 125978 79792
rect 125501 79734 125978 79736
rect 126192 79734 126284 79794
rect 125501 79731 125567 79734
rect 126278 79732 126284 79734
rect 126348 79732 126354 79796
rect 126838 79794 126898 79867
rect 127065 79794 127131 79797
rect 126838 79792 127131 79794
rect 126838 79736 127070 79792
rect 127126 79736 127131 79792
rect 126838 79734 127131 79736
rect 126283 79731 126349 79732
rect 127065 79731 127131 79734
rect 124949 79658 125015 79661
rect 126973 79658 127039 79661
rect 124949 79656 127039 79658
rect 124949 79600 124954 79656
rect 125010 79600 126978 79656
rect 127034 79600 127039 79656
rect 124949 79598 127039 79600
rect 127344 79658 127404 79867
rect 127574 79794 127634 79867
rect 127709 79794 127775 79797
rect 127574 79792 127775 79794
rect 127574 79736 127714 79792
rect 127770 79736 127775 79792
rect 127574 79734 127775 79736
rect 127709 79731 127775 79734
rect 127525 79658 127591 79661
rect 127344 79656 127591 79658
rect 127344 79600 127530 79656
rect 127586 79600 127591 79656
rect 127344 79598 127591 79600
rect 124949 79595 125015 79598
rect 126973 79595 127039 79598
rect 127525 79595 127591 79598
rect 127985 79658 128051 79661
rect 128126 79658 128186 79901
rect 127985 79656 128186 79658
rect 127985 79600 127990 79656
rect 128046 79600 128186 79656
rect 127985 79598 128186 79600
rect 128310 79658 128370 80142
rect 145414 80140 145420 80204
rect 145484 80202 145490 80204
rect 145484 80142 146264 80202
rect 145484 80140 145490 80142
rect 140446 80066 140452 80068
rect 140408 80004 140452 80066
rect 140516 80004 140522 80068
rect 128951 79964 129017 79967
rect 129503 79964 129569 79967
rect 128951 79962 129244 79964
rect 128486 79868 128492 79932
rect 128556 79930 128562 79932
rect 128675 79930 128741 79933
rect 128556 79928 128741 79930
rect 128556 79872 128680 79928
rect 128736 79872 128741 79928
rect 128951 79906 128956 79962
rect 129012 79906 129244 79962
rect 129460 79962 129569 79964
rect 129460 79932 129508 79962
rect 128951 79904 129244 79906
rect 128951 79901 129017 79904
rect 128556 79870 128741 79872
rect 128556 79868 128562 79870
rect 128675 79867 128741 79870
rect 129184 79797 129244 79904
rect 129406 79868 129412 79932
rect 129476 79906 129508 79932
rect 129564 79906 129569 79962
rect 130331 79962 130397 79967
rect 129476 79901 129569 79906
rect 129687 79928 129753 79933
rect 129476 79870 129520 79901
rect 129687 79872 129692 79928
rect 129748 79872 129753 79928
rect 129476 79868 129482 79870
rect 129687 79867 129753 79872
rect 129871 79930 129937 79933
rect 130331 79932 130336 79962
rect 130392 79932 130397 79962
rect 132539 79962 132605 79967
rect 129871 79928 130072 79930
rect 129871 79872 129876 79928
rect 129932 79872 130072 79928
rect 129871 79870 130072 79872
rect 129871 79867 129937 79870
rect 128859 79796 128925 79797
rect 128854 79794 128860 79796
rect 128768 79734 128860 79794
rect 128854 79732 128860 79734
rect 128924 79732 128930 79796
rect 129181 79792 129247 79797
rect 129181 79736 129186 79792
rect 129242 79736 129247 79792
rect 128859 79731 128925 79732
rect 129181 79731 129247 79736
rect 129365 79658 129431 79661
rect 128310 79656 129431 79658
rect 128310 79600 129370 79656
rect 129426 79600 129431 79656
rect 128310 79598 129431 79600
rect 129690 79658 129750 79867
rect 130012 79796 130072 79870
rect 130326 79868 130332 79932
rect 130396 79930 130402 79932
rect 130396 79870 130454 79930
rect 130396 79868 130402 79870
rect 130694 79868 130700 79932
rect 130764 79930 130770 79932
rect 131619 79930 131685 79933
rect 132355 79930 132421 79933
rect 130764 79928 131685 79930
rect 130764 79872 131624 79928
rect 131680 79872 131685 79928
rect 130764 79870 131685 79872
rect 130764 79868 130770 79870
rect 131619 79867 131685 79870
rect 131806 79928 132421 79930
rect 131806 79872 132360 79928
rect 132416 79872 132421 79928
rect 132539 79906 132544 79962
rect 132600 79930 132605 79962
rect 134931 79962 134997 79967
rect 133454 79930 133460 79932
rect 132600 79906 133460 79930
rect 132539 79901 133460 79906
rect 131806 79870 132421 79872
rect 132542 79870 133460 79901
rect 131435 79796 131501 79797
rect 129958 79732 129964 79796
rect 130028 79734 130072 79796
rect 130028 79732 130034 79734
rect 131430 79732 131436 79796
rect 131500 79794 131506 79796
rect 131500 79734 131592 79794
rect 131500 79732 131506 79734
rect 131435 79731 131501 79732
rect 129825 79658 129891 79661
rect 129690 79656 129891 79658
rect 129690 79600 129830 79656
rect 129886 79600 129891 79656
rect 129690 79598 129891 79600
rect 127985 79595 128051 79598
rect 129365 79595 129431 79598
rect 129825 79595 129891 79598
rect 131205 79658 131271 79661
rect 131806 79658 131866 79870
rect 132355 79867 132421 79870
rect 133454 79868 133460 79870
rect 133524 79868 133530 79932
rect 134287 79930 134353 79933
rect 134655 79930 134721 79933
rect 133876 79928 134353 79930
rect 133876 79872 134292 79928
rect 134348 79872 134353 79928
rect 133876 79870 134353 79872
rect 133876 79797 133936 79870
rect 134287 79867 134353 79870
rect 134612 79928 134721 79930
rect 134612 79872 134660 79928
rect 134716 79872 134721 79928
rect 134931 79906 134936 79962
rect 134992 79906 134997 79962
rect 134931 79901 134997 79906
rect 135483 79962 135549 79967
rect 135483 79906 135488 79962
rect 135544 79930 135549 79962
rect 135851 79962 135917 79967
rect 135662 79930 135668 79932
rect 135544 79906 135668 79930
rect 135483 79901 135668 79906
rect 134612 79867 134721 79872
rect 133873 79792 133939 79797
rect 133873 79736 133878 79792
rect 133934 79736 133939 79792
rect 133873 79731 133939 79736
rect 131205 79656 131866 79658
rect 131205 79600 131210 79656
rect 131266 79600 131866 79656
rect 131205 79598 131866 79600
rect 134333 79658 134399 79661
rect 134612 79658 134672 79867
rect 134333 79656 134672 79658
rect 134333 79600 134338 79656
rect 134394 79600 134672 79656
rect 134333 79598 134672 79600
rect 134793 79658 134859 79661
rect 134934 79658 134994 79901
rect 135486 79870 135668 79901
rect 135662 79868 135668 79870
rect 135732 79868 135738 79932
rect 135851 79906 135856 79962
rect 135912 79906 135917 79962
rect 136587 79962 136653 79967
rect 136403 79930 136469 79933
rect 136587 79932 136592 79962
rect 136648 79932 136653 79962
rect 136955 79962 137021 79967
rect 136955 79932 136960 79962
rect 137016 79932 137021 79962
rect 137967 79962 138033 79967
rect 135851 79901 135917 79906
rect 136222 79928 136469 79930
rect 135345 79796 135411 79797
rect 135529 79796 135595 79797
rect 135294 79794 135300 79796
rect 135254 79734 135300 79794
rect 135364 79792 135411 79796
rect 135406 79736 135411 79792
rect 135294 79732 135300 79734
rect 135364 79732 135411 79736
rect 135478 79732 135484 79796
rect 135548 79794 135595 79796
rect 135548 79792 135640 79794
rect 135590 79736 135640 79792
rect 135548 79734 135640 79736
rect 135548 79732 135595 79734
rect 135345 79731 135411 79732
rect 135529 79731 135595 79732
rect 134793 79656 134994 79658
rect 134793 79600 134798 79656
rect 134854 79600 134994 79656
rect 134793 79598 134994 79600
rect 135345 79658 135411 79661
rect 135854 79658 135914 79901
rect 135345 79656 135914 79658
rect 135345 79600 135350 79656
rect 135406 79600 135914 79656
rect 135345 79598 135914 79600
rect 136222 79872 136408 79928
rect 136464 79872 136469 79928
rect 136222 79870 136469 79872
rect 136222 79661 136282 79870
rect 136403 79867 136469 79870
rect 136582 79868 136588 79932
rect 136652 79930 136658 79932
rect 136652 79870 136710 79930
rect 136652 79868 136658 79870
rect 136950 79868 136956 79932
rect 137020 79930 137026 79932
rect 137020 79870 137078 79930
rect 137020 79868 137026 79870
rect 137686 79868 137692 79932
rect 137756 79930 137762 79932
rect 137967 79930 137972 79962
rect 137756 79906 137972 79930
rect 138028 79906 138033 79962
rect 137756 79901 138033 79906
rect 138151 79964 138217 79967
rect 139439 79964 139505 79967
rect 138151 79962 138352 79964
rect 138151 79906 138156 79962
rect 138212 79906 138352 79962
rect 139396 79962 139505 79964
rect 138151 79904 138352 79906
rect 138151 79901 138217 79904
rect 137756 79870 138030 79901
rect 137756 79868 137762 79870
rect 138292 79797 138352 79904
rect 138611 79928 138677 79933
rect 138611 79872 138616 79928
rect 138672 79872 138677 79928
rect 138611 79867 138677 79872
rect 138790 79868 138796 79932
rect 138860 79930 138866 79932
rect 139163 79930 139229 79933
rect 138860 79928 139229 79930
rect 138860 79872 139168 79928
rect 139224 79872 139229 79928
rect 138860 79870 139229 79872
rect 138860 79868 138866 79870
rect 139163 79867 139229 79870
rect 139396 79906 139444 79962
rect 139500 79906 139505 79962
rect 139396 79901 139505 79906
rect 140408 79930 140468 80004
rect 146204 79967 146264 80142
rect 156270 80140 156276 80204
rect 156340 80202 156346 80204
rect 156340 80142 162594 80202
rect 156340 80140 156346 80142
rect 157558 80004 157564 80068
rect 157628 80066 157634 80068
rect 157628 80006 157810 80066
rect 157628 80004 157634 80006
rect 140727 79964 140793 79967
rect 140911 79964 140977 79967
rect 140684 79962 140793 79964
rect 140543 79930 140609 79933
rect 140408 79928 140609 79930
rect 136398 79732 136404 79796
rect 136468 79794 136474 79796
rect 138059 79794 138125 79797
rect 136468 79792 138125 79794
rect 136468 79736 138064 79792
rect 138120 79736 138125 79792
rect 136468 79734 138125 79736
rect 136468 79732 136474 79734
rect 138059 79731 138125 79734
rect 138289 79792 138355 79797
rect 138289 79736 138294 79792
rect 138350 79736 138355 79792
rect 138289 79731 138355 79736
rect 136222 79656 136331 79661
rect 136222 79600 136270 79656
rect 136326 79600 136331 79656
rect 136222 79598 136331 79600
rect 138614 79658 138674 79867
rect 138841 79658 138907 79661
rect 138614 79656 138907 79658
rect 138614 79600 138846 79656
rect 138902 79600 138907 79656
rect 138614 79598 138907 79600
rect 131205 79595 131271 79598
rect 134333 79595 134399 79598
rect 134793 79595 134859 79598
rect 135345 79595 135411 79598
rect 136265 79595 136331 79598
rect 138841 79595 138907 79598
rect 139117 79660 139183 79661
rect 139117 79656 139164 79660
rect 139228 79658 139234 79660
rect 139396 79658 139456 79901
rect 140408 79872 140548 79928
rect 140604 79872 140609 79928
rect 140408 79870 140609 79872
rect 140543 79867 140609 79870
rect 140684 79906 140732 79962
rect 140788 79906 140793 79962
rect 140684 79901 140793 79906
rect 140868 79962 140977 79964
rect 140868 79906 140916 79962
rect 140972 79906 140977 79962
rect 141371 79962 141437 79967
rect 142015 79964 142081 79967
rect 141371 79932 141376 79962
rect 141432 79932 141437 79962
rect 141972 79962 142081 79964
rect 141972 79932 142020 79962
rect 140868 79901 140977 79906
rect 139577 79794 139643 79797
rect 139894 79794 139900 79796
rect 139577 79792 139900 79794
rect 139577 79736 139582 79792
rect 139638 79736 139900 79792
rect 139577 79734 139900 79736
rect 139577 79731 139643 79734
rect 139894 79732 139900 79734
rect 139964 79732 139970 79796
rect 139669 79658 139735 79661
rect 139117 79600 139122 79656
rect 139117 79596 139164 79600
rect 139228 79598 139274 79658
rect 139396 79656 139735 79658
rect 139396 79600 139674 79656
rect 139730 79600 139735 79656
rect 139396 79598 139735 79600
rect 139228 79596 139234 79598
rect 139117 79595 139183 79596
rect 139669 79595 139735 79598
rect 140078 79596 140084 79660
rect 140148 79658 140154 79660
rect 140684 79658 140744 79901
rect 140148 79598 140744 79658
rect 140868 79658 140928 79901
rect 141366 79868 141372 79932
rect 141436 79930 141442 79932
rect 141436 79870 141494 79930
rect 141436 79868 141442 79870
rect 141918 79868 141924 79932
rect 141988 79906 142020 79932
rect 142076 79906 142081 79962
rect 143395 79962 143461 79967
rect 142291 79932 142357 79933
rect 142286 79930 142292 79932
rect 141988 79901 142081 79906
rect 141988 79870 142032 79901
rect 142200 79870 142292 79930
rect 141988 79868 141994 79870
rect 142286 79868 142292 79870
rect 142356 79868 142362 79932
rect 142843 79930 142909 79933
rect 142662 79928 142909 79930
rect 142662 79872 142848 79928
rect 142904 79872 142909 79928
rect 142662 79870 142909 79872
rect 142291 79867 142357 79868
rect 140998 79732 141004 79796
rect 141068 79794 141074 79796
rect 142107 79794 142173 79797
rect 141068 79792 142173 79794
rect 141068 79736 142112 79792
rect 142168 79736 142173 79792
rect 141068 79734 142173 79736
rect 141068 79732 141074 79734
rect 142107 79731 142173 79734
rect 142061 79658 142127 79661
rect 140868 79656 142127 79658
rect 140868 79600 142066 79656
rect 142122 79600 142127 79656
rect 140868 79598 142127 79600
rect 142662 79658 142722 79870
rect 142843 79867 142909 79870
rect 143022 79868 143028 79932
rect 143092 79930 143098 79932
rect 143211 79930 143277 79933
rect 143092 79928 143277 79930
rect 143092 79872 143216 79928
rect 143272 79872 143277 79928
rect 143395 79906 143400 79962
rect 143456 79906 143461 79962
rect 143395 79901 143461 79906
rect 143763 79962 143829 79967
rect 143763 79906 143768 79962
rect 143824 79906 143829 79962
rect 144867 79962 144933 79967
rect 143763 79901 143829 79906
rect 143092 79870 143277 79872
rect 143092 79868 143098 79870
rect 143211 79867 143277 79870
rect 142838 79732 142844 79796
rect 142908 79794 142914 79796
rect 142908 79734 143090 79794
rect 142908 79732 142914 79734
rect 142889 79658 142955 79661
rect 142662 79656 142955 79658
rect 142662 79600 142894 79656
rect 142950 79600 142955 79656
rect 142662 79598 142955 79600
rect 143030 79658 143090 79734
rect 143206 79732 143212 79796
rect 143276 79794 143282 79796
rect 143398 79794 143458 79901
rect 143276 79734 143458 79794
rect 143276 79732 143282 79734
rect 143165 79658 143231 79661
rect 143030 79656 143231 79658
rect 143030 79600 143170 79656
rect 143226 79600 143231 79656
rect 143030 79598 143231 79600
rect 140148 79596 140154 79598
rect 142061 79595 142127 79598
rect 142889 79595 142955 79598
rect 143165 79595 143231 79598
rect 143625 79658 143691 79661
rect 143766 79658 143826 79901
rect 144126 79868 144132 79932
rect 144196 79930 144202 79932
rect 144867 79930 144872 79962
rect 144196 79906 144872 79930
rect 144928 79906 144933 79962
rect 144196 79901 144933 79906
rect 145603 79962 145669 79967
rect 145603 79906 145608 79962
rect 145664 79906 145669 79962
rect 145603 79901 145669 79906
rect 146204 79962 146313 79967
rect 146204 79906 146252 79962
rect 146308 79906 146313 79962
rect 147443 79962 147509 79967
rect 146204 79904 146313 79906
rect 146247 79901 146313 79904
rect 144196 79870 144930 79901
rect 144196 79868 144202 79870
rect 144499 79794 144565 79797
rect 144821 79794 144887 79797
rect 144499 79792 144887 79794
rect 144499 79736 144504 79792
rect 144560 79736 144826 79792
rect 144882 79736 144887 79792
rect 144499 79734 144887 79736
rect 144499 79731 144565 79734
rect 144821 79731 144887 79734
rect 143625 79656 143826 79658
rect 143625 79600 143630 79656
rect 143686 79600 143826 79656
rect 143625 79598 143826 79600
rect 144453 79660 144519 79661
rect 144453 79656 144500 79660
rect 144564 79658 144570 79660
rect 145465 79658 145531 79661
rect 145606 79658 145666 79901
rect 147070 79868 147076 79932
rect 147140 79930 147146 79932
rect 147443 79930 147448 79962
rect 147140 79906 147448 79930
rect 147504 79906 147509 79962
rect 148179 79962 148245 79967
rect 148639 79964 148705 79967
rect 147140 79901 147509 79906
rect 147627 79928 147693 79933
rect 147140 79870 147506 79901
rect 147627 79872 147632 79928
rect 147688 79872 147693 79928
rect 148179 79906 148184 79962
rect 148240 79906 148245 79962
rect 148596 79962 148705 79964
rect 148596 79932 148644 79962
rect 148179 79901 148245 79906
rect 147140 79868 147146 79870
rect 147627 79867 147693 79872
rect 145833 79794 145899 79797
rect 147305 79794 147371 79797
rect 145833 79792 147371 79794
rect 145833 79736 145838 79792
rect 145894 79736 147310 79792
rect 147366 79736 147371 79792
rect 145833 79734 147371 79736
rect 145833 79731 145899 79734
rect 147305 79731 147371 79734
rect 144453 79600 144458 79656
rect 143625 79595 143691 79598
rect 144453 79596 144500 79600
rect 144564 79598 144610 79658
rect 145465 79656 145666 79658
rect 145465 79600 145470 79656
rect 145526 79600 145666 79656
rect 145465 79598 145666 79600
rect 144564 79596 144570 79598
rect 144453 79595 144519 79596
rect 145465 79595 145531 79598
rect 145782 79596 145788 79660
rect 145852 79658 145858 79660
rect 146201 79658 146267 79661
rect 145852 79656 146267 79658
rect 145852 79600 146206 79656
rect 146262 79600 146267 79656
rect 145852 79598 146267 79600
rect 145852 79596 145858 79598
rect 146201 79595 146267 79598
rect 146886 79596 146892 79660
rect 146956 79658 146962 79660
rect 147630 79658 147690 79867
rect 147811 79792 147877 79797
rect 147811 79736 147816 79792
rect 147872 79736 147877 79792
rect 147811 79731 147877 79736
rect 146956 79598 147690 79658
rect 147814 79658 147874 79731
rect 148182 79661 148242 79901
rect 148542 79868 148548 79932
rect 148612 79906 148644 79932
rect 148700 79906 148705 79962
rect 149743 79964 149809 79967
rect 150111 79964 150177 79967
rect 149743 79962 149852 79964
rect 148823 79930 148889 79933
rect 149283 79932 149349 79933
rect 149278 79930 149284 79932
rect 148612 79901 148705 79906
rect 148780 79928 148889 79930
rect 148612 79870 148656 79901
rect 148780 79872 148828 79928
rect 148884 79872 148889 79928
rect 148612 79868 148618 79870
rect 148780 79867 148889 79872
rect 149192 79870 149284 79930
rect 149278 79868 149284 79870
rect 149348 79868 149354 79932
rect 149559 79930 149625 79933
rect 149559 79928 149668 79930
rect 149559 79872 149564 79928
rect 149620 79872 149668 79928
rect 149743 79906 149748 79962
rect 149804 79906 149852 79962
rect 150068 79962 150177 79964
rect 150068 79932 150116 79962
rect 149743 79901 149852 79906
rect 149283 79867 149349 79868
rect 149559 79867 149668 79872
rect 148780 79796 148840 79867
rect 148726 79732 148732 79796
rect 148796 79734 148840 79796
rect 148796 79732 148802 79734
rect 147949 79658 148015 79661
rect 147814 79656 148015 79658
rect 147814 79600 147954 79656
rect 148010 79600 148015 79656
rect 147814 79598 148015 79600
rect 146956 79596 146962 79598
rect 147949 79595 148015 79598
rect 148133 79656 148242 79661
rect 148133 79600 148138 79656
rect 148194 79600 148242 79656
rect 148133 79598 148242 79600
rect 149421 79658 149487 79661
rect 149608 79658 149668 79867
rect 149421 79656 149668 79658
rect 149421 79600 149426 79656
rect 149482 79600 149668 79656
rect 149421 79598 149668 79600
rect 149792 79658 149852 79901
rect 150014 79868 150020 79932
rect 150084 79906 150116 79932
rect 150172 79906 150177 79962
rect 150084 79901 150177 79906
rect 150479 79964 150545 79967
rect 150479 79962 150818 79964
rect 150479 79906 150484 79962
rect 150540 79906 150818 79962
rect 151675 79962 151741 79967
rect 150479 79904 150818 79906
rect 150479 79901 150545 79904
rect 150084 79870 150128 79901
rect 150084 79868 150090 79870
rect 150203 79826 150269 79831
rect 150014 79732 150020 79796
rect 150084 79794 150090 79796
rect 150203 79794 150208 79826
rect 150084 79770 150208 79794
rect 150264 79770 150269 79826
rect 150084 79765 150269 79770
rect 150084 79734 150266 79765
rect 150084 79732 150090 79734
rect 150758 79661 150818 79904
rect 151123 79928 151189 79933
rect 151123 79872 151128 79928
rect 151184 79872 151189 79928
rect 151123 79867 151189 79872
rect 151486 79868 151492 79932
rect 151556 79930 151562 79932
rect 151675 79930 151680 79962
rect 151556 79906 151680 79930
rect 151736 79906 151741 79962
rect 152779 79962 152845 79967
rect 153055 79964 153121 79967
rect 152043 79932 152109 79933
rect 151556 79901 151741 79906
rect 151556 79870 151738 79901
rect 151556 79868 151562 79870
rect 152038 79868 152044 79932
rect 152108 79930 152114 79932
rect 152108 79870 152200 79930
rect 152411 79928 152477 79933
rect 152779 79932 152784 79962
rect 152840 79932 152845 79962
rect 153012 79962 153121 79964
rect 152411 79872 152416 79928
rect 152472 79872 152477 79928
rect 152108 79868 152114 79870
rect 152043 79867 152109 79868
rect 152411 79867 152477 79872
rect 152774 79868 152780 79932
rect 152844 79930 152850 79932
rect 152844 79870 152902 79930
rect 153012 79906 153060 79962
rect 153116 79906 153121 79962
rect 153699 79962 153765 79967
rect 153012 79901 153121 79906
rect 152844 79868 152850 79870
rect 150065 79658 150131 79661
rect 149792 79656 150131 79658
rect 149792 79600 150070 79656
rect 150126 79600 150131 79656
rect 149792 79598 150131 79600
rect 148133 79595 148199 79598
rect 149421 79595 149487 79598
rect 150065 79595 150131 79598
rect 150709 79656 150818 79661
rect 150709 79600 150714 79656
rect 150770 79600 150818 79656
rect 150709 79598 150818 79600
rect 151126 79661 151186 79867
rect 151767 79794 151833 79797
rect 151632 79792 151833 79794
rect 151632 79736 151772 79792
rect 151828 79736 151833 79792
rect 151632 79734 151833 79736
rect 151126 79656 151235 79661
rect 151126 79600 151174 79656
rect 151230 79600 151235 79656
rect 151126 79598 151235 79600
rect 151632 79660 151692 79734
rect 151767 79731 151833 79734
rect 151632 79598 151676 79660
rect 150709 79595 150775 79598
rect 151169 79595 151235 79598
rect 151670 79596 151676 79598
rect 151740 79596 151746 79660
rect 151813 79658 151879 79661
rect 152414 79658 152474 79867
rect 153012 79796 153072 79901
rect 153326 79868 153332 79932
rect 153396 79930 153402 79932
rect 153699 79930 153704 79962
rect 153396 79906 153704 79930
rect 153760 79906 153765 79962
rect 153883 79962 153949 79967
rect 153883 79932 153888 79962
rect 153944 79932 153949 79962
rect 154803 79962 154869 79967
rect 153396 79901 153765 79906
rect 153396 79870 153762 79901
rect 153396 79868 153402 79870
rect 153878 79868 153884 79932
rect 153948 79930 153954 79932
rect 154159 79930 154225 79933
rect 153948 79870 154006 79930
rect 154116 79928 154225 79930
rect 154116 79872 154164 79928
rect 154220 79872 154225 79928
rect 153948 79868 153954 79870
rect 154116 79867 154225 79872
rect 154343 79930 154409 79933
rect 154343 79928 154452 79930
rect 154343 79872 154348 79928
rect 154404 79872 154452 79928
rect 154803 79906 154808 79962
rect 154864 79906 154869 79962
rect 154803 79901 154869 79906
rect 154987 79962 155053 79967
rect 154987 79906 154992 79962
rect 155048 79906 155053 79962
rect 154987 79901 155053 79906
rect 155631 79964 155697 79967
rect 155631 79962 155740 79964
rect 155631 79906 155636 79962
rect 155692 79932 155740 79962
rect 156459 79962 156525 79967
rect 156091 79932 156157 79933
rect 156459 79932 156464 79962
rect 156520 79932 156525 79962
rect 157103 79964 157169 79967
rect 157103 79962 157212 79964
rect 155692 79906 155724 79932
rect 155631 79901 155724 79906
rect 154343 79867 154452 79872
rect 154116 79796 154176 79867
rect 152958 79732 152964 79796
rect 153028 79734 153072 79796
rect 153028 79732 153034 79734
rect 154062 79732 154068 79796
rect 154132 79734 154176 79796
rect 154392 79796 154452 79867
rect 154392 79734 154436 79796
rect 154132 79732 154138 79734
rect 154430 79732 154436 79734
rect 154500 79732 154506 79796
rect 154806 79661 154866 79901
rect 154990 79797 155050 79901
rect 155680 79870 155724 79901
rect 155718 79868 155724 79870
rect 155788 79868 155794 79932
rect 156086 79930 156092 79932
rect 156000 79870 156092 79930
rect 156086 79868 156092 79870
rect 156156 79868 156162 79932
rect 156454 79868 156460 79932
rect 156524 79930 156530 79932
rect 156524 79870 156582 79930
rect 156643 79928 156709 79933
rect 156643 79872 156648 79928
rect 156704 79872 156709 79928
rect 156524 79868 156530 79870
rect 156091 79867 156157 79868
rect 156643 79867 156709 79872
rect 156919 79930 156985 79933
rect 156919 79928 157028 79930
rect 156919 79872 156924 79928
rect 156980 79872 157028 79928
rect 157103 79906 157108 79962
rect 157164 79932 157212 79962
rect 157750 79933 157810 80006
rect 158846 80004 158852 80068
rect 158916 80066 158922 80068
rect 158916 80006 160018 80066
rect 158916 80004 158922 80006
rect 159958 79933 160018 80006
rect 162534 79967 162594 80142
rect 166574 80140 166580 80204
rect 166644 80202 166650 80204
rect 166644 80142 167010 80202
rect 166644 80140 166650 80142
rect 166950 79967 167010 80142
rect 168698 79967 168758 80278
rect 554773 80275 554839 80278
rect 171734 80142 182190 80202
rect 171734 79967 171794 80142
rect 173198 80066 173204 80068
rect 173068 80006 173204 80066
rect 160691 79962 160757 79967
rect 157164 79906 157196 79932
rect 157103 79901 157196 79906
rect 156919 79867 157028 79872
rect 157152 79870 157196 79901
rect 157190 79868 157196 79870
rect 157260 79868 157266 79932
rect 157747 79928 157813 79933
rect 157747 79872 157752 79928
rect 157808 79872 157813 79928
rect 157747 79867 157813 79872
rect 158207 79930 158273 79933
rect 158943 79930 159009 79933
rect 159771 79932 159837 79933
rect 159766 79930 159772 79932
rect 158207 79928 158408 79930
rect 158207 79872 158212 79928
rect 158268 79872 158408 79928
rect 158943 79928 159328 79930
rect 158207 79870 158408 79872
rect 158207 79867 158273 79870
rect 154941 79792 155050 79797
rect 154941 79736 154946 79792
rect 155002 79736 155050 79792
rect 154941 79734 155050 79736
rect 155677 79794 155743 79797
rect 155902 79794 155908 79796
rect 155677 79792 155908 79794
rect 155677 79736 155682 79792
rect 155738 79736 155908 79792
rect 155677 79734 155908 79736
rect 154941 79731 155007 79734
rect 155677 79731 155743 79734
rect 155902 79732 155908 79734
rect 155972 79732 155978 79796
rect 153929 79660 153995 79661
rect 151813 79656 152474 79658
rect 151813 79600 151818 79656
rect 151874 79600 152474 79656
rect 151813 79598 152474 79600
rect 151813 79595 151879 79598
rect 153878 79596 153884 79660
rect 153948 79658 153995 79660
rect 154205 79660 154271 79661
rect 153948 79656 154040 79658
rect 153990 79600 154040 79656
rect 153948 79598 154040 79600
rect 154205 79656 154252 79660
rect 154316 79658 154322 79660
rect 154205 79600 154210 79656
rect 153948 79596 153995 79598
rect 153929 79595 153995 79596
rect 154205 79596 154252 79600
rect 154316 79598 154362 79658
rect 154757 79656 154866 79661
rect 154757 79600 154762 79656
rect 154818 79600 154866 79656
rect 154757 79598 154866 79600
rect 156646 79658 156706 79867
rect 156968 79796 157028 79867
rect 156968 79734 157012 79796
rect 157006 79732 157012 79734
rect 157076 79732 157082 79796
rect 157425 79794 157491 79797
rect 157793 79794 157859 79797
rect 157931 79796 157997 79797
rect 158348 79796 158408 79870
rect 158483 79894 158549 79899
rect 158483 79838 158488 79894
rect 158544 79838 158549 79894
rect 158943 79872 158948 79928
rect 159004 79872 159328 79928
rect 158943 79870 159328 79872
rect 159680 79870 159772 79930
rect 158943 79867 159009 79870
rect 158483 79833 158549 79838
rect 157425 79792 157859 79794
rect 157425 79736 157430 79792
rect 157486 79736 157798 79792
rect 157854 79736 157859 79792
rect 157425 79734 157859 79736
rect 157425 79731 157491 79734
rect 157793 79731 157859 79734
rect 157926 79732 157932 79796
rect 157996 79794 158002 79796
rect 157996 79734 158088 79794
rect 157996 79732 158002 79734
rect 158294 79732 158300 79796
rect 158364 79734 158408 79796
rect 158364 79732 158370 79734
rect 157931 79731 157997 79732
rect 156781 79658 156847 79661
rect 156646 79656 156847 79658
rect 156646 79600 156786 79656
rect 156842 79600 156847 79656
rect 156646 79598 156847 79600
rect 154316 79596 154322 79598
rect 154205 79595 154271 79596
rect 154757 79595 154823 79598
rect 156781 79595 156847 79598
rect 158110 79596 158116 79660
rect 158180 79658 158186 79660
rect 158486 79658 158546 79833
rect 159268 79797 159328 79870
rect 159766 79868 159772 79870
rect 159836 79868 159842 79932
rect 159955 79928 160021 79933
rect 160691 79930 160696 79962
rect 159955 79872 159960 79928
rect 160016 79872 160021 79928
rect 159771 79867 159837 79868
rect 159955 79867 160021 79872
rect 160510 79906 160696 79930
rect 160752 79906 160757 79962
rect 161059 79962 161125 79967
rect 160510 79901 160757 79906
rect 160510 79870 160754 79901
rect 159403 79828 159469 79831
rect 159403 79826 159526 79828
rect 159265 79792 159331 79797
rect 159403 79796 159408 79826
rect 159464 79796 159526 79826
rect 159265 79736 159270 79792
rect 159326 79736 159331 79792
rect 159265 79731 159331 79736
rect 159398 79732 159404 79796
rect 159468 79768 159526 79796
rect 159863 79794 159929 79797
rect 160134 79794 160140 79796
rect 159863 79792 160140 79794
rect 159468 79732 159474 79768
rect 159863 79736 159868 79792
rect 159924 79736 160140 79792
rect 159863 79734 160140 79736
rect 159863 79731 159929 79734
rect 160134 79732 160140 79734
rect 160204 79732 160210 79796
rect 158180 79598 158546 79658
rect 158180 79596 158186 79598
rect 159030 79596 159036 79660
rect 159100 79658 159106 79660
rect 160001 79658 160067 79661
rect 159100 79656 160067 79658
rect 159100 79600 160006 79656
rect 160062 79600 160067 79656
rect 159100 79598 160067 79600
rect 160510 79658 160570 79870
rect 160870 79868 160876 79932
rect 160940 79930 160946 79932
rect 161059 79930 161064 79962
rect 160940 79906 161064 79930
rect 161120 79906 161125 79962
rect 161427 79964 161493 79967
rect 161427 79962 161550 79964
rect 161427 79932 161432 79962
rect 161488 79932 161550 79962
rect 160940 79901 161125 79906
rect 160940 79870 161122 79901
rect 160940 79868 160946 79870
rect 161422 79868 161428 79932
rect 161492 79904 161550 79932
rect 161611 79962 161677 79967
rect 161611 79906 161616 79962
rect 161672 79906 161677 79962
rect 162163 79962 162229 79967
rect 161795 79932 161861 79933
rect 161492 79868 161498 79904
rect 161611 79901 161677 79906
rect 160686 79732 160692 79796
rect 160756 79794 160762 79796
rect 160875 79794 160941 79797
rect 160756 79792 160941 79794
rect 160756 79736 160880 79792
rect 160936 79736 160941 79792
rect 160756 79734 160941 79736
rect 160756 79732 160762 79734
rect 160875 79731 160941 79734
rect 160645 79658 160711 79661
rect 160510 79656 160711 79658
rect 160510 79600 160650 79656
rect 160706 79600 160711 79656
rect 160510 79598 160711 79600
rect 161614 79658 161674 79901
rect 161790 79868 161796 79932
rect 161860 79930 161866 79932
rect 161860 79870 161952 79930
rect 162163 79906 162168 79962
rect 162224 79906 162229 79962
rect 162163 79901 162229 79906
rect 162531 79962 162597 79967
rect 162531 79906 162536 79962
rect 162592 79906 162597 79962
rect 162715 79962 162781 79967
rect 162715 79932 162720 79962
rect 162776 79932 162781 79962
rect 166671 79964 166737 79967
rect 166671 79962 166780 79964
rect 162531 79901 162597 79906
rect 161860 79868 161866 79870
rect 161795 79867 161861 79868
rect 161974 79732 161980 79796
rect 162044 79794 162050 79796
rect 162166 79794 162226 79901
rect 162710 79868 162716 79932
rect 162780 79930 162786 79932
rect 162780 79870 162838 79930
rect 163267 79928 163333 79933
rect 163267 79872 163272 79928
rect 163328 79872 163333 79928
rect 162780 79868 162786 79870
rect 163267 79867 163333 79872
rect 163635 79928 163701 79933
rect 163635 79872 163640 79928
rect 163696 79872 163701 79928
rect 163635 79867 163701 79872
rect 163819 79928 163885 79933
rect 163819 79872 163824 79928
rect 163880 79872 163885 79928
rect 165107 79930 165173 79933
rect 165470 79930 165476 79932
rect 165107 79928 165476 79930
rect 163819 79867 163885 79872
rect 164555 79894 164621 79899
rect 162044 79734 162226 79794
rect 162044 79732 162050 79734
rect 163270 79661 163330 79867
rect 163638 79797 163698 79867
rect 163589 79792 163698 79797
rect 163589 79736 163594 79792
rect 163650 79736 163698 79792
rect 163589 79734 163698 79736
rect 163589 79731 163655 79734
rect 163822 79661 163882 79867
rect 164555 79838 164560 79894
rect 164616 79838 164621 79894
rect 165107 79872 165112 79928
rect 165168 79872 165476 79928
rect 165107 79870 165476 79872
rect 165107 79867 165173 79870
rect 165470 79868 165476 79870
rect 165540 79868 165546 79932
rect 165935 79930 166001 79933
rect 166206 79930 166212 79932
rect 165935 79928 166212 79930
rect 165935 79872 165940 79928
rect 165996 79872 166212 79928
rect 165935 79870 166212 79872
rect 165935 79867 166001 79870
rect 166206 79868 166212 79870
rect 166276 79868 166282 79932
rect 166395 79928 166461 79933
rect 166395 79872 166400 79928
rect 166456 79872 166461 79928
rect 166671 79906 166676 79962
rect 166732 79932 166780 79962
rect 166947 79962 167013 79967
rect 166732 79906 166764 79932
rect 166671 79901 166764 79906
rect 166395 79867 166461 79872
rect 166720 79870 166764 79901
rect 166758 79868 166764 79870
rect 166828 79868 166834 79932
rect 166947 79906 166952 79962
rect 167008 79906 167013 79962
rect 168695 79962 168761 79967
rect 167223 79930 167289 79933
rect 166947 79901 167013 79906
rect 167180 79928 167289 79930
rect 167180 79872 167228 79928
rect 167284 79872 167289 79928
rect 167180 79867 167289 79872
rect 167591 79930 167657 79933
rect 168046 79930 168052 79932
rect 167591 79928 168052 79930
rect 167591 79872 167596 79928
rect 167652 79872 168052 79928
rect 167591 79870 168052 79872
rect 167591 79867 167657 79870
rect 168046 79868 168052 79870
rect 168116 79868 168122 79932
rect 168327 79928 168393 79933
rect 168327 79872 168332 79928
rect 168388 79872 168393 79928
rect 168695 79906 168700 79962
rect 168756 79906 168761 79962
rect 169707 79962 169773 79967
rect 170351 79964 170417 79967
rect 168695 79901 168761 79906
rect 168327 79867 168393 79872
rect 169150 79868 169156 79932
rect 169220 79930 169226 79932
rect 169431 79930 169497 79933
rect 169220 79928 169497 79930
rect 169220 79872 169436 79928
rect 169492 79872 169497 79928
rect 169707 79906 169712 79962
rect 169768 79906 169773 79962
rect 170308 79962 170417 79964
rect 170075 79932 170141 79933
rect 170070 79930 170076 79932
rect 169707 79901 169773 79906
rect 169220 79870 169497 79872
rect 169220 79868 169226 79870
rect 169431 79867 169497 79870
rect 164555 79833 164621 79838
rect 161841 79658 161907 79661
rect 161614 79656 161907 79658
rect 161614 79600 161846 79656
rect 161902 79600 161907 79656
rect 161614 79598 161907 79600
rect 159100 79596 159106 79598
rect 160001 79595 160067 79598
rect 160645 79595 160711 79598
rect 161841 79595 161907 79598
rect 162158 79596 162164 79660
rect 162228 79658 162234 79660
rect 162301 79658 162367 79661
rect 162228 79656 162367 79658
rect 162228 79600 162306 79656
rect 162362 79600 162367 79656
rect 162228 79598 162367 79600
rect 162228 79596 162234 79598
rect 162301 79595 162367 79598
rect 162577 79658 162643 79661
rect 162710 79658 162716 79660
rect 162577 79656 162716 79658
rect 162577 79600 162582 79656
rect 162638 79600 162716 79656
rect 162577 79598 162716 79600
rect 162577 79595 162643 79598
rect 162710 79596 162716 79598
rect 162780 79596 162786 79660
rect 163270 79656 163379 79661
rect 163270 79600 163318 79656
rect 163374 79600 163379 79656
rect 163270 79598 163379 79600
rect 163313 79595 163379 79598
rect 163773 79656 163882 79661
rect 163773 79600 163778 79656
rect 163834 79600 163882 79656
rect 163773 79598 163882 79600
rect 164558 79658 164618 79833
rect 165705 79794 165771 79797
rect 166398 79794 166458 79867
rect 165705 79792 166458 79794
rect 165705 79736 165710 79792
rect 165766 79736 166458 79792
rect 165705 79734 166458 79736
rect 166579 79792 166645 79797
rect 166579 79736 166584 79792
rect 166640 79736 166645 79792
rect 165705 79731 165771 79734
rect 166579 79731 166645 79736
rect 167180 79794 167240 79867
rect 167310 79794 167316 79796
rect 167180 79734 167316 79794
rect 167310 79732 167316 79734
rect 167380 79732 167386 79796
rect 167678 79732 167684 79796
rect 167748 79794 167754 79796
rect 168143 79794 168209 79797
rect 167748 79792 168209 79794
rect 167748 79736 168148 79792
rect 168204 79736 168209 79792
rect 167748 79734 168209 79736
rect 167748 79732 167754 79734
rect 168143 79731 168209 79734
rect 165061 79658 165127 79661
rect 164558 79656 165127 79658
rect 164558 79600 165066 79656
rect 165122 79600 165127 79656
rect 164558 79598 165127 79600
rect 163773 79595 163839 79598
rect 165061 79595 165127 79598
rect 165286 79596 165292 79660
rect 165356 79658 165362 79660
rect 165429 79658 165495 79661
rect 165356 79656 165495 79658
rect 165356 79600 165434 79656
rect 165490 79600 165495 79656
rect 165356 79598 165495 79600
rect 165356 79596 165362 79598
rect 165429 79595 165495 79598
rect 166022 79596 166028 79660
rect 166092 79658 166098 79660
rect 166582 79658 166642 79731
rect 166092 79598 166642 79658
rect 168330 79658 168390 79867
rect 169518 79732 169524 79796
rect 169588 79794 169594 79796
rect 169710 79794 169770 79901
rect 169984 79870 170076 79930
rect 170070 79868 170076 79870
rect 170140 79868 170146 79932
rect 170308 79906 170356 79962
rect 170412 79930 170417 79962
rect 171731 79962 171797 79967
rect 170995 79932 171061 79933
rect 170622 79930 170628 79932
rect 170412 79906 170628 79930
rect 170308 79870 170628 79906
rect 170622 79868 170628 79870
rect 170692 79868 170698 79932
rect 170990 79868 170996 79932
rect 171060 79930 171066 79932
rect 171271 79930 171337 79933
rect 171542 79930 171548 79932
rect 171060 79870 171152 79930
rect 171271 79928 171548 79930
rect 171271 79872 171276 79928
rect 171332 79872 171548 79928
rect 171271 79870 171548 79872
rect 171060 79868 171066 79870
rect 170075 79867 170141 79868
rect 170995 79867 171061 79868
rect 171271 79867 171337 79870
rect 171542 79868 171548 79870
rect 171612 79868 171618 79932
rect 171731 79906 171736 79962
rect 171792 79906 171797 79962
rect 171731 79901 171797 79906
rect 172191 79964 172257 79967
rect 172191 79962 172300 79964
rect 172191 79906 172196 79962
rect 172252 79930 172300 79962
rect 172646 79930 172652 79932
rect 172252 79906 172652 79930
rect 172191 79901 172652 79906
rect 172240 79870 172652 79901
rect 172646 79868 172652 79870
rect 172716 79868 172722 79932
rect 172835 79930 172901 79933
rect 173068 79930 173128 80006
rect 173198 80004 173204 80006
rect 173268 80004 173274 80068
rect 173566 80004 173572 80068
rect 173636 80066 173642 80068
rect 176101 80066 176167 80069
rect 173636 80064 176167 80066
rect 173636 80008 176106 80064
rect 176162 80008 176167 80064
rect 173636 80006 176167 80008
rect 173636 80004 173642 80006
rect 176101 80003 176167 80006
rect 173387 79962 173453 79967
rect 172835 79928 173128 79930
rect 172835 79872 172840 79928
rect 172896 79872 173128 79928
rect 172835 79870 173128 79872
rect 173203 79928 173269 79933
rect 173203 79872 173208 79928
rect 173264 79872 173269 79928
rect 173387 79906 173392 79962
rect 173448 79906 173453 79962
rect 173387 79901 173453 79906
rect 172835 79867 172901 79870
rect 173203 79867 173269 79872
rect 169588 79734 169770 79794
rect 169588 79732 169594 79734
rect 170438 79732 170444 79796
rect 170508 79794 170514 79796
rect 170903 79794 170969 79797
rect 173206 79794 173266 79867
rect 173390 79797 173450 79901
rect 170508 79792 170969 79794
rect 170508 79736 170908 79792
rect 170964 79736 170969 79792
rect 170508 79734 170969 79736
rect 170508 79732 170514 79734
rect 170903 79731 170969 79734
rect 171090 79734 173266 79794
rect 173341 79792 173450 79797
rect 173341 79736 173346 79792
rect 173402 79736 173450 79792
rect 173341 79734 173450 79736
rect 182130 79794 182190 80142
rect 580441 79794 580507 79797
rect 182130 79792 580507 79794
rect 182130 79736 580446 79792
rect 580502 79736 580507 79792
rect 182130 79734 580507 79736
rect 168966 79658 168972 79660
rect 168330 79598 168972 79658
rect 166092 79596 166098 79598
rect 168966 79596 168972 79598
rect 169036 79596 169042 79660
rect 170029 79658 170095 79661
rect 171090 79658 171150 79734
rect 173341 79731 173407 79734
rect 580441 79731 580507 79734
rect 170029 79656 171150 79658
rect 170029 79600 170034 79656
rect 170090 79600 171150 79656
rect 170029 79598 171150 79600
rect 171869 79660 171935 79661
rect 171869 79656 171916 79660
rect 171980 79658 171986 79660
rect 171869 79600 171874 79656
rect 170029 79595 170095 79598
rect 171869 79596 171916 79600
rect 171980 79598 172026 79658
rect 171980 79596 171986 79598
rect 172094 79596 172100 79660
rect 172164 79658 172170 79660
rect 174997 79658 175063 79661
rect 172164 79656 175063 79658
rect 172164 79600 175002 79656
rect 175058 79600 175063 79656
rect 172164 79598 175063 79600
rect 172164 79596 172170 79598
rect 171869 79595 171935 79596
rect 174997 79595 175063 79598
rect 3969 79522 4035 79525
rect 162669 79522 162735 79525
rect 173157 79522 173223 79525
rect 3969 79520 162594 79522
rect 3969 79464 3974 79520
rect 4030 79464 162594 79520
rect 3969 79462 162594 79464
rect 3969 79459 4035 79462
rect 3785 79386 3851 79389
rect 162534 79386 162594 79462
rect 162669 79520 173223 79522
rect 162669 79464 162674 79520
rect 162730 79464 173162 79520
rect 173218 79464 173223 79520
rect 162669 79462 173223 79464
rect 162669 79459 162735 79462
rect 173157 79459 173223 79462
rect 173341 79386 173407 79389
rect 580257 79386 580323 79389
rect 3785 79384 162410 79386
rect 3785 79328 3790 79384
rect 3846 79328 162410 79384
rect 3785 79326 162410 79328
rect 162534 79384 173407 79386
rect 162534 79328 173346 79384
rect 173402 79328 173407 79384
rect 162534 79326 173407 79328
rect 3785 79323 3851 79326
rect 3601 79250 3667 79253
rect 162350 79250 162410 79326
rect 173341 79323 173407 79326
rect 180750 79384 580323 79386
rect 180750 79328 580262 79384
rect 580318 79328 580323 79384
rect 180750 79326 580323 79328
rect 173249 79250 173315 79253
rect 3601 79248 162272 79250
rect 3601 79192 3606 79248
rect 3662 79192 162272 79248
rect 3601 79190 162272 79192
rect 162350 79248 173315 79250
rect 162350 79192 173254 79248
rect 173310 79192 173315 79248
rect 162350 79190 173315 79192
rect 3601 79187 3667 79190
rect 3417 79114 3483 79117
rect 162212 79114 162272 79190
rect 173249 79187 173315 79190
rect 173382 79188 173388 79252
rect 173452 79250 173458 79252
rect 180750 79250 180810 79326
rect 580257 79323 580323 79326
rect 173452 79190 180810 79250
rect 173452 79188 173458 79190
rect 170029 79114 170095 79117
rect 170949 79116 171015 79117
rect 170949 79114 170996 79116
rect 3417 79112 162042 79114
rect 3417 79056 3422 79112
rect 3478 79056 162042 79112
rect 3417 79054 162042 79056
rect 162212 79112 170095 79114
rect 162212 79056 170034 79112
rect 170090 79056 170095 79112
rect 162212 79054 170095 79056
rect 170904 79112 170996 79114
rect 170904 79056 170954 79112
rect 170904 79054 170996 79056
rect 3417 79051 3483 79054
rect 3233 78978 3299 78981
rect 161473 78978 161539 78981
rect 3233 78976 161539 78978
rect 3233 78920 3238 78976
rect 3294 78920 161478 78976
rect 161534 78920 161539 78976
rect 3233 78918 161539 78920
rect 161982 78978 162042 79054
rect 170029 79051 170095 79054
rect 170949 79052 170996 79054
rect 171060 79052 171066 79116
rect 171501 79114 171567 79117
rect 176193 79114 176259 79117
rect 171501 79112 176259 79114
rect 171501 79056 171506 79112
rect 171562 79056 176198 79112
rect 176254 79056 176259 79112
rect 171501 79054 176259 79056
rect 170949 79051 171015 79052
rect 171501 79051 171567 79054
rect 176193 79051 176259 79054
rect 170857 78978 170923 78981
rect 173709 78978 173775 78981
rect 161982 78918 170506 78978
rect 3233 78915 3299 78918
rect 161473 78915 161539 78918
rect 3049 78842 3115 78845
rect 169661 78844 169727 78845
rect 3049 78840 169218 78842
rect 3049 78784 3054 78840
rect 3110 78784 169218 78840
rect 3049 78782 169218 78784
rect 3049 78779 3115 78782
rect 125685 78708 125751 78709
rect 125869 78708 125935 78709
rect 125685 78706 125732 78708
rect 125640 78704 125732 78706
rect 125640 78648 125690 78704
rect 125640 78646 125732 78648
rect 125685 78644 125732 78646
rect 125796 78644 125802 78708
rect 125869 78704 125916 78708
rect 125980 78706 125986 78708
rect 126145 78706 126211 78709
rect 126278 78706 126284 78708
rect 125869 78648 125874 78704
rect 125869 78644 125916 78648
rect 125980 78646 126026 78706
rect 126145 78704 126284 78706
rect 126145 78648 126150 78704
rect 126206 78648 126284 78704
rect 126145 78646 126284 78648
rect 125980 78644 125986 78646
rect 125685 78643 125751 78644
rect 125869 78643 125935 78644
rect 126145 78643 126211 78646
rect 126278 78644 126284 78646
rect 126348 78644 126354 78708
rect 126421 78706 126487 78709
rect 156689 78708 156755 78709
rect 126646 78706 126652 78708
rect 126421 78704 126652 78706
rect 126421 78648 126426 78704
rect 126482 78648 126652 78704
rect 126421 78646 126652 78648
rect 126421 78643 126487 78646
rect 126646 78644 126652 78646
rect 126716 78644 126722 78708
rect 127566 78644 127572 78708
rect 127636 78706 127642 78708
rect 156270 78706 156276 78708
rect 127636 78646 156276 78706
rect 127636 78644 127642 78646
rect 156270 78644 156276 78646
rect 156340 78644 156346 78708
rect 156638 78644 156644 78708
rect 156708 78706 156755 78708
rect 157149 78706 157215 78709
rect 157374 78706 157380 78708
rect 156708 78704 156800 78706
rect 156750 78648 156800 78704
rect 156708 78646 156800 78648
rect 157149 78704 157380 78706
rect 157149 78648 157154 78704
rect 157210 78648 157380 78704
rect 157149 78646 157380 78648
rect 156708 78644 156755 78646
rect 156689 78643 156755 78644
rect 157149 78643 157215 78646
rect 157374 78644 157380 78646
rect 157444 78644 157450 78708
rect 161565 78706 161631 78709
rect 168373 78706 168439 78709
rect 161565 78704 168439 78706
rect 161565 78648 161570 78704
rect 161626 78648 168378 78704
rect 168434 78648 168439 78704
rect 161565 78646 168439 78648
rect 169158 78706 169218 78782
rect 169661 78840 169708 78844
rect 169772 78842 169778 78844
rect 170446 78842 170506 78918
rect 170857 78976 173775 78978
rect 170857 78920 170862 78976
rect 170918 78920 173714 78976
rect 173770 78920 173775 78976
rect 170857 78918 173775 78920
rect 170857 78915 170923 78918
rect 173709 78915 173775 78918
rect 173433 78842 173499 78845
rect 169661 78784 169666 78840
rect 169661 78780 169708 78784
rect 169772 78782 169818 78842
rect 170446 78840 173499 78842
rect 170446 78784 173438 78840
rect 173494 78784 173499 78840
rect 170446 78782 173499 78784
rect 169772 78780 169778 78782
rect 169661 78779 169727 78780
rect 173433 78779 173499 78782
rect 173617 78706 173683 78709
rect 169158 78704 173683 78706
rect 169158 78648 173622 78704
rect 173678 78648 173683 78704
rect 169158 78646 173683 78648
rect 161565 78643 161631 78646
rect 168373 78643 168439 78646
rect 173617 78643 173683 78646
rect 119337 78570 119403 78573
rect 173893 78570 173959 78573
rect 119337 78568 173959 78570
rect 119337 78512 119342 78568
rect 119398 78512 173898 78568
rect 173954 78512 173959 78568
rect 119337 78510 173959 78512
rect 119337 78507 119403 78510
rect 173893 78507 173959 78510
rect 127985 78436 128051 78437
rect 128721 78436 128787 78437
rect 127934 78372 127940 78436
rect 128004 78434 128051 78436
rect 128004 78432 128096 78434
rect 128046 78376 128096 78432
rect 128004 78374 128096 78376
rect 128004 78372 128051 78374
rect 128670 78372 128676 78436
rect 128740 78434 128787 78436
rect 129365 78436 129431 78437
rect 129733 78436 129799 78437
rect 129365 78434 129412 78436
rect 128740 78432 128832 78434
rect 128782 78376 128832 78432
rect 128740 78374 128832 78376
rect 129320 78432 129412 78434
rect 129320 78376 129370 78432
rect 129320 78374 129412 78376
rect 128740 78372 128787 78374
rect 127985 78371 128051 78372
rect 128721 78371 128787 78372
rect 129365 78372 129412 78374
rect 129476 78372 129482 78436
rect 129733 78432 129780 78436
rect 129844 78434 129850 78436
rect 130193 78434 130259 78437
rect 130326 78434 130332 78436
rect 129733 78376 129738 78432
rect 129733 78372 129780 78376
rect 129844 78374 129890 78434
rect 130193 78432 130332 78434
rect 130193 78376 130198 78432
rect 130254 78376 130332 78432
rect 130193 78374 130332 78376
rect 129844 78372 129850 78374
rect 129365 78371 129431 78372
rect 129733 78371 129799 78372
rect 130193 78371 130259 78374
rect 130326 78372 130332 78374
rect 130396 78372 130402 78436
rect 131113 78434 131179 78437
rect 135529 78436 135595 78437
rect 131614 78434 131620 78436
rect 131113 78432 131620 78434
rect 131113 78376 131118 78432
rect 131174 78376 131620 78432
rect 131113 78374 131620 78376
rect 131113 78371 131179 78374
rect 131614 78372 131620 78374
rect 131684 78372 131690 78436
rect 135478 78372 135484 78436
rect 135548 78434 135595 78436
rect 136541 78436 136607 78437
rect 137921 78436 137987 78437
rect 136541 78434 136588 78436
rect 135548 78432 135640 78434
rect 135590 78376 135640 78432
rect 135548 78374 135640 78376
rect 136496 78432 136588 78434
rect 136496 78376 136546 78432
rect 136496 78374 136588 78376
rect 135548 78372 135595 78374
rect 135529 78371 135595 78372
rect 136541 78372 136588 78374
rect 136652 78372 136658 78436
rect 137870 78434 137876 78436
rect 137830 78374 137876 78434
rect 137940 78432 137987 78436
rect 137982 78376 137987 78432
rect 137870 78372 137876 78374
rect 137940 78372 137987 78376
rect 138974 78372 138980 78436
rect 139044 78434 139050 78436
rect 139393 78434 139459 78437
rect 139044 78432 139459 78434
rect 139044 78376 139398 78432
rect 139454 78376 139459 78432
rect 139044 78374 139459 78376
rect 139044 78372 139050 78374
rect 136541 78371 136607 78372
rect 137921 78371 137987 78372
rect 139393 78371 139459 78374
rect 143349 78436 143415 78437
rect 144637 78436 144703 78437
rect 143349 78432 143396 78436
rect 143460 78434 143466 78436
rect 143349 78376 143354 78432
rect 143349 78372 143396 78376
rect 143460 78374 143506 78434
rect 144637 78432 144684 78436
rect 144748 78434 144754 78436
rect 144637 78376 144642 78432
rect 143460 78372 143466 78374
rect 144637 78372 144684 78376
rect 144748 78374 144794 78434
rect 144748 78372 144754 78374
rect 147254 78372 147260 78436
rect 147324 78434 147330 78436
rect 147581 78434 147647 78437
rect 147324 78432 147647 78434
rect 147324 78376 147586 78432
rect 147642 78376 147647 78432
rect 147324 78374 147647 78376
rect 147324 78372 147330 78374
rect 143349 78371 143415 78372
rect 144637 78371 144703 78372
rect 147581 78371 147647 78374
rect 147949 78434 148015 78437
rect 148358 78434 148364 78436
rect 147949 78432 148364 78434
rect 147949 78376 147954 78432
rect 148010 78376 148364 78432
rect 147949 78374 148364 78376
rect 147949 78371 148015 78374
rect 148358 78372 148364 78374
rect 148428 78372 148434 78436
rect 149278 78372 149284 78436
rect 149348 78434 149354 78436
rect 149605 78434 149671 78437
rect 149348 78432 149671 78434
rect 149348 78376 149610 78432
rect 149666 78376 149671 78432
rect 149348 78374 149671 78376
rect 149348 78372 149354 78374
rect 149605 78371 149671 78374
rect 149830 78372 149836 78436
rect 149900 78434 149906 78436
rect 149973 78434 150039 78437
rect 149900 78432 150039 78434
rect 149900 78376 149978 78432
rect 150034 78376 150039 78432
rect 149900 78374 150039 78376
rect 149900 78372 149906 78374
rect 149973 78371 150039 78374
rect 152406 78372 152412 78436
rect 152476 78434 152482 78436
rect 152733 78434 152799 78437
rect 152476 78432 152799 78434
rect 152476 78376 152738 78432
rect 152794 78376 152799 78432
rect 152476 78374 152799 78376
rect 152476 78372 152482 78374
rect 152733 78371 152799 78374
rect 153193 78434 153259 78437
rect 157425 78434 157491 78437
rect 153193 78432 157491 78434
rect 153193 78376 153198 78432
rect 153254 78376 157430 78432
rect 157486 78376 157491 78432
rect 153193 78374 157491 78376
rect 153193 78371 153259 78374
rect 157425 78371 157491 78374
rect 157558 78372 157564 78436
rect 157628 78434 157634 78436
rect 157701 78434 157767 78437
rect 157628 78432 157767 78434
rect 157628 78376 157706 78432
rect 157762 78376 157767 78432
rect 157628 78374 157767 78376
rect 157628 78372 157634 78374
rect 157701 78371 157767 78374
rect 157926 78372 157932 78436
rect 157996 78434 158002 78436
rect 158161 78434 158227 78437
rect 157996 78432 158227 78434
rect 157996 78376 158166 78432
rect 158222 78376 158227 78432
rect 157996 78374 158227 78376
rect 157996 78372 158002 78374
rect 158161 78371 158227 78374
rect 165102 78372 165108 78436
rect 165172 78434 165178 78436
rect 165521 78434 165587 78437
rect 165172 78432 165587 78434
rect 165172 78376 165526 78432
rect 165582 78376 165587 78432
rect 165172 78374 165587 78376
rect 165172 78372 165178 78374
rect 165521 78371 165587 78374
rect 166390 78372 166396 78436
rect 166460 78434 166466 78436
rect 166809 78434 166875 78437
rect 166460 78432 166875 78434
rect 166460 78376 166814 78432
rect 166870 78376 166875 78432
rect 166460 78374 166875 78376
rect 166460 78372 166466 78374
rect 166809 78371 166875 78374
rect 168373 78434 168439 78437
rect 170990 78434 170996 78436
rect 168373 78432 170996 78434
rect 168373 78376 168378 78432
rect 168434 78376 170996 78432
rect 168373 78374 170996 78376
rect 168373 78371 168439 78374
rect 170990 78372 170996 78374
rect 171060 78372 171066 78436
rect 171777 78434 171843 78437
rect 174169 78434 174235 78437
rect 171777 78432 174235 78434
rect 171777 78376 171782 78432
rect 171838 78376 174174 78432
rect 174230 78376 174235 78432
rect 171777 78374 174235 78376
rect 171777 78371 171843 78374
rect 174169 78371 174235 78374
rect 130009 78298 130075 78301
rect 130326 78298 130332 78300
rect 130009 78296 130332 78298
rect 130009 78240 130014 78296
rect 130070 78240 130332 78296
rect 130009 78238 130332 78240
rect 130009 78235 130075 78238
rect 130326 78236 130332 78238
rect 130396 78236 130402 78300
rect 130929 78298 130995 78301
rect 131062 78298 131068 78300
rect 130929 78296 131068 78298
rect 130929 78240 130934 78296
rect 130990 78240 131068 78296
rect 130929 78238 131068 78240
rect 130929 78235 130995 78238
rect 131062 78236 131068 78238
rect 131132 78236 131138 78300
rect 135437 78298 135503 78301
rect 135662 78298 135668 78300
rect 135437 78296 135668 78298
rect 135437 78240 135442 78296
rect 135498 78240 135668 78296
rect 135437 78238 135668 78240
rect 135437 78235 135503 78238
rect 135662 78236 135668 78238
rect 135732 78236 135738 78300
rect 138606 78236 138612 78300
rect 138676 78298 138682 78300
rect 139025 78298 139091 78301
rect 138676 78296 139091 78298
rect 138676 78240 139030 78296
rect 139086 78240 139091 78296
rect 138676 78238 139091 78240
rect 138676 78236 138682 78238
rect 139025 78235 139091 78238
rect 140405 78300 140471 78301
rect 140405 78296 140452 78300
rect 140516 78298 140522 78300
rect 140405 78240 140410 78296
rect 140405 78236 140452 78240
rect 140516 78238 140562 78298
rect 140516 78236 140522 78238
rect 148358 78236 148364 78300
rect 148428 78298 148434 78300
rect 148869 78298 148935 78301
rect 148428 78296 148935 78298
rect 148428 78240 148874 78296
rect 148930 78240 148935 78296
rect 148428 78238 148935 78240
rect 148428 78236 148434 78238
rect 140405 78235 140471 78236
rect 148869 78235 148935 78238
rect 149462 78236 149468 78300
rect 149532 78298 149538 78300
rect 150249 78298 150315 78301
rect 149532 78296 150315 78298
rect 149532 78240 150254 78296
rect 150310 78240 150315 78296
rect 149532 78238 150315 78240
rect 149532 78236 149538 78238
rect 150249 78235 150315 78238
rect 152590 78236 152596 78300
rect 152660 78298 152666 78300
rect 153009 78298 153075 78301
rect 152660 78296 153075 78298
rect 152660 78240 153014 78296
rect 153070 78240 153075 78296
rect 152660 78238 153075 78240
rect 152660 78236 152666 78238
rect 153009 78235 153075 78238
rect 154062 78236 154068 78300
rect 154132 78298 154138 78300
rect 154389 78298 154455 78301
rect 154132 78296 154455 78298
rect 154132 78240 154394 78296
rect 154450 78240 154455 78296
rect 154132 78238 154455 78240
rect 154132 78236 154138 78238
rect 154389 78235 154455 78238
rect 157333 78298 157399 78301
rect 158294 78298 158300 78300
rect 157333 78296 158300 78298
rect 157333 78240 157338 78296
rect 157394 78240 158300 78296
rect 157333 78238 158300 78240
rect 157333 78235 157399 78238
rect 158294 78236 158300 78238
rect 158364 78236 158370 78300
rect 158805 78298 158871 78301
rect 170765 78300 170831 78301
rect 159398 78298 159404 78300
rect 158805 78296 159404 78298
rect 158805 78240 158810 78296
rect 158866 78240 159404 78296
rect 158805 78238 159404 78240
rect 158805 78235 158871 78238
rect 159398 78236 159404 78238
rect 159468 78236 159474 78300
rect 159766 78236 159772 78300
rect 159836 78298 159842 78300
rect 159836 78238 168574 78298
rect 159836 78236 159842 78238
rect 136950 78100 136956 78164
rect 137020 78162 137026 78164
rect 140497 78162 140563 78165
rect 137020 78160 140563 78162
rect 137020 78104 140502 78160
rect 140558 78104 140563 78160
rect 137020 78102 140563 78104
rect 137020 78100 137026 78102
rect 140497 78099 140563 78102
rect 140681 78162 140747 78165
rect 141366 78162 141372 78164
rect 140681 78160 141372 78162
rect 140681 78104 140686 78160
rect 140742 78104 141372 78160
rect 140681 78102 141372 78104
rect 140681 78099 140747 78102
rect 141366 78100 141372 78102
rect 141436 78100 141442 78164
rect 148542 78100 148548 78164
rect 148612 78162 148618 78164
rect 149053 78162 149119 78165
rect 148612 78160 149119 78162
rect 148612 78104 149058 78160
rect 149114 78104 149119 78160
rect 148612 78102 149119 78104
rect 148612 78100 148618 78102
rect 149053 78099 149119 78102
rect 151302 78100 151308 78164
rect 151372 78162 151378 78164
rect 151629 78162 151695 78165
rect 151372 78160 151695 78162
rect 151372 78104 151634 78160
rect 151690 78104 151695 78160
rect 151372 78102 151695 78104
rect 151372 78100 151378 78102
rect 151629 78099 151695 78102
rect 152038 78100 152044 78164
rect 152108 78162 152114 78164
rect 153193 78162 153259 78165
rect 152108 78160 153259 78162
rect 152108 78104 153198 78160
rect 153254 78104 153259 78160
rect 152108 78102 153259 78104
rect 152108 78100 152114 78102
rect 153193 78099 153259 78102
rect 153878 78100 153884 78164
rect 153948 78162 153954 78164
rect 154573 78162 154639 78165
rect 160737 78164 160803 78165
rect 153948 78160 154639 78162
rect 153948 78104 154578 78160
rect 154634 78104 154639 78160
rect 153948 78102 154639 78104
rect 153948 78100 153954 78102
rect 154573 78099 154639 78102
rect 160686 78100 160692 78164
rect 160756 78162 160803 78164
rect 160756 78160 160848 78162
rect 160798 78104 160848 78160
rect 160756 78102 160848 78104
rect 160756 78100 160803 78102
rect 161790 78100 161796 78164
rect 161860 78162 161866 78164
rect 162761 78162 162827 78165
rect 168373 78162 168439 78165
rect 161860 78160 162827 78162
rect 161860 78104 162766 78160
rect 162822 78104 162827 78160
rect 161860 78102 162827 78104
rect 161860 78100 161866 78102
rect 160737 78099 160803 78100
rect 162761 78099 162827 78102
rect 166950 78160 168439 78162
rect 166950 78104 168378 78160
rect 168434 78104 168439 78160
rect 166950 78102 168439 78104
rect 168514 78162 168574 78238
rect 170765 78296 170812 78300
rect 170876 78298 170882 78300
rect 171133 78298 171199 78301
rect 180149 78298 180215 78301
rect 170765 78240 170770 78296
rect 170765 78236 170812 78240
rect 170876 78238 170922 78298
rect 171133 78296 180215 78298
rect 171133 78240 171138 78296
rect 171194 78240 180154 78296
rect 180210 78240 180215 78296
rect 171133 78238 180215 78240
rect 170876 78236 170882 78238
rect 170765 78235 170831 78236
rect 171133 78235 171199 78238
rect 180149 78235 180215 78238
rect 171726 78162 171732 78164
rect 168514 78102 171732 78162
rect 131297 78028 131363 78029
rect 131246 78026 131252 78028
rect 131206 77966 131252 78026
rect 131316 78024 131363 78028
rect 131358 77968 131363 78024
rect 131246 77964 131252 77966
rect 131316 77964 131363 77968
rect 131297 77963 131363 77964
rect 132677 78026 132743 78029
rect 133086 78026 133092 78028
rect 132677 78024 133092 78026
rect 132677 77968 132682 78024
rect 132738 77968 133092 78024
rect 132677 77966 133092 77968
rect 132677 77963 132743 77966
rect 133086 77964 133092 77966
rect 133156 77964 133162 78028
rect 134006 77964 134012 78028
rect 134076 78026 134082 78028
rect 134149 78026 134215 78029
rect 134076 78024 134215 78026
rect 134076 77968 134154 78024
rect 134210 77968 134215 78024
rect 134076 77966 134215 77968
rect 134076 77964 134082 77966
rect 134149 77963 134215 77966
rect 140589 78028 140655 78029
rect 140589 78024 140636 78028
rect 140700 78026 140706 78028
rect 140589 77968 140594 78024
rect 140589 77964 140636 77968
rect 140700 77966 140746 78026
rect 140700 77964 140706 77966
rect 142286 77964 142292 78028
rect 142356 78026 142362 78028
rect 142429 78026 142495 78029
rect 142356 78024 142495 78026
rect 142356 77968 142434 78024
rect 142490 77968 142495 78024
rect 142356 77966 142495 77968
rect 142356 77964 142362 77966
rect 140589 77963 140655 77964
rect 142429 77963 142495 77966
rect 148777 78026 148843 78029
rect 148910 78026 148916 78028
rect 148777 78024 148916 78026
rect 148777 77968 148782 78024
rect 148838 77968 148916 78024
rect 148777 77966 148916 77968
rect 148777 77963 148843 77966
rect 148910 77964 148916 77966
rect 148980 77964 148986 78028
rect 153326 77964 153332 78028
rect 153396 78026 153402 78028
rect 154113 78026 154179 78029
rect 156137 78028 156203 78029
rect 153396 78024 154179 78026
rect 153396 77968 154118 78024
rect 154174 77968 154179 78024
rect 153396 77966 154179 77968
rect 153396 77964 153402 77966
rect 154113 77963 154179 77966
rect 156086 77964 156092 78028
rect 156156 78026 156203 78028
rect 156156 78024 156248 78026
rect 156198 77968 156248 78024
rect 156156 77966 156248 77968
rect 156156 77964 156203 77966
rect 157742 77964 157748 78028
rect 157812 78026 157818 78028
rect 158437 78026 158503 78029
rect 157812 78024 158503 78026
rect 157812 77968 158442 78024
rect 158498 77968 158503 78024
rect 157812 77966 158503 77968
rect 157812 77964 157818 77966
rect 156137 77963 156203 77964
rect 158437 77963 158503 77966
rect 159725 78026 159791 78029
rect 166950 78026 167010 78102
rect 168373 78099 168439 78102
rect 171726 78100 171732 78102
rect 171796 78100 171802 78164
rect 171910 78100 171916 78164
rect 171980 78162 171986 78164
rect 176193 78162 176259 78165
rect 171980 78160 176259 78162
rect 171980 78104 176198 78160
rect 176254 78104 176259 78160
rect 171980 78102 176259 78104
rect 171980 78100 171986 78102
rect 176193 78099 176259 78102
rect 168005 78028 168071 78029
rect 168005 78026 168052 78028
rect 159725 78024 167010 78026
rect 159725 77968 159730 78024
rect 159786 77968 167010 78024
rect 159725 77966 167010 77968
rect 167960 78024 168052 78026
rect 167960 77968 168010 78024
rect 167960 77966 168052 77968
rect 159725 77963 159791 77966
rect 168005 77964 168052 77966
rect 168116 77964 168122 78028
rect 169334 77964 169340 78028
rect 169404 78026 169410 78028
rect 170765 78026 170831 78029
rect 169404 78024 170831 78026
rect 169404 77968 170770 78024
rect 170826 77968 170831 78024
rect 169404 77966 170831 77968
rect 169404 77964 169410 77966
rect 168005 77963 168071 77964
rect 170765 77963 170831 77966
rect 175457 78026 175523 78029
rect 462313 78026 462379 78029
rect 175457 78024 462379 78026
rect 175457 77968 175462 78024
rect 175518 77968 462318 78024
rect 462374 77968 462379 78024
rect 175457 77966 462379 77968
rect 175457 77963 175523 77966
rect 462313 77963 462379 77966
rect 133137 77890 133203 77893
rect 133270 77890 133276 77892
rect 133137 77888 133276 77890
rect 133137 77832 133142 77888
rect 133198 77832 133276 77888
rect 133137 77830 133276 77832
rect 133137 77827 133203 77830
rect 133270 77828 133276 77830
rect 133340 77828 133346 77892
rect 134057 77890 134123 77893
rect 139945 77892 140011 77893
rect 134190 77890 134196 77892
rect 134057 77888 134196 77890
rect 134057 77832 134062 77888
rect 134118 77832 134196 77888
rect 134057 77830 134196 77832
rect 134057 77827 134123 77830
rect 134190 77828 134196 77830
rect 134260 77828 134266 77892
rect 139894 77828 139900 77892
rect 139964 77890 140011 77892
rect 154021 77892 154087 77893
rect 139964 77888 140056 77890
rect 140006 77832 140056 77888
rect 139964 77830 140056 77832
rect 154021 77888 154068 77892
rect 154132 77890 154138 77892
rect 162393 77890 162459 77893
rect 162526 77890 162532 77892
rect 154021 77832 154026 77888
rect 139964 77828 140011 77830
rect 139945 77827 140011 77828
rect 154021 77828 154068 77832
rect 154132 77830 154178 77890
rect 162393 77888 162532 77890
rect 162393 77832 162398 77888
rect 162454 77832 162532 77888
rect 162393 77830 162532 77832
rect 154132 77828 154138 77830
rect 154021 77827 154087 77828
rect 162393 77827 162459 77830
rect 162526 77828 162532 77830
rect 162596 77828 162602 77892
rect 164918 77828 164924 77892
rect 164988 77890 164994 77892
rect 165245 77890 165311 77893
rect 165521 77892 165587 77893
rect 165470 77890 165476 77892
rect 164988 77888 165311 77890
rect 164988 77832 165250 77888
rect 165306 77832 165311 77888
rect 164988 77830 165311 77832
rect 165430 77830 165476 77890
rect 165540 77888 165587 77892
rect 171869 77890 171935 77893
rect 165582 77832 165587 77888
rect 164988 77828 164994 77830
rect 165245 77827 165311 77830
rect 165470 77828 165476 77830
rect 165540 77828 165587 77832
rect 165521 77827 165587 77828
rect 166950 77888 171935 77890
rect 166950 77832 171874 77888
rect 171930 77832 171935 77888
rect 166950 77830 171935 77832
rect 129181 77754 129247 77757
rect 130694 77754 130700 77756
rect 129181 77752 130700 77754
rect 129181 77696 129186 77752
rect 129242 77696 130700 77752
rect 129181 77694 130700 77696
rect 129181 77691 129247 77694
rect 130694 77692 130700 77694
rect 130764 77692 130770 77756
rect 156454 77692 156460 77756
rect 156524 77754 156530 77756
rect 166950 77754 167010 77830
rect 171869 77827 171935 77830
rect 156524 77694 167010 77754
rect 167177 77754 167243 77757
rect 172094 77754 172100 77756
rect 167177 77752 172100 77754
rect 167177 77696 167182 77752
rect 167238 77696 172100 77752
rect 167177 77694 172100 77696
rect 156524 77692 156530 77694
rect 167177 77691 167243 77694
rect 172094 77692 172100 77694
rect 172164 77692 172170 77756
rect 145230 77556 145236 77620
rect 145300 77618 145306 77620
rect 146017 77618 146083 77621
rect 145300 77616 146083 77618
rect 145300 77560 146022 77616
rect 146078 77560 146083 77616
rect 145300 77558 146083 77560
rect 145300 77556 145306 77558
rect 146017 77555 146083 77558
rect 157057 77618 157123 77621
rect 157057 77616 167194 77618
rect 157057 77560 157062 77616
rect 157118 77560 167194 77616
rect 157057 77558 167194 77560
rect 157057 77555 157123 77558
rect 160686 77420 160692 77484
rect 160756 77482 160762 77484
rect 161197 77482 161263 77485
rect 160756 77480 161263 77482
rect 160756 77424 161202 77480
rect 161258 77424 161263 77480
rect 160756 77422 161263 77424
rect 160756 77420 160762 77422
rect 161197 77419 161263 77422
rect 162342 77420 162348 77484
rect 162412 77482 162418 77484
rect 162577 77482 162643 77485
rect 162412 77480 162643 77482
rect 162412 77424 162582 77480
rect 162638 77424 162643 77480
rect 162412 77422 162643 77424
rect 162412 77420 162418 77422
rect 162577 77419 162643 77422
rect 165337 77482 165403 77485
rect 165470 77482 165476 77484
rect 165337 77480 165476 77482
rect 165337 77424 165342 77480
rect 165398 77424 165476 77480
rect 165337 77422 165476 77424
rect 165337 77419 165403 77422
rect 165470 77420 165476 77422
rect 165540 77420 165546 77484
rect 166206 77420 166212 77484
rect 166276 77482 166282 77484
rect 166809 77482 166875 77485
rect 166276 77480 166875 77482
rect 166276 77424 166814 77480
rect 166870 77424 166875 77480
rect 166276 77422 166875 77424
rect 167134 77482 167194 77558
rect 167862 77556 167868 77620
rect 167932 77618 167938 77620
rect 168097 77618 168163 77621
rect 172237 77618 172303 77621
rect 167932 77616 168163 77618
rect 167932 77560 168102 77616
rect 168158 77560 168163 77616
rect 167932 77558 168163 77560
rect 167932 77556 167938 77558
rect 168097 77555 168163 77558
rect 168238 77616 172303 77618
rect 168238 77560 172242 77616
rect 172298 77560 172303 77616
rect 168238 77558 172303 77560
rect 168238 77482 168298 77558
rect 172237 77555 172303 77558
rect 167134 77422 168298 77482
rect 168649 77482 168715 77485
rect 171910 77482 171916 77484
rect 168649 77480 171916 77482
rect 168649 77424 168654 77480
rect 168710 77424 171916 77480
rect 168649 77422 171916 77424
rect 166276 77420 166282 77422
rect 166809 77419 166875 77422
rect 168649 77419 168715 77422
rect 171910 77420 171916 77422
rect 171980 77420 171986 77484
rect 125542 77284 125548 77348
rect 125612 77346 125618 77348
rect 126094 77346 126100 77348
rect 125612 77286 126100 77346
rect 125612 77284 125618 77286
rect 126094 77284 126100 77286
rect 126164 77284 126170 77348
rect 166206 77284 166212 77348
rect 166276 77346 166282 77348
rect 166717 77346 166783 77349
rect 166276 77344 166783 77346
rect 166276 77288 166722 77344
rect 166778 77288 166783 77344
rect 166276 77286 166783 77288
rect 166276 77284 166282 77286
rect 166717 77283 166783 77286
rect 167310 77284 167316 77348
rect 167380 77346 167386 77348
rect 167545 77346 167611 77349
rect 167380 77344 167611 77346
rect 167380 77288 167550 77344
rect 167606 77288 167611 77344
rect 167380 77286 167611 77288
rect 167380 77284 167386 77286
rect 167545 77283 167611 77286
rect 168046 77284 168052 77348
rect 168116 77346 168122 77348
rect 168189 77346 168255 77349
rect 168116 77344 168255 77346
rect 168116 77288 168194 77344
rect 168250 77288 168255 77344
rect 168116 77286 168255 77288
rect 168116 77284 168122 77286
rect 168189 77283 168255 77286
rect 170070 77284 170076 77348
rect 170140 77346 170146 77348
rect 170213 77346 170279 77349
rect 170140 77344 170279 77346
rect 170140 77288 170218 77344
rect 170274 77288 170279 77344
rect 170140 77286 170279 77288
rect 170140 77284 170146 77286
rect 170213 77283 170279 77286
rect 171174 77284 171180 77348
rect 171244 77346 171250 77348
rect 172278 77346 172284 77348
rect 171244 77286 172284 77346
rect 171244 77284 171250 77286
rect 172278 77284 172284 77286
rect 172348 77284 172354 77348
rect 178769 77346 178835 77349
rect 182817 77346 182883 77349
rect 178769 77344 182883 77346
rect 178769 77288 178774 77344
rect 178830 77288 182822 77344
rect 182878 77288 182883 77344
rect 178769 77286 182883 77288
rect 178769 77283 178835 77286
rect 182817 77283 182883 77286
rect 71773 77210 71839 77213
rect 172881 77210 172947 77213
rect 71773 77208 172947 77210
rect 71773 77152 71778 77208
rect 71834 77152 172886 77208
rect 172942 77152 172947 77208
rect 71773 77150 172947 77152
rect 71773 77147 71839 77150
rect 172881 77147 172947 77150
rect 129641 77074 129707 77077
rect 130142 77074 130148 77076
rect 129641 77072 130148 77074
rect 129641 77016 129646 77072
rect 129702 77016 130148 77072
rect 129641 77014 130148 77016
rect 129641 77011 129707 77014
rect 130142 77012 130148 77014
rect 130212 77012 130218 77076
rect 158345 77074 158411 77077
rect 158478 77074 158484 77076
rect 158345 77072 158484 77074
rect 158345 77016 158350 77072
rect 158406 77016 158484 77072
rect 158345 77014 158484 77016
rect 158345 77011 158411 77014
rect 158478 77012 158484 77014
rect 158548 77012 158554 77076
rect 161422 77012 161428 77076
rect 161492 77074 161498 77076
rect 173157 77074 173223 77077
rect 161492 77072 173223 77074
rect 161492 77016 173162 77072
rect 173218 77016 173223 77072
rect 161492 77014 173223 77016
rect 161492 77012 161498 77014
rect 173157 77011 173223 77014
rect 142102 76876 142108 76940
rect 142172 76938 142178 76940
rect 173341 76938 173407 76941
rect 142172 76936 173407 76938
rect 142172 76880 173346 76936
rect 173402 76880 173407 76936
rect 142172 76878 173407 76880
rect 142172 76876 142178 76878
rect 173341 76875 173407 76878
rect 111793 76802 111859 76805
rect 133873 76802 133939 76805
rect 111793 76800 133939 76802
rect 111793 76744 111798 76800
rect 111854 76744 133878 76800
rect 133934 76744 133939 76800
rect 111793 76742 133939 76744
rect 111793 76739 111859 76742
rect 133873 76739 133939 76742
rect 146385 76802 146451 76805
rect 247033 76802 247099 76805
rect 146385 76800 247099 76802
rect 146385 76744 146390 76800
rect 146446 76744 247038 76800
rect 247094 76744 247099 76800
rect 146385 76742 247099 76744
rect 146385 76739 146451 76742
rect 247033 76739 247099 76742
rect 37273 76666 37339 76669
rect 128445 76666 128511 76669
rect 37273 76664 128511 76666
rect 37273 76608 37278 76664
rect 37334 76608 128450 76664
rect 128506 76608 128511 76664
rect 37273 76606 128511 76608
rect 37273 76603 37339 76606
rect 128445 76603 128511 76606
rect 147673 76666 147739 76669
rect 282913 76666 282979 76669
rect 147673 76664 282979 76666
rect 147673 76608 147678 76664
rect 147734 76608 282918 76664
rect 282974 76608 282979 76664
rect 147673 76606 282979 76608
rect 147673 76603 147739 76606
rect 282913 76603 282979 76606
rect 20713 76530 20779 76533
rect 127249 76530 127315 76533
rect 166073 76532 166139 76533
rect 20713 76528 127315 76530
rect 20713 76472 20718 76528
rect 20774 76472 127254 76528
rect 127310 76472 127315 76528
rect 20713 76470 127315 76472
rect 20713 76467 20779 76470
rect 127249 76467 127315 76470
rect 166022 76468 166028 76532
rect 166092 76530 166139 76532
rect 166092 76528 166184 76530
rect 166134 76472 166184 76528
rect 166092 76470 166184 76472
rect 166092 76468 166139 76470
rect 169702 76468 169708 76532
rect 169772 76530 169778 76532
rect 565813 76530 565879 76533
rect 169772 76528 565879 76530
rect 169772 76472 565818 76528
rect 565874 76472 565879 76528
rect 169772 76470 565879 76472
rect 169772 76468 169778 76470
rect 166073 76467 166139 76468
rect 565813 76467 565879 76470
rect 170489 76394 170555 76397
rect 170990 76394 170996 76396
rect 170489 76392 170996 76394
rect 170489 76336 170494 76392
rect 170550 76336 170996 76392
rect 170489 76334 170996 76336
rect 170489 76331 170555 76334
rect 170990 76332 170996 76334
rect 171060 76332 171066 76396
rect 170622 76196 170628 76260
rect 170692 76258 170698 76260
rect 171041 76258 171107 76261
rect 170692 76256 171107 76258
rect 170692 76200 171046 76256
rect 171102 76200 171107 76256
rect 170692 76198 171107 76200
rect 170692 76196 170698 76198
rect 171041 76195 171107 76198
rect 163446 75924 163452 75988
rect 163516 75986 163522 75988
rect 164417 75986 164483 75989
rect 163516 75984 164483 75986
rect 163516 75928 164422 75984
rect 164478 75928 164483 75984
rect 163516 75926 164483 75928
rect 163516 75924 163522 75926
rect 164417 75923 164483 75926
rect 138606 75788 138612 75852
rect 138676 75850 138682 75852
rect 173893 75850 173959 75853
rect 138676 75848 173959 75850
rect 138676 75792 173898 75848
rect 173954 75792 173959 75848
rect 138676 75790 173959 75792
rect 138676 75788 138682 75790
rect 173893 75787 173959 75790
rect 151670 75652 151676 75716
rect 151740 75714 151746 75716
rect 193857 75714 193923 75717
rect 151740 75712 193923 75714
rect 151740 75656 193862 75712
rect 193918 75656 193923 75712
rect 151740 75654 193923 75656
rect 151740 75652 151746 75654
rect 193857 75651 193923 75654
rect 89713 75578 89779 75581
rect 133454 75578 133460 75580
rect 89713 75576 133460 75578
rect 89713 75520 89718 75576
rect 89774 75520 133460 75576
rect 89713 75518 133460 75520
rect 89713 75515 89779 75518
rect 133454 75516 133460 75518
rect 133524 75516 133530 75580
rect 151302 75516 151308 75580
rect 151372 75578 151378 75580
rect 154665 75578 154731 75581
rect 151372 75576 154731 75578
rect 151372 75520 154670 75576
rect 154726 75520 154731 75576
rect 151372 75518 154731 75520
rect 151372 75516 151378 75518
rect 154665 75515 154731 75518
rect 157190 75516 157196 75580
rect 157260 75578 157266 75580
rect 339125 75578 339191 75581
rect 157260 75576 339191 75578
rect 157260 75520 339130 75576
rect 339186 75520 339191 75576
rect 157260 75518 339191 75520
rect 157260 75516 157266 75518
rect 339125 75515 339191 75518
rect 75913 75442 75979 75445
rect 131430 75442 131436 75444
rect 75913 75440 131436 75442
rect 75913 75384 75918 75440
rect 75974 75384 131436 75440
rect 75913 75382 131436 75384
rect 75913 75379 75979 75382
rect 131430 75380 131436 75382
rect 131500 75380 131506 75444
rect 155718 75380 155724 75444
rect 155788 75442 155794 75444
rect 369117 75442 369183 75445
rect 155788 75440 369183 75442
rect 155788 75384 369122 75440
rect 369178 75384 369183 75440
rect 155788 75382 369183 75384
rect 155788 75380 155794 75382
rect 369117 75379 369183 75382
rect 2773 75306 2839 75309
rect 125542 75306 125548 75308
rect 2773 75304 125548 75306
rect 2773 75248 2778 75304
rect 2834 75248 125548 75304
rect 2773 75246 125548 75248
rect 2773 75243 2839 75246
rect 125542 75244 125548 75246
rect 125612 75244 125618 75308
rect 133965 75306 134031 75309
rect 134374 75306 134380 75308
rect 133965 75304 134380 75306
rect 133965 75248 133970 75304
rect 134026 75248 134380 75304
rect 133965 75246 134380 75248
rect 133965 75243 134031 75246
rect 134374 75244 134380 75246
rect 134444 75244 134450 75308
rect 135437 75306 135503 75309
rect 135662 75306 135668 75308
rect 135437 75304 135668 75306
rect 135437 75248 135442 75304
rect 135498 75248 135668 75304
rect 135437 75246 135668 75248
rect 135437 75243 135503 75246
rect 135662 75244 135668 75246
rect 135732 75244 135738 75308
rect 158294 75244 158300 75308
rect 158364 75306 158370 75308
rect 158437 75306 158503 75309
rect 161105 75308 161171 75309
rect 158364 75304 158503 75306
rect 158364 75248 158442 75304
rect 158498 75248 158503 75304
rect 158364 75246 158503 75248
rect 158364 75244 158370 75246
rect 158437 75243 158503 75246
rect 161054 75244 161060 75308
rect 161124 75306 161171 75308
rect 161749 75306 161815 75309
rect 161974 75306 161980 75308
rect 161124 75304 161216 75306
rect 161166 75248 161216 75304
rect 161124 75246 161216 75248
rect 161749 75304 161980 75306
rect 161749 75248 161754 75304
rect 161810 75248 161980 75304
rect 161749 75246 161980 75248
rect 161124 75244 161171 75246
rect 161105 75243 161171 75244
rect 161749 75243 161815 75246
rect 161974 75244 161980 75246
rect 162044 75244 162050 75308
rect 162342 75244 162348 75308
rect 162412 75306 162418 75308
rect 162577 75306 162643 75309
rect 162412 75304 162643 75306
rect 162412 75248 162582 75304
rect 162638 75248 162643 75304
rect 162412 75246 162643 75248
rect 162412 75244 162418 75246
rect 162577 75243 162643 75246
rect 163630 75244 163636 75308
rect 163700 75306 163706 75308
rect 163957 75306 164023 75309
rect 163700 75304 164023 75306
rect 163700 75248 163962 75304
rect 164018 75248 164023 75304
rect 163700 75246 164023 75248
rect 163700 75244 163706 75246
rect 163957 75243 164023 75246
rect 164141 75306 164207 75309
rect 496813 75306 496879 75309
rect 164141 75304 496879 75306
rect 164141 75248 164146 75304
rect 164202 75248 496818 75304
rect 496874 75248 496879 75304
rect 164141 75246 496879 75248
rect 164141 75243 164207 75246
rect 496813 75243 496879 75246
rect 1393 75170 1459 75173
rect 125726 75170 125732 75172
rect 1393 75168 125732 75170
rect 1393 75112 1398 75168
rect 1454 75112 125732 75168
rect 1393 75110 125732 75112
rect 1393 75107 1459 75110
rect 125726 75108 125732 75110
rect 125796 75108 125802 75172
rect 130377 75170 130443 75173
rect 135294 75170 135300 75172
rect 130377 75168 135300 75170
rect 130377 75112 130382 75168
rect 130438 75112 135300 75168
rect 130377 75110 135300 75112
rect 130377 75107 130443 75110
rect 135294 75108 135300 75110
rect 135364 75108 135370 75172
rect 160001 75170 160067 75173
rect 160134 75170 160140 75172
rect 160001 75168 160140 75170
rect 160001 75112 160006 75168
rect 160062 75112 160140 75168
rect 160001 75110 160140 75112
rect 160001 75107 160067 75110
rect 160134 75108 160140 75110
rect 160204 75108 160210 75172
rect 170438 75108 170444 75172
rect 170508 75170 170514 75172
rect 171961 75170 172027 75173
rect 549253 75170 549319 75173
rect 170508 75168 172027 75170
rect 170508 75112 171966 75168
rect 172022 75112 172027 75168
rect 170508 75110 172027 75112
rect 170508 75108 170514 75110
rect 171961 75107 172027 75110
rect 176610 75168 549319 75170
rect 176610 75112 549258 75168
rect 549314 75112 549319 75168
rect 176610 75110 549319 75112
rect 169150 74972 169156 75036
rect 169220 75034 169226 75036
rect 176610 75034 176670 75110
rect 549253 75107 549319 75110
rect 169220 74974 176670 75034
rect 169220 74972 169226 74974
rect 140078 74428 140084 74492
rect 140148 74490 140154 74492
rect 194593 74490 194659 74493
rect 140148 74488 194659 74490
rect 140148 74432 194598 74488
rect 194654 74432 194659 74488
rect 140148 74430 194659 74432
rect 140148 74428 140154 74430
rect 194593 74427 194659 74430
rect 142838 74292 142844 74356
rect 142908 74354 142914 74356
rect 230473 74354 230539 74357
rect 142908 74352 230539 74354
rect 142908 74296 230478 74352
rect 230534 74296 230539 74352
rect 142908 74294 230539 74296
rect 142908 74292 142914 74294
rect 230473 74291 230539 74294
rect 144678 74156 144684 74220
rect 144748 74218 144754 74220
rect 244273 74218 244339 74221
rect 144748 74216 244339 74218
rect 144748 74160 244278 74216
rect 244334 74160 244339 74216
rect 144748 74158 244339 74160
rect 144748 74156 144754 74158
rect 244273 74155 244339 74158
rect 71773 74082 71839 74085
rect 131614 74082 131620 74084
rect 71773 74080 131620 74082
rect 71773 74024 71778 74080
rect 71834 74024 131620 74080
rect 71773 74022 131620 74024
rect 71773 74019 71839 74022
rect 131614 74020 131620 74022
rect 131684 74020 131690 74084
rect 155902 74020 155908 74084
rect 155972 74082 155978 74084
rect 156873 74082 156939 74085
rect 155972 74080 156939 74082
rect 155972 74024 156878 74080
rect 156934 74024 156939 74080
rect 155972 74022 156939 74024
rect 155972 74020 155978 74022
rect 156873 74019 156939 74022
rect 157006 74020 157012 74084
rect 157076 74082 157082 74084
rect 349797 74082 349863 74085
rect 157076 74080 349863 74082
rect 157076 74024 349802 74080
rect 349858 74024 349863 74080
rect 157076 74022 349863 74024
rect 157076 74020 157082 74022
rect 349797 74019 349863 74022
rect 57973 73946 58039 73949
rect 130142 73946 130148 73948
rect 57973 73944 130148 73946
rect 57973 73888 57978 73944
rect 58034 73888 130148 73944
rect 57973 73886 130148 73888
rect 57973 73883 58039 73886
rect 130142 73884 130148 73886
rect 130212 73884 130218 73948
rect 156822 73884 156828 73948
rect 156892 73946 156898 73948
rect 378409 73946 378475 73949
rect 156892 73944 378475 73946
rect 156892 73888 378414 73944
rect 378470 73888 378475 73944
rect 156892 73886 378475 73888
rect 156892 73884 156898 73886
rect 378409 73883 378475 73886
rect 53833 73810 53899 73813
rect 129774 73810 129780 73812
rect 53833 73808 129780 73810
rect 53833 73752 53838 73808
rect 53894 73752 129780 73808
rect 53833 73750 129780 73752
rect 53833 73747 53899 73750
rect 129774 73748 129780 73750
rect 129844 73748 129850 73812
rect 170305 73810 170371 73813
rect 578233 73810 578299 73813
rect 170305 73808 578299 73810
rect 170305 73752 170310 73808
rect 170366 73752 578238 73808
rect 578294 73752 578299 73808
rect 170305 73750 578299 73752
rect 170305 73747 170371 73750
rect 578233 73747 578299 73750
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect 156638 72524 156644 72588
rect 156708 72586 156714 72588
rect 296069 72586 296135 72589
rect 156708 72584 296135 72586
rect 156708 72528 296074 72584
rect 296130 72528 296135 72584
rect 156708 72526 296135 72528
rect 156708 72524 156714 72526
rect 296069 72523 296135 72526
rect 148910 72388 148916 72452
rect 148980 72450 148986 72452
rect 298093 72450 298159 72453
rect 148980 72448 298159 72450
rect 148980 72392 298098 72448
rect 298154 72392 298159 72448
rect 148980 72390 298159 72392
rect 148980 72388 148986 72390
rect 298093 72387 298159 72390
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 151486 71028 151492 71092
rect 151556 71090 151562 71092
rect 306925 71090 306991 71093
rect 151556 71088 306991 71090
rect 151556 71032 306930 71088
rect 306986 71032 306991 71088
rect 151556 71030 306991 71032
rect 151556 71028 151562 71030
rect 306925 71027 306991 71030
rect 138790 68444 138796 68508
rect 138860 68506 138866 68508
rect 175273 68506 175339 68509
rect 138860 68504 175339 68506
rect 138860 68448 175278 68504
rect 175334 68448 175339 68504
rect 138860 68446 175339 68448
rect 138860 68444 138866 68446
rect 175273 68443 175339 68446
rect 140262 68308 140268 68372
rect 140332 68370 140338 68372
rect 193213 68370 193279 68373
rect 140332 68368 193279 68370
rect 140332 68312 193218 68368
rect 193274 68312 193279 68368
rect 140332 68310 193279 68312
rect 140332 68308 140338 68310
rect 193213 68307 193279 68310
rect 152958 68172 152964 68236
rect 153028 68234 153034 68236
rect 353293 68234 353359 68237
rect 153028 68232 353359 68234
rect 153028 68176 353298 68232
rect 353354 68176 353359 68232
rect 153028 68174 353359 68176
rect 153028 68172 153034 68174
rect 353293 68171 353359 68174
rect 166206 66948 166212 67012
rect 166276 67010 166282 67012
rect 529933 67010 529999 67013
rect 166276 67008 529999 67010
rect 166276 66952 529938 67008
rect 529994 66952 529999 67008
rect 166276 66950 529999 66952
rect 166276 66948 166282 66950
rect 529933 66947 529999 66950
rect 167678 66812 167684 66876
rect 167748 66874 167754 66876
rect 547873 66874 547939 66877
rect 167748 66872 547939 66874
rect 167748 66816 547878 66872
rect 547934 66816 547939 66872
rect 167748 66814 547939 66816
rect 167748 66812 167754 66814
rect 547873 66811 547939 66814
rect 163446 65452 163452 65516
rect 163516 65514 163522 65516
rect 494053 65514 494119 65517
rect 163516 65512 494119 65514
rect 163516 65456 494058 65512
rect 494114 65456 494119 65512
rect 163516 65454 494119 65456
rect 163516 65452 163522 65454
rect 494053 65451 494119 65454
rect 164918 64092 164924 64156
rect 164988 64154 164994 64156
rect 511993 64154 512059 64157
rect 164988 64152 512059 64154
rect 164988 64096 511998 64152
rect 512054 64096 512059 64152
rect 164988 64094 512059 64096
rect 164988 64092 164994 64094
rect 511993 64091 512059 64094
rect 145230 62732 145236 62796
rect 145300 62794 145306 62796
rect 263593 62794 263659 62797
rect 145300 62792 263659 62794
rect 145300 62736 263598 62792
rect 263654 62736 263659 62792
rect 145300 62734 263659 62736
rect 145300 62732 145306 62734
rect 263593 62731 263659 62734
rect 172278 61372 172284 61436
rect 172348 61434 172354 61436
rect 431953 61434 432019 61437
rect 172348 61432 432019 61434
rect 172348 61376 431958 61432
rect 432014 61376 432019 61432
rect 172348 61374 432019 61376
rect 172348 61372 172354 61374
rect 431953 61371 432019 61374
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 144494 58516 144500 58580
rect 144564 58578 144570 58580
rect 245653 58578 245719 58581
rect 144564 58576 245719 58578
rect 144564 58520 245658 58576
rect 245714 58520 245719 58576
rect 144564 58518 245719 58520
rect 144564 58516 144570 58518
rect 245653 58515 245719 58518
rect 152590 51716 152596 51780
rect 152660 51778 152666 51780
rect 351913 51778 351979 51781
rect 152660 51776 351979 51778
rect 152660 51720 351918 51776
rect 351974 51720 351979 51776
rect 152660 51718 351979 51720
rect 152660 51716 152666 51718
rect 351913 51715 351979 51718
rect 172094 48860 172100 48924
rect 172164 48922 172170 48924
rect 425053 48922 425119 48925
rect 172164 48920 425119 48922
rect 172164 48864 425058 48920
rect 425114 48864 425119 48920
rect 172164 48862 425119 48864
rect 172164 48860 172170 48862
rect 425053 48859 425119 48862
rect 171910 47500 171916 47564
rect 171980 47562 171986 47564
rect 550633 47562 550699 47565
rect 171980 47560 550699 47562
rect 171980 47504 550638 47560
rect 550694 47504 550699 47560
rect 171980 47502 550699 47504
rect 171980 47500 171986 47502
rect 550633 47499 550699 47502
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 91093 44842 91159 44845
rect 133270 44842 133276 44844
rect 91093 44840 133276 44842
rect 91093 44784 91098 44840
rect 91154 44784 133276 44840
rect 91093 44782 133276 44784
rect 91093 44779 91159 44782
rect 133270 44780 133276 44782
rect 133340 44780 133346 44844
rect 171726 42060 171732 42124
rect 171796 42122 171802 42124
rect 440233 42122 440299 42125
rect 171796 42120 440299 42122
rect 171796 42064 440238 42120
rect 440294 42064 440299 42120
rect 171796 42062 440299 42064
rect 171796 42060 171802 42062
rect 440233 42059 440299 42062
rect 153878 35124 153884 35188
rect 153948 35186 153954 35188
rect 372613 35186 372679 35189
rect 153948 35184 372679 35186
rect 153948 35128 372618 35184
rect 372674 35128 372679 35184
rect 153948 35126 372679 35128
rect 153948 35124 153954 35126
rect 372613 35123 372679 35126
rect 140446 34036 140452 34100
rect 140516 34098 140522 34100
rect 191833 34098 191899 34101
rect 140516 34096 191899 34098
rect 140516 34040 191838 34096
rect 191894 34040 191899 34096
rect 140516 34038 191899 34040
rect 140516 34036 140522 34038
rect 191833 34035 191899 34038
rect 143022 33900 143028 33964
rect 143092 33962 143098 33964
rect 226425 33962 226491 33965
rect 143092 33960 226491 33962
rect 143092 33904 226430 33960
rect 226486 33904 226491 33960
rect 143092 33902 226491 33904
rect 143092 33900 143098 33902
rect 226425 33899 226491 33902
rect 145414 33764 145420 33828
rect 145484 33826 145490 33828
rect 266353 33826 266419 33829
rect 145484 33824 266419 33826
rect 145484 33768 266358 33824
rect 266414 33768 266419 33824
rect 145484 33766 266419 33768
rect 145484 33764 145490 33766
rect 266353 33763 266419 33766
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 138974 32540 138980 32604
rect 139044 32602 139050 32604
rect 176653 32602 176719 32605
rect 139044 32600 176719 32602
rect 139044 32544 176658 32600
rect 176714 32544 176719 32600
rect 139044 32542 176719 32544
rect 139044 32540 139050 32542
rect 176653 32539 176719 32542
rect 3417 32466 3483 32469
rect -960 32464 3483 32466
rect -960 32408 3422 32464
rect 3478 32408 3483 32464
rect -960 32406 3483 32408
rect -960 32316 480 32406
rect 3417 32403 3483 32406
rect 165102 32404 165108 32468
rect 165172 32466 165178 32468
rect 514845 32466 514911 32469
rect 165172 32464 514911 32466
rect 165172 32408 514850 32464
rect 514906 32408 514911 32464
rect 165172 32406 514911 32408
rect 165172 32404 165178 32406
rect 514845 32403 514911 32406
rect 149462 29820 149468 29884
rect 149532 29882 149538 29884
rect 317413 29882 317479 29885
rect 149532 29880 317479 29882
rect 149532 29824 317418 29880
rect 317474 29824 317479 29880
rect 149532 29822 317479 29824
rect 149532 29820 149538 29822
rect 317413 29819 317479 29822
rect 152774 29684 152780 29748
rect 152844 29746 152850 29748
rect 349153 29746 349219 29749
rect 152844 29744 349219 29746
rect 152844 29688 349158 29744
rect 349214 29688 349219 29744
rect 152844 29686 349219 29688
rect 152844 29684 152850 29686
rect 349153 29683 349219 29686
rect 169518 29548 169524 29612
rect 169588 29610 169594 29612
rect 567193 29610 567259 29613
rect 169588 29608 567259 29610
rect 169588 29552 567198 29608
rect 567254 29552 567259 29608
rect 169588 29550 567259 29552
rect 169588 29548 169594 29550
rect 567193 29547 567259 29550
rect 140630 25468 140636 25532
rect 140700 25530 140706 25532
rect 193305 25530 193371 25533
rect 140700 25528 193371 25530
rect 140700 25472 193310 25528
rect 193366 25472 193371 25528
rect 140700 25470 193371 25472
rect 140700 25468 140706 25470
rect 193305 25467 193371 25470
rect 127617 22674 127683 22677
rect 135662 22674 135668 22676
rect 127617 22672 135668 22674
rect 127617 22616 127622 22672
rect 127678 22616 135668 22672
rect 127617 22614 135668 22616
rect 127617 22611 127683 22614
rect 135662 22612 135668 22614
rect 135732 22612 135738 22676
rect 157926 22612 157932 22676
rect 157996 22674 158002 22676
rect 422293 22674 422359 22677
rect 157996 22672 422359 22674
rect 157996 22616 422298 22672
rect 422354 22616 422359 22672
rect 157996 22614 422359 22616
rect 157996 22612 158002 22614
rect 422293 22611 422359 22614
rect 166390 21252 166396 21316
rect 166460 21314 166466 21316
rect 531313 21314 531379 21317
rect 166460 21312 531379 21314
rect 166460 21256 531318 21312
rect 531374 21256 531379 21312
rect 166460 21254 531379 21256
rect 166460 21252 166466 21254
rect 531313 21251 531379 21254
rect 144126 20028 144132 20092
rect 144196 20090 144202 20092
rect 248413 20090 248479 20093
rect 144196 20088 248479 20090
rect 144196 20032 248418 20088
rect 248474 20032 248479 20088
rect 144196 20030 248479 20032
rect 144196 20028 144202 20030
rect 248413 20027 248479 20030
rect 42793 19954 42859 19957
rect 128854 19954 128860 19956
rect 42793 19952 128860 19954
rect 42793 19896 42798 19952
rect 42854 19896 128860 19952
rect 42793 19894 128860 19896
rect 42793 19891 42859 19894
rect 128854 19892 128860 19894
rect 128924 19892 128930 19956
rect 137686 19892 137692 19956
rect 137756 19954 137762 19956
rect 160093 19954 160159 19957
rect 137756 19952 160159 19954
rect 137756 19896 160098 19952
rect 160154 19896 160159 19952
rect 137756 19894 160159 19896
rect 137756 19892 137762 19894
rect 160093 19891 160159 19894
rect 165286 19892 165292 19956
rect 165356 19954 165362 19956
rect 513373 19954 513439 19957
rect 165356 19952 513439 19954
rect 165356 19896 513378 19952
rect 513434 19896 513439 19952
rect 165356 19894 513439 19896
rect 165356 19892 165362 19894
rect 513373 19891 513439 19894
rect 579613 19818 579679 19821
rect 583520 19818 584960 19908
rect 579613 19816 584960 19818
rect 579613 19760 579618 19816
rect 579674 19760 584960 19816
rect 579613 19758 584960 19760
rect 579613 19755 579679 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3325 19410 3391 19413
rect -960 19408 3391 19410
rect -960 19352 3330 19408
rect 3386 19352 3391 19408
rect -960 19350 3391 19352
rect -960 19260 480 19350
rect 3325 19347 3391 19350
rect 167862 18532 167868 18596
rect 167932 18594 167938 18596
rect 546493 18594 546559 18597
rect 167932 18592 546559 18594
rect 167932 18536 546498 18592
rect 546554 18536 546559 18592
rect 167932 18534 546559 18536
rect 167932 18532 167938 18534
rect 546493 18531 546559 18534
rect 140998 17580 141004 17644
rect 141068 17642 141074 17644
rect 212533 17642 212599 17645
rect 141068 17640 212599 17642
rect 141068 17584 212538 17640
rect 212594 17584 212599 17640
rect 141068 17582 212599 17584
rect 141068 17580 141074 17582
rect 212533 17579 212599 17582
rect 148542 17444 148548 17508
rect 148612 17506 148618 17508
rect 300853 17506 300919 17509
rect 148612 17504 300919 17506
rect 148612 17448 300858 17504
rect 300914 17448 300919 17504
rect 148612 17446 300919 17448
rect 148612 17444 148618 17446
rect 300853 17443 300919 17446
rect 158110 17308 158116 17372
rect 158180 17370 158186 17372
rect 423673 17370 423739 17373
rect 158180 17368 423739 17370
rect 158180 17312 423678 17368
rect 423734 17312 423739 17368
rect 158180 17310 423739 17312
rect 158180 17308 158186 17310
rect 423673 17307 423739 17310
rect 163630 17172 163636 17236
rect 163700 17234 163706 17236
rect 495433 17234 495499 17237
rect 163700 17232 495499 17234
rect 163700 17176 495438 17232
rect 495494 17176 495499 17232
rect 163700 17174 495499 17176
rect 163700 17172 163706 17174
rect 495433 17171 495499 17174
rect 154062 15812 154068 15876
rect 154132 15874 154138 15876
rect 365713 15874 365779 15877
rect 154132 15872 365779 15874
rect 154132 15816 365718 15872
rect 365774 15816 365779 15872
rect 154132 15814 365779 15816
rect 154132 15812 154138 15814
rect 365713 15811 365779 15814
rect 158846 14724 158852 14788
rect 158916 14786 158922 14788
rect 442625 14786 442691 14789
rect 158916 14784 442691 14786
rect 158916 14728 442630 14784
rect 442686 14728 442691 14784
rect 158916 14726 442691 14728
rect 158916 14724 158922 14726
rect 442625 14723 442691 14726
rect 159030 14588 159036 14652
rect 159100 14650 159106 14652
rect 443361 14650 443427 14653
rect 159100 14648 443427 14650
rect 159100 14592 443366 14648
rect 443422 14592 443427 14648
rect 159100 14590 443427 14592
rect 159100 14588 159106 14590
rect 443361 14587 443427 14590
rect 165470 14452 165476 14516
rect 165540 14514 165546 14516
rect 511257 14514 511323 14517
rect 165540 14512 511323 14514
rect 165540 14456 511262 14512
rect 511318 14456 511323 14512
rect 165540 14454 511323 14456
rect 165540 14452 165546 14454
rect 511257 14451 511323 14454
rect 143206 13364 143212 13428
rect 143276 13426 143282 13428
rect 229369 13426 229435 13429
rect 143276 13424 229435 13426
rect 143276 13368 229374 13424
rect 229430 13368 229435 13424
rect 143276 13366 229435 13368
rect 143276 13364 143282 13366
rect 229369 13363 229435 13366
rect 154430 13228 154436 13292
rect 154500 13290 154506 13292
rect 370129 13290 370195 13293
rect 154500 13288 370195 13290
rect 154500 13232 370134 13288
rect 370190 13232 370195 13288
rect 154500 13230 370195 13232
rect 154500 13228 154506 13230
rect 370129 13227 370195 13230
rect 154246 13092 154252 13156
rect 154316 13154 154322 13156
rect 371233 13154 371299 13157
rect 154316 13152 371299 13154
rect 154316 13096 371238 13152
rect 371294 13096 371299 13152
rect 154316 13094 371299 13096
rect 154316 13092 154322 13094
rect 371233 13091 371299 13094
rect 166574 12956 166580 13020
rect 166644 13018 166650 13020
rect 532049 13018 532115 13021
rect 166644 13016 532115 13018
rect 166644 12960 532054 13016
rect 532110 12960 532115 13016
rect 166644 12958 532115 12960
rect 166644 12956 166650 12958
rect 532049 12955 532115 12958
rect 158294 11868 158300 11932
rect 158364 11930 158370 11932
rect 423765 11930 423831 11933
rect 158364 11928 423831 11930
rect 158364 11872 423770 11928
rect 423826 11872 423831 11928
rect 158364 11870 423831 11872
rect 158364 11868 158370 11870
rect 423765 11867 423831 11870
rect 162158 11732 162164 11796
rect 162228 11794 162234 11796
rect 473905 11794 473971 11797
rect 162228 11792 473971 11794
rect 162228 11736 473910 11792
rect 473966 11736 473971 11792
rect 162228 11734 473971 11736
rect 162228 11732 162234 11734
rect 473905 11731 473971 11734
rect 162342 11596 162348 11660
rect 162412 11658 162418 11660
rect 478137 11658 478203 11661
rect 162412 11656 478203 11658
rect 162412 11600 478142 11656
rect 478198 11600 478203 11656
rect 162412 11598 478203 11600
rect 162412 11596 162418 11598
rect 478137 11595 478203 11598
rect 110505 10570 110571 10573
rect 134190 10570 134196 10572
rect 110505 10568 134196 10570
rect 110505 10512 110510 10568
rect 110566 10512 134196 10568
rect 110505 10510 134196 10512
rect 110505 10507 110571 10510
rect 134190 10508 134196 10510
rect 134260 10508 134266 10572
rect 92473 10434 92539 10437
rect 133086 10434 133092 10436
rect 92473 10432 133092 10434
rect 92473 10376 92478 10432
rect 92534 10376 133092 10432
rect 92473 10374 133092 10376
rect 92473 10371 92539 10374
rect 133086 10372 133092 10374
rect 133156 10372 133162 10436
rect 149646 10372 149652 10436
rect 149716 10434 149722 10436
rect 316033 10434 316099 10437
rect 149716 10432 316099 10434
rect 149716 10376 316038 10432
rect 316094 10376 316099 10432
rect 149716 10374 316099 10376
rect 149716 10372 149722 10374
rect 316033 10371 316099 10374
rect 74993 10298 75059 10301
rect 131246 10298 131252 10300
rect 74993 10296 131252 10298
rect 74993 10240 74998 10296
rect 75054 10240 131252 10296
rect 74993 10238 131252 10240
rect 74993 10235 75059 10238
rect 131246 10236 131252 10238
rect 131316 10236 131322 10300
rect 158478 10236 158484 10300
rect 158548 10298 158554 10300
rect 420913 10298 420979 10301
rect 158548 10296 420979 10298
rect 158548 10240 420918 10296
rect 420974 10240 420979 10296
rect 158548 10238 420979 10240
rect 158548 10236 158554 10238
rect 420913 10235 420979 10238
rect 145598 9556 145604 9620
rect 145668 9618 145674 9620
rect 265341 9618 265407 9621
rect 145668 9616 265407 9618
rect 145668 9560 265346 9616
rect 265402 9560 265407 9616
rect 145668 9558 265407 9560
rect 145668 9556 145674 9558
rect 265341 9555 265407 9558
rect 147070 9420 147076 9484
rect 147140 9482 147146 9484
rect 281901 9482 281967 9485
rect 147140 9480 281967 9482
rect 147140 9424 281906 9480
rect 281962 9424 281967 9480
rect 147140 9422 281967 9424
rect 147140 9420 147146 9422
rect 281901 9419 281967 9422
rect 148726 9284 148732 9348
rect 148796 9346 148802 9348
rect 299657 9346 299723 9349
rect 148796 9344 299723 9346
rect 148796 9288 299662 9344
rect 299718 9288 299723 9344
rect 148796 9286 299723 9288
rect 148796 9284 148802 9286
rect 299657 9283 299723 9286
rect 57237 9210 57303 9213
rect 130326 9210 130332 9212
rect 57237 9208 130332 9210
rect 57237 9152 57242 9208
rect 57298 9152 130332 9208
rect 57237 9150 130332 9152
rect 57237 9147 57303 9150
rect 130326 9148 130332 9150
rect 130396 9148 130402 9212
rect 149830 9148 149836 9212
rect 149900 9210 149906 9212
rect 315021 9210 315087 9213
rect 149900 9208 315087 9210
rect 149900 9152 315026 9208
rect 315082 9152 315087 9208
rect 149900 9150 315087 9152
rect 149900 9148 149906 9150
rect 315021 9147 315087 9150
rect 56041 9074 56107 9077
rect 129958 9074 129964 9076
rect 56041 9072 129964 9074
rect 56041 9016 56046 9072
rect 56102 9016 129964 9072
rect 56041 9014 129964 9016
rect 56041 9011 56107 9014
rect 129958 9012 129964 9014
rect 130028 9012 130034 9076
rect 160870 9012 160876 9076
rect 160940 9074 160946 9076
rect 456885 9074 456951 9077
rect 160940 9072 456951 9074
rect 160940 9016 456890 9072
rect 456946 9016 456951 9072
rect 160940 9014 456951 9016
rect 160940 9012 160946 9014
rect 456885 9011 456951 9014
rect 41873 8938 41939 8941
rect 128670 8938 128676 8940
rect 41873 8936 128676 8938
rect 41873 8880 41878 8936
rect 41934 8880 128676 8936
rect 41873 8878 128676 8880
rect 41873 8875 41939 8878
rect 128670 8876 128676 8878
rect 128740 8876 128746 8940
rect 161054 8876 161060 8940
rect 161124 8938 161130 8940
rect 459185 8938 459251 8941
rect 161124 8936 459251 8938
rect 161124 8880 459190 8936
rect 459246 8880 459251 8936
rect 161124 8878 459251 8880
rect 161124 8876 161130 8878
rect 459185 8875 459251 8878
rect 111609 7714 111675 7717
rect 134006 7714 134012 7716
rect 111609 7712 134012 7714
rect 111609 7656 111614 7712
rect 111670 7656 134012 7712
rect 111609 7654 134012 7656
rect 111609 7651 111675 7654
rect 134006 7652 134012 7654
rect 134076 7652 134082 7716
rect 109309 7578 109375 7581
rect 134374 7578 134380 7580
rect 109309 7576 134380 7578
rect 109309 7520 109314 7576
rect 109370 7520 134380 7576
rect 109309 7518 134380 7520
rect 109309 7515 109375 7518
rect 134374 7516 134380 7518
rect 134444 7516 134450 7580
rect 150014 7516 150020 7580
rect 150084 7578 150090 7580
rect 316217 7578 316283 7581
rect 150084 7576 316283 7578
rect 150084 7520 316222 7576
rect 316278 7520 316283 7576
rect 150084 7518 316283 7520
rect 150084 7516 150090 7518
rect 316217 7515 316283 7518
rect 147254 6836 147260 6900
rect 147324 6898 147330 6900
rect 280705 6898 280771 6901
rect 147324 6896 280771 6898
rect 147324 6840 280710 6896
rect 280766 6840 280771 6896
rect 147324 6838 280771 6840
rect 147324 6836 147330 6838
rect 280705 6835 280771 6838
rect 146886 6700 146892 6764
rect 146956 6762 146962 6764
rect 284293 6762 284359 6765
rect 146956 6760 284359 6762
rect 146956 6704 284298 6760
rect 284354 6704 284359 6760
rect 146956 6702 284359 6704
rect 146956 6700 146962 6702
rect 284293 6699 284359 6702
rect -960 6490 480 6580
rect 148358 6564 148364 6628
rect 148428 6626 148434 6628
rect 300761 6626 300827 6629
rect 148428 6624 300827 6626
rect 148428 6568 300766 6624
rect 300822 6568 300827 6624
rect 148428 6566 300827 6568
rect 148428 6564 148434 6566
rect 300761 6563 300827 6566
rect 580257 6626 580323 6629
rect 583520 6626 584960 6716
rect 580257 6624 584960 6626
rect 580257 6568 580262 6624
rect 580318 6568 584960 6624
rect 580257 6566 584960 6568
rect 580257 6563 580323 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 152406 6428 152412 6492
rect 152476 6490 152482 6492
rect 351637 6490 351703 6493
rect 152476 6488 351703 6490
rect 152476 6432 351642 6488
rect 351698 6432 351703 6488
rect 583520 6476 584960 6566
rect 152476 6430 351703 6432
rect 152476 6428 152482 6430
rect 351637 6427 351703 6430
rect 73797 6354 73863 6357
rect 131062 6354 131068 6356
rect 73797 6352 131068 6354
rect 73797 6296 73802 6352
rect 73858 6296 131068 6352
rect 73797 6294 131068 6296
rect 73797 6291 73863 6294
rect 131062 6292 131068 6294
rect 131132 6292 131138 6356
rect 160686 6292 160692 6356
rect 160756 6354 160762 6356
rect 460381 6354 460447 6357
rect 160756 6352 460447 6354
rect 160756 6296 460386 6352
rect 460442 6296 460447 6352
rect 160756 6294 460447 6296
rect 160756 6292 160762 6294
rect 460381 6291 460447 6294
rect 40677 6218 40743 6221
rect 128670 6218 128676 6220
rect 40677 6216 128676 6218
rect 40677 6160 40682 6216
rect 40738 6160 128676 6216
rect 40677 6158 128676 6160
rect 40677 6155 40743 6158
rect 128670 6156 128676 6158
rect 128740 6156 128746 6220
rect 168046 6156 168052 6220
rect 168116 6218 168122 6220
rect 549069 6218 549135 6221
rect 168116 6216 549135 6218
rect 168116 6160 549074 6216
rect 549130 6160 549135 6216
rect 168116 6158 549135 6160
rect 168116 6156 168122 6158
rect 549069 6155 549135 6158
rect 143390 6020 143396 6084
rect 143460 6082 143466 6084
rect 228725 6082 228791 6085
rect 143460 6080 228791 6082
rect 143460 6024 228730 6080
rect 228786 6024 228791 6080
rect 143460 6022 228791 6024
rect 143460 6020 143466 6022
rect 228725 6019 228791 6022
rect 166758 5068 166764 5132
rect 166828 5130 166834 5132
rect 529013 5130 529079 5133
rect 166828 5128 529079 5130
rect 166828 5072 529018 5128
rect 529074 5072 529079 5128
rect 166828 5070 529079 5072
rect 166828 5068 166834 5070
rect 529013 5067 529079 5070
rect 20621 4994 20687 4997
rect 127014 4994 127020 4996
rect 20621 4992 127020 4994
rect 20621 4936 20626 4992
rect 20682 4936 127020 4992
rect 20621 4934 127020 4936
rect 20621 4931 20687 4934
rect 127014 4932 127020 4934
rect 127084 4932 127090 4996
rect 139158 4932 139164 4996
rect 139228 4994 139234 4996
rect 154481 4994 154547 4997
rect 139228 4992 154547 4994
rect 139228 4936 154486 4992
rect 154542 4936 154547 4992
rect 139228 4934 154547 4936
rect 139228 4932 139234 4934
rect 154481 4931 154547 4934
rect 170990 4932 170996 4996
rect 171060 4994 171066 4996
rect 577405 4994 577471 4997
rect 171060 4992 577471 4994
rect 171060 4936 577410 4992
rect 577466 4936 577471 4992
rect 171060 4934 577471 4936
rect 171060 4932 171066 4934
rect 577405 4931 577471 4934
rect 4061 4858 4127 4861
rect 125910 4858 125916 4860
rect 4061 4856 125916 4858
rect 4061 4800 4066 4856
rect 4122 4800 125916 4856
rect 4061 4798 125916 4800
rect 4061 4795 4127 4798
rect 125910 4796 125916 4798
rect 125980 4796 125986 4860
rect 137870 4796 137876 4860
rect 137940 4858 137946 4860
rect 158897 4858 158963 4861
rect 137940 4856 158963 4858
rect 137940 4800 158902 4856
rect 158958 4800 158963 4856
rect 137940 4798 158963 4800
rect 137940 4796 137946 4798
rect 158897 4795 158963 4798
rect 170806 4796 170812 4860
rect 170876 4858 170882 4860
rect 583385 4858 583451 4861
rect 170876 4856 583451 4858
rect 170876 4800 583390 4856
rect 583446 4800 583451 4856
rect 170876 4798 583451 4800
rect 170876 4796 170882 4798
rect 583385 4795 583451 4798
rect 161565 3906 161631 3909
rect 469857 3906 469923 3909
rect 161565 3904 469923 3906
rect 161565 3848 161570 3904
rect 161626 3848 469862 3904
rect 469918 3848 469923 3904
rect 161565 3846 469923 3848
rect 161565 3843 161631 3846
rect 469857 3843 469923 3846
rect 162526 3708 162532 3772
rect 162596 3770 162602 3772
rect 473445 3770 473511 3773
rect 162596 3768 473511 3770
rect 162596 3712 473450 3768
rect 473506 3712 473511 3768
rect 162596 3710 473511 3712
rect 162596 3708 162602 3710
rect 473445 3707 473511 3710
rect 162710 3572 162716 3636
rect 162780 3634 162786 3636
rect 476941 3634 477007 3637
rect 162780 3632 477007 3634
rect 162780 3576 476946 3632
rect 477002 3576 477007 3632
rect 162780 3574 477007 3576
rect 162780 3572 162786 3574
rect 476941 3571 477007 3574
rect 136398 3436 136404 3500
rect 136468 3498 136474 3500
rect 161289 3498 161355 3501
rect 136468 3496 161355 3498
rect 136468 3440 161294 3496
rect 161350 3440 161355 3496
rect 136468 3438 161355 3440
rect 136468 3436 136474 3438
rect 161289 3435 161355 3438
rect 170397 3498 170463 3501
rect 491109 3498 491175 3501
rect 170397 3496 491175 3498
rect 170397 3440 170402 3496
rect 170458 3440 491114 3496
rect 491170 3440 491175 3496
rect 170397 3438 491175 3440
rect 170397 3435 170463 3438
rect 491109 3435 491175 3438
rect 127566 3300 127572 3364
rect 127636 3362 127642 3364
rect 475745 3362 475811 3365
rect 127636 3360 475811 3362
rect 127636 3304 475750 3360
rect 475806 3304 475811 3360
rect 127636 3302 475811 3304
rect 127636 3300 127642 3302
rect 475745 3299 475811 3302
<< via3 >>
rect 125732 79906 125736 79932
rect 125736 79906 125792 79932
rect 125792 79906 125796 79932
rect 125732 79868 125796 79906
rect 126652 79868 126716 79932
rect 127020 79868 127084 79932
rect 127940 79906 127944 79932
rect 127944 79906 128000 79932
rect 128000 79906 128004 79932
rect 127940 79868 128004 79906
rect 126284 79792 126348 79796
rect 126284 79736 126288 79792
rect 126288 79736 126344 79792
rect 126344 79736 126348 79792
rect 126284 79732 126348 79736
rect 145420 80140 145484 80204
rect 140452 80004 140516 80068
rect 128492 79868 128556 79932
rect 129412 79868 129476 79932
rect 128860 79792 128924 79796
rect 128860 79736 128864 79792
rect 128864 79736 128920 79792
rect 128920 79736 128924 79792
rect 128860 79732 128924 79736
rect 130332 79906 130336 79932
rect 130336 79906 130392 79932
rect 130392 79906 130396 79932
rect 130332 79868 130396 79906
rect 130700 79868 130764 79932
rect 129964 79732 130028 79796
rect 131436 79792 131500 79796
rect 131436 79736 131440 79792
rect 131440 79736 131496 79792
rect 131496 79736 131500 79792
rect 131436 79732 131500 79736
rect 133460 79868 133524 79932
rect 135668 79868 135732 79932
rect 135300 79792 135364 79796
rect 135300 79736 135350 79792
rect 135350 79736 135364 79792
rect 135300 79732 135364 79736
rect 135484 79792 135548 79796
rect 135484 79736 135534 79792
rect 135534 79736 135548 79792
rect 135484 79732 135548 79736
rect 136588 79906 136592 79932
rect 136592 79906 136648 79932
rect 136648 79906 136652 79932
rect 136588 79868 136652 79906
rect 136956 79906 136960 79932
rect 136960 79906 137016 79932
rect 137016 79906 137020 79932
rect 136956 79868 137020 79906
rect 137692 79868 137756 79932
rect 138796 79868 138860 79932
rect 156276 80140 156340 80204
rect 157564 80004 157628 80068
rect 136404 79732 136468 79796
rect 139164 79656 139228 79660
rect 139900 79732 139964 79796
rect 139164 79600 139178 79656
rect 139178 79600 139228 79656
rect 139164 79596 139228 79600
rect 140084 79596 140148 79660
rect 141372 79906 141376 79932
rect 141376 79906 141432 79932
rect 141432 79906 141436 79932
rect 141372 79868 141436 79906
rect 141924 79868 141988 79932
rect 142292 79928 142356 79932
rect 142292 79872 142296 79928
rect 142296 79872 142352 79928
rect 142352 79872 142356 79928
rect 142292 79868 142356 79872
rect 141004 79732 141068 79796
rect 143028 79868 143092 79932
rect 142844 79732 142908 79796
rect 143212 79732 143276 79796
rect 144132 79868 144196 79932
rect 144500 79656 144564 79660
rect 147076 79868 147140 79932
rect 144500 79600 144514 79656
rect 144514 79600 144564 79656
rect 144500 79596 144564 79600
rect 145788 79596 145852 79660
rect 146892 79596 146956 79660
rect 148548 79868 148612 79932
rect 149284 79928 149348 79932
rect 149284 79872 149288 79928
rect 149288 79872 149344 79928
rect 149344 79872 149348 79928
rect 149284 79868 149348 79872
rect 148732 79732 148796 79796
rect 150020 79868 150084 79932
rect 150020 79732 150084 79796
rect 151492 79868 151556 79932
rect 152044 79928 152108 79932
rect 152044 79872 152048 79928
rect 152048 79872 152104 79928
rect 152104 79872 152108 79928
rect 152044 79868 152108 79872
rect 152780 79906 152784 79932
rect 152784 79906 152840 79932
rect 152840 79906 152844 79932
rect 152780 79868 152844 79906
rect 151676 79596 151740 79660
rect 153332 79868 153396 79932
rect 153884 79906 153888 79932
rect 153888 79906 153944 79932
rect 153944 79906 153948 79932
rect 153884 79868 153948 79906
rect 152964 79732 153028 79796
rect 154068 79732 154132 79796
rect 154436 79732 154500 79796
rect 155724 79868 155788 79932
rect 156092 79928 156156 79932
rect 156092 79872 156096 79928
rect 156096 79872 156152 79928
rect 156152 79872 156156 79928
rect 156092 79868 156156 79872
rect 156460 79906 156464 79932
rect 156464 79906 156520 79932
rect 156520 79906 156524 79932
rect 156460 79868 156524 79906
rect 158852 80004 158916 80068
rect 166580 80140 166644 80204
rect 157196 79868 157260 79932
rect 155908 79732 155972 79796
rect 153884 79656 153948 79660
rect 153884 79600 153934 79656
rect 153934 79600 153948 79656
rect 153884 79596 153948 79600
rect 154252 79656 154316 79660
rect 154252 79600 154266 79656
rect 154266 79600 154316 79656
rect 154252 79596 154316 79600
rect 157012 79732 157076 79796
rect 159772 79928 159836 79932
rect 159772 79872 159776 79928
rect 159776 79872 159832 79928
rect 159832 79872 159836 79928
rect 157932 79792 157996 79796
rect 157932 79736 157936 79792
rect 157936 79736 157992 79792
rect 157992 79736 157996 79792
rect 157932 79732 157996 79736
rect 158300 79732 158364 79796
rect 158116 79596 158180 79660
rect 159772 79868 159836 79872
rect 159404 79770 159408 79796
rect 159408 79770 159464 79796
rect 159464 79770 159468 79796
rect 159404 79732 159468 79770
rect 160140 79732 160204 79796
rect 159036 79596 159100 79660
rect 160876 79868 160940 79932
rect 161428 79906 161432 79932
rect 161432 79906 161488 79932
rect 161488 79906 161492 79932
rect 161428 79868 161492 79906
rect 160692 79732 160756 79796
rect 161796 79928 161860 79932
rect 161796 79872 161800 79928
rect 161800 79872 161856 79928
rect 161856 79872 161860 79928
rect 161796 79868 161860 79872
rect 161980 79732 162044 79796
rect 162716 79906 162720 79932
rect 162720 79906 162776 79932
rect 162776 79906 162780 79932
rect 162716 79868 162780 79906
rect 165476 79868 165540 79932
rect 166212 79868 166276 79932
rect 166764 79868 166828 79932
rect 168052 79868 168116 79932
rect 169156 79868 169220 79932
rect 162164 79596 162228 79660
rect 162716 79596 162780 79660
rect 167316 79732 167380 79796
rect 167684 79732 167748 79796
rect 165292 79596 165356 79660
rect 166028 79596 166092 79660
rect 169524 79732 169588 79796
rect 170076 79928 170140 79932
rect 170076 79872 170080 79928
rect 170080 79872 170136 79928
rect 170136 79872 170140 79928
rect 170076 79868 170140 79872
rect 170628 79868 170692 79932
rect 170996 79928 171060 79932
rect 170996 79872 171000 79928
rect 171000 79872 171056 79928
rect 171056 79872 171060 79928
rect 170996 79868 171060 79872
rect 171548 79868 171612 79932
rect 172652 79868 172716 79932
rect 173204 80004 173268 80068
rect 173572 80004 173636 80068
rect 170444 79732 170508 79796
rect 168972 79596 169036 79660
rect 171916 79656 171980 79660
rect 171916 79600 171930 79656
rect 171930 79600 171980 79656
rect 171916 79596 171980 79600
rect 172100 79596 172164 79660
rect 173388 79188 173452 79252
rect 170996 79112 171060 79116
rect 170996 79056 171010 79112
rect 171010 79056 171060 79112
rect 170996 79052 171060 79056
rect 125732 78704 125796 78708
rect 125732 78648 125746 78704
rect 125746 78648 125796 78704
rect 125732 78644 125796 78648
rect 125916 78704 125980 78708
rect 125916 78648 125930 78704
rect 125930 78648 125980 78704
rect 125916 78644 125980 78648
rect 126284 78644 126348 78708
rect 126652 78644 126716 78708
rect 127572 78644 127636 78708
rect 156276 78644 156340 78708
rect 156644 78704 156708 78708
rect 156644 78648 156694 78704
rect 156694 78648 156708 78704
rect 156644 78644 156708 78648
rect 157380 78644 157444 78708
rect 169708 78840 169772 78844
rect 169708 78784 169722 78840
rect 169722 78784 169772 78840
rect 169708 78780 169772 78784
rect 127940 78432 128004 78436
rect 127940 78376 127990 78432
rect 127990 78376 128004 78432
rect 127940 78372 128004 78376
rect 128676 78432 128740 78436
rect 128676 78376 128726 78432
rect 128726 78376 128740 78432
rect 128676 78372 128740 78376
rect 129412 78432 129476 78436
rect 129412 78376 129426 78432
rect 129426 78376 129476 78432
rect 129412 78372 129476 78376
rect 129780 78432 129844 78436
rect 129780 78376 129794 78432
rect 129794 78376 129844 78432
rect 129780 78372 129844 78376
rect 130332 78372 130396 78436
rect 131620 78372 131684 78436
rect 135484 78432 135548 78436
rect 135484 78376 135534 78432
rect 135534 78376 135548 78432
rect 135484 78372 135548 78376
rect 136588 78432 136652 78436
rect 136588 78376 136602 78432
rect 136602 78376 136652 78432
rect 136588 78372 136652 78376
rect 137876 78432 137940 78436
rect 137876 78376 137926 78432
rect 137926 78376 137940 78432
rect 137876 78372 137940 78376
rect 138980 78372 139044 78436
rect 143396 78432 143460 78436
rect 143396 78376 143410 78432
rect 143410 78376 143460 78432
rect 143396 78372 143460 78376
rect 144684 78432 144748 78436
rect 144684 78376 144698 78432
rect 144698 78376 144748 78432
rect 144684 78372 144748 78376
rect 147260 78372 147324 78436
rect 148364 78372 148428 78436
rect 149284 78372 149348 78436
rect 149836 78372 149900 78436
rect 152412 78372 152476 78436
rect 157564 78372 157628 78436
rect 157932 78372 157996 78436
rect 165108 78372 165172 78436
rect 166396 78372 166460 78436
rect 170996 78372 171060 78436
rect 130332 78236 130396 78300
rect 131068 78236 131132 78300
rect 135668 78236 135732 78300
rect 138612 78236 138676 78300
rect 140452 78296 140516 78300
rect 140452 78240 140466 78296
rect 140466 78240 140516 78296
rect 140452 78236 140516 78240
rect 148364 78236 148428 78300
rect 149468 78236 149532 78300
rect 152596 78236 152660 78300
rect 154068 78236 154132 78300
rect 158300 78236 158364 78300
rect 159404 78236 159468 78300
rect 159772 78236 159836 78300
rect 136956 78100 137020 78164
rect 141372 78100 141436 78164
rect 148548 78100 148612 78164
rect 151308 78100 151372 78164
rect 152044 78100 152108 78164
rect 153884 78100 153948 78164
rect 160692 78160 160756 78164
rect 160692 78104 160742 78160
rect 160742 78104 160756 78160
rect 160692 78100 160756 78104
rect 161796 78100 161860 78164
rect 170812 78296 170876 78300
rect 170812 78240 170826 78296
rect 170826 78240 170876 78296
rect 170812 78236 170876 78240
rect 131252 78024 131316 78028
rect 131252 77968 131302 78024
rect 131302 77968 131316 78024
rect 131252 77964 131316 77968
rect 133092 77964 133156 78028
rect 134012 77964 134076 78028
rect 140636 78024 140700 78028
rect 140636 77968 140650 78024
rect 140650 77968 140700 78024
rect 140636 77964 140700 77968
rect 142292 77964 142356 78028
rect 148916 77964 148980 78028
rect 153332 77964 153396 78028
rect 156092 78024 156156 78028
rect 156092 77968 156142 78024
rect 156142 77968 156156 78024
rect 156092 77964 156156 77968
rect 157748 77964 157812 78028
rect 171732 78100 171796 78164
rect 171916 78100 171980 78164
rect 168052 78024 168116 78028
rect 168052 77968 168066 78024
rect 168066 77968 168116 78024
rect 168052 77964 168116 77968
rect 169340 77964 169404 78028
rect 133276 77828 133340 77892
rect 134196 77828 134260 77892
rect 139900 77888 139964 77892
rect 139900 77832 139950 77888
rect 139950 77832 139964 77888
rect 139900 77828 139964 77832
rect 154068 77888 154132 77892
rect 154068 77832 154082 77888
rect 154082 77832 154132 77888
rect 154068 77828 154132 77832
rect 162532 77828 162596 77892
rect 164924 77828 164988 77892
rect 165476 77888 165540 77892
rect 165476 77832 165526 77888
rect 165526 77832 165540 77888
rect 165476 77828 165540 77832
rect 130700 77692 130764 77756
rect 156460 77692 156524 77756
rect 172100 77692 172164 77756
rect 145236 77556 145300 77620
rect 160692 77420 160756 77484
rect 162348 77420 162412 77484
rect 165476 77420 165540 77484
rect 166212 77420 166276 77484
rect 167868 77556 167932 77620
rect 171916 77420 171980 77484
rect 125548 77284 125612 77348
rect 126100 77284 126164 77348
rect 166212 77284 166276 77348
rect 167316 77284 167380 77348
rect 168052 77284 168116 77348
rect 170076 77284 170140 77348
rect 171180 77284 171244 77348
rect 172284 77284 172348 77348
rect 130148 77012 130212 77076
rect 158484 77012 158548 77076
rect 161428 77012 161492 77076
rect 142108 76876 142172 76940
rect 166028 76528 166092 76532
rect 166028 76472 166078 76528
rect 166078 76472 166092 76528
rect 166028 76468 166092 76472
rect 169708 76468 169772 76532
rect 170996 76332 171060 76396
rect 170628 76196 170692 76260
rect 163452 75924 163516 75988
rect 138612 75788 138676 75852
rect 151676 75652 151740 75716
rect 133460 75516 133524 75580
rect 151308 75516 151372 75580
rect 157196 75516 157260 75580
rect 131436 75380 131500 75444
rect 155724 75380 155788 75444
rect 125548 75244 125612 75308
rect 134380 75244 134444 75308
rect 135668 75244 135732 75308
rect 158300 75244 158364 75308
rect 161060 75304 161124 75308
rect 161060 75248 161110 75304
rect 161110 75248 161124 75304
rect 161060 75244 161124 75248
rect 161980 75244 162044 75308
rect 162348 75244 162412 75308
rect 163636 75244 163700 75308
rect 125732 75108 125796 75172
rect 135300 75108 135364 75172
rect 160140 75108 160204 75172
rect 170444 75108 170508 75172
rect 169156 74972 169220 75036
rect 140084 74428 140148 74492
rect 142844 74292 142908 74356
rect 144684 74156 144748 74220
rect 131620 74020 131684 74084
rect 155908 74020 155972 74084
rect 157012 74020 157076 74084
rect 130148 73884 130212 73948
rect 156828 73884 156892 73948
rect 129780 73748 129844 73812
rect 156644 72524 156708 72588
rect 148916 72388 148980 72452
rect 151492 71028 151556 71092
rect 138796 68444 138860 68508
rect 140268 68308 140332 68372
rect 152964 68172 153028 68236
rect 166212 66948 166276 67012
rect 167684 66812 167748 66876
rect 163452 65452 163516 65516
rect 164924 64092 164988 64156
rect 145236 62732 145300 62796
rect 172284 61372 172348 61436
rect 144500 58516 144564 58580
rect 152596 51716 152660 51780
rect 172100 48860 172164 48924
rect 171916 47500 171980 47564
rect 133276 44780 133340 44844
rect 171732 42060 171796 42124
rect 153884 35124 153948 35188
rect 140452 34036 140516 34100
rect 143028 33900 143092 33964
rect 145420 33764 145484 33828
rect 138980 32540 139044 32604
rect 165108 32404 165172 32468
rect 149468 29820 149532 29884
rect 152780 29684 152844 29748
rect 169524 29548 169588 29612
rect 140636 25468 140700 25532
rect 135668 22612 135732 22676
rect 157932 22612 157996 22676
rect 166396 21252 166460 21316
rect 144132 20028 144196 20092
rect 128860 19892 128924 19956
rect 137692 19892 137756 19956
rect 165292 19892 165356 19956
rect 167868 18532 167932 18596
rect 141004 17580 141068 17644
rect 148548 17444 148612 17508
rect 158116 17308 158180 17372
rect 163636 17172 163700 17236
rect 154068 15812 154132 15876
rect 158852 14724 158916 14788
rect 159036 14588 159100 14652
rect 165476 14452 165540 14516
rect 143212 13364 143276 13428
rect 154436 13228 154500 13292
rect 154252 13092 154316 13156
rect 166580 12956 166644 13020
rect 158300 11868 158364 11932
rect 162164 11732 162228 11796
rect 162348 11596 162412 11660
rect 134196 10508 134260 10572
rect 133092 10372 133156 10436
rect 149652 10372 149716 10436
rect 131252 10236 131316 10300
rect 158484 10236 158548 10300
rect 145604 9556 145668 9620
rect 147076 9420 147140 9484
rect 148732 9284 148796 9348
rect 130332 9148 130396 9212
rect 149836 9148 149900 9212
rect 129964 9012 130028 9076
rect 160876 9012 160940 9076
rect 128676 8876 128740 8940
rect 161060 8876 161124 8940
rect 134012 7652 134076 7716
rect 134380 7516 134444 7580
rect 150020 7516 150084 7580
rect 147260 6836 147324 6900
rect 146892 6700 146956 6764
rect 148364 6564 148428 6628
rect 152412 6428 152476 6492
rect 131068 6292 131132 6356
rect 160692 6292 160756 6356
rect 128676 6156 128740 6220
rect 168052 6156 168116 6220
rect 143396 6020 143460 6084
rect 166764 5068 166828 5132
rect 127020 4932 127084 4996
rect 139164 4932 139228 4996
rect 170996 4932 171060 4996
rect 125916 4796 125980 4860
rect 137876 4796 137940 4860
rect 170812 4796 170876 4860
rect 162532 3708 162596 3772
rect 162716 3572 162780 3636
rect 136404 3436 136468 3500
rect 127572 3300 127636 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 214954 69914 250398
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 205954 96914 241398
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 246454 101414 281898
rect 100794 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 101414 246454
rect 100794 246134 101414 246218
rect 100794 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 101414 246134
rect 100794 210454 101414 245898
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100794 174454 101414 209898
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 214954 105914 250398
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 259954 114914 295398
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 223954 114914 259398
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114294 115954 114914 151398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 228454 119414 263898
rect 118794 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 119414 228454
rect 118794 228134 119414 228218
rect 118794 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 119414 228134
rect 118794 192454 119414 227898
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 142000 119414 155898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 232954 123914 268398
rect 123294 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 123914 232954
rect 123294 232634 123914 232718
rect 123294 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 123914 232634
rect 123294 196954 123914 232398
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 142000 123914 160398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 142000 128414 164898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 241954 132914 277398
rect 132294 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 132914 241954
rect 132294 241634 132914 241718
rect 132294 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 132914 241634
rect 132294 205954 132914 241398
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 132294 169954 132914 205398
rect 132294 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 132914 169954
rect 132294 169634 132914 169718
rect 132294 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 132914 169634
rect 132294 142000 132914 169398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 246454 137414 281898
rect 136794 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 137414 246454
rect 136794 246134 137414 246218
rect 136794 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 137414 246134
rect 136794 210454 137414 245898
rect 136794 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 137414 210454
rect 136794 210134 137414 210218
rect 136794 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 137414 210134
rect 136794 174454 137414 209898
rect 136794 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 137414 174454
rect 136794 174134 137414 174218
rect 136794 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 137414 174134
rect 136794 142000 137414 173898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 214954 141914 250398
rect 141294 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 141914 214954
rect 141294 214634 141914 214718
rect 141294 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 141914 214634
rect 141294 178954 141914 214398
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 141294 142954 141914 178398
rect 141294 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 141914 142954
rect 141294 142634 141914 142718
rect 141294 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 141914 142634
rect 141294 142000 141914 142398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 142000 146414 146898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 223954 150914 259398
rect 150294 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 150914 223954
rect 150294 223634 150914 223718
rect 150294 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 150914 223634
rect 150294 187954 150914 223398
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 150294 151954 150914 187398
rect 150294 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 150914 151954
rect 150294 151634 150914 151718
rect 150294 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 150914 151634
rect 150294 142000 150914 151398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 228454 155414 263898
rect 154794 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 155414 228454
rect 154794 228134 155414 228218
rect 154794 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 155414 228134
rect 154794 192454 155414 227898
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154794 156454 155414 191898
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154794 142000 155414 155898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 232954 159914 268398
rect 159294 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 159914 232954
rect 159294 232634 159914 232718
rect 159294 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 159914 232634
rect 159294 196954 159914 232398
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 159294 160954 159914 196398
rect 159294 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 159914 160954
rect 159294 160634 159914 160718
rect 159294 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 159914 160634
rect 159294 142000 159914 160398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 142000 164414 164898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 241954 168914 277398
rect 168294 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 168914 241954
rect 168294 241634 168914 241718
rect 168294 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 168914 241634
rect 168294 205954 168914 241398
rect 168294 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 168914 205954
rect 168294 205634 168914 205718
rect 168294 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 168914 205634
rect 168294 169954 168914 205398
rect 168294 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 168914 169954
rect 168294 169634 168914 169718
rect 168294 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 168914 169634
rect 168294 142000 168914 169398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 246454 173414 281898
rect 172794 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 173414 246454
rect 172794 246134 173414 246218
rect 172794 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 173414 246134
rect 172794 210454 173414 245898
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 172794 142000 173414 173898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 214954 177914 250398
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 142000 177914 142398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 142000 182414 146898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 223954 186914 259398
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 139568 115954 139888 115986
rect 139568 115718 139610 115954
rect 139846 115718 139888 115954
rect 139568 115634 139888 115718
rect 139568 115398 139610 115634
rect 139846 115398 139888 115634
rect 139568 115366 139888 115398
rect 170288 115954 170608 115986
rect 170288 115718 170330 115954
rect 170566 115718 170608 115954
rect 170288 115634 170608 115718
rect 170288 115398 170330 115634
rect 170566 115398 170608 115634
rect 170288 115366 170608 115398
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 124208 111454 124528 111486
rect 124208 111218 124250 111454
rect 124486 111218 124528 111454
rect 124208 111134 124528 111218
rect 124208 110898 124250 111134
rect 124486 110898 124528 111134
rect 124208 110866 124528 110898
rect 154928 111454 155248 111486
rect 154928 111218 154970 111454
rect 155206 111218 155248 111454
rect 154928 111134 155248 111218
rect 154928 110898 154970 111134
rect 155206 110898 155248 111134
rect 154928 110866 155248 110898
rect 145419 80204 145485 80205
rect 145419 80140 145420 80204
rect 145484 80140 145485 80204
rect 145419 80139 145485 80140
rect 156275 80204 156341 80205
rect 156275 80140 156276 80204
rect 156340 80140 156341 80204
rect 156275 80139 156341 80140
rect 166579 80204 166645 80205
rect 166579 80140 166580 80204
rect 166644 80140 166645 80204
rect 166579 80139 166645 80140
rect 140451 80068 140517 80069
rect 140451 80004 140452 80068
rect 140516 80004 140517 80068
rect 140451 80003 140517 80004
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 125731 79932 125797 79933
rect 125731 79868 125732 79932
rect 125796 79930 125797 79932
rect 126651 79932 126717 79933
rect 125796 79870 126162 79930
rect 125796 79868 125797 79870
rect 125731 79867 125797 79868
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 125731 78708 125797 78709
rect 125731 78644 125732 78708
rect 125796 78644 125797 78708
rect 125731 78643 125797 78644
rect 125915 78708 125981 78709
rect 125915 78644 125916 78708
rect 125980 78644 125981 78708
rect 125915 78643 125981 78644
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 48454 119414 78000
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 52954 123914 78000
rect 125547 77348 125613 77349
rect 125547 77284 125548 77348
rect 125612 77284 125613 77348
rect 125547 77283 125613 77284
rect 125550 75309 125610 77283
rect 125547 75308 125613 75309
rect 125547 75244 125548 75308
rect 125612 75244 125613 75308
rect 125547 75243 125613 75244
rect 125734 75173 125794 78643
rect 125731 75172 125797 75173
rect 125731 75108 125732 75172
rect 125796 75108 125797 75172
rect 125731 75107 125797 75108
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 125918 4861 125978 78643
rect 126102 77349 126162 79870
rect 126651 79868 126652 79932
rect 126716 79868 126717 79932
rect 126651 79867 126717 79868
rect 127019 79932 127085 79933
rect 127019 79868 127020 79932
rect 127084 79868 127085 79932
rect 127019 79867 127085 79868
rect 127939 79932 128005 79933
rect 127939 79868 127940 79932
rect 128004 79868 128005 79932
rect 127939 79867 128005 79868
rect 128491 79932 128557 79933
rect 128491 79868 128492 79932
rect 128556 79868 128557 79932
rect 128491 79867 128557 79868
rect 129411 79932 129477 79933
rect 129411 79868 129412 79932
rect 129476 79868 129477 79932
rect 129411 79867 129477 79868
rect 130331 79932 130397 79933
rect 130331 79868 130332 79932
rect 130396 79868 130397 79932
rect 130331 79867 130397 79868
rect 130699 79932 130765 79933
rect 130699 79868 130700 79932
rect 130764 79868 130765 79932
rect 130699 79867 130765 79868
rect 133459 79932 133525 79933
rect 133459 79868 133460 79932
rect 133524 79868 133525 79932
rect 133459 79867 133525 79868
rect 135667 79932 135733 79933
rect 135667 79868 135668 79932
rect 135732 79868 135733 79932
rect 135667 79867 135733 79868
rect 136587 79932 136653 79933
rect 136587 79868 136588 79932
rect 136652 79868 136653 79932
rect 136587 79867 136653 79868
rect 136955 79932 137021 79933
rect 136955 79868 136956 79932
rect 137020 79868 137021 79932
rect 136955 79867 137021 79868
rect 137691 79932 137757 79933
rect 137691 79868 137692 79932
rect 137756 79868 137757 79932
rect 137691 79867 137757 79868
rect 138795 79932 138861 79933
rect 138795 79868 138796 79932
rect 138860 79868 138861 79932
rect 138795 79867 138861 79868
rect 126283 79796 126349 79797
rect 126283 79732 126284 79796
rect 126348 79732 126349 79796
rect 126283 79731 126349 79732
rect 126286 78709 126346 79731
rect 126654 78709 126714 79867
rect 126283 78708 126349 78709
rect 126283 78644 126284 78708
rect 126348 78644 126349 78708
rect 126283 78643 126349 78644
rect 126651 78708 126717 78709
rect 126651 78644 126652 78708
rect 126716 78644 126717 78708
rect 126651 78643 126717 78644
rect 126099 77348 126165 77349
rect 126099 77284 126100 77348
rect 126164 77284 126165 77348
rect 126099 77283 126165 77284
rect 127022 4997 127082 79867
rect 127571 78708 127637 78709
rect 127571 78644 127572 78708
rect 127636 78644 127637 78708
rect 127571 78643 127637 78644
rect 127019 4996 127085 4997
rect 127019 4932 127020 4996
rect 127084 4932 127085 4996
rect 127019 4931 127085 4932
rect 125915 4860 125981 4861
rect 125915 4796 125916 4860
rect 125980 4796 125981 4860
rect 125915 4795 125981 4796
rect 127574 3365 127634 78643
rect 127942 78437 128002 79867
rect 127939 78436 128005 78437
rect 127939 78372 127940 78436
rect 128004 78372 128005 78436
rect 127939 78371 128005 78372
rect 127794 57454 128414 78000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127571 3364 127637 3365
rect 127571 3300 127572 3364
rect 127636 3300 127637 3364
rect 127571 3299 127637 3300
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 -4186 128414 20898
rect 128494 6930 128554 79867
rect 128859 79796 128925 79797
rect 128859 79732 128860 79796
rect 128924 79732 128925 79796
rect 128859 79731 128925 79732
rect 128675 78436 128741 78437
rect 128675 78372 128676 78436
rect 128740 78372 128741 78436
rect 128675 78371 128741 78372
rect 128678 8941 128738 78371
rect 128862 19957 128922 79731
rect 129414 78437 129474 79867
rect 129963 79796 130029 79797
rect 129963 79732 129964 79796
rect 130028 79732 130029 79796
rect 129963 79731 130029 79732
rect 129411 78436 129477 78437
rect 129411 78372 129412 78436
rect 129476 78372 129477 78436
rect 129411 78371 129477 78372
rect 129779 78436 129845 78437
rect 129779 78372 129780 78436
rect 129844 78372 129845 78436
rect 129779 78371 129845 78372
rect 129782 73813 129842 78371
rect 129779 73812 129845 73813
rect 129779 73748 129780 73812
rect 129844 73748 129845 73812
rect 129779 73747 129845 73748
rect 128859 19956 128925 19957
rect 128859 19892 128860 19956
rect 128924 19892 128925 19956
rect 128859 19891 128925 19892
rect 129966 9077 130026 79731
rect 130334 78437 130394 79867
rect 130331 78436 130397 78437
rect 130331 78372 130332 78436
rect 130396 78372 130397 78436
rect 130331 78371 130397 78372
rect 130331 78300 130397 78301
rect 130331 78236 130332 78300
rect 130396 78236 130397 78300
rect 130331 78235 130397 78236
rect 130147 77076 130213 77077
rect 130147 77012 130148 77076
rect 130212 77012 130213 77076
rect 130147 77011 130213 77012
rect 130150 73949 130210 77011
rect 130147 73948 130213 73949
rect 130147 73884 130148 73948
rect 130212 73884 130213 73948
rect 130147 73883 130213 73884
rect 130334 9213 130394 78235
rect 130702 77757 130762 79867
rect 131435 79796 131501 79797
rect 131435 79732 131436 79796
rect 131500 79732 131501 79796
rect 131435 79731 131501 79732
rect 131067 78300 131133 78301
rect 131067 78236 131068 78300
rect 131132 78236 131133 78300
rect 131067 78235 131133 78236
rect 130699 77756 130765 77757
rect 130699 77692 130700 77756
rect 130764 77692 130765 77756
rect 130699 77691 130765 77692
rect 130331 9212 130397 9213
rect 130331 9148 130332 9212
rect 130396 9148 130397 9212
rect 130331 9147 130397 9148
rect 129963 9076 130029 9077
rect 129963 9012 129964 9076
rect 130028 9012 130029 9076
rect 129963 9011 130029 9012
rect 128675 8940 128741 8941
rect 128675 8876 128676 8940
rect 128740 8876 128741 8940
rect 128675 8875 128741 8876
rect 128494 6870 128738 6930
rect 128678 6221 128738 6870
rect 131070 6357 131130 78235
rect 131251 78028 131317 78029
rect 131251 77964 131252 78028
rect 131316 77964 131317 78028
rect 131251 77963 131317 77964
rect 131254 10301 131314 77963
rect 131438 75445 131498 79731
rect 131619 78436 131685 78437
rect 131619 78372 131620 78436
rect 131684 78372 131685 78436
rect 131619 78371 131685 78372
rect 131435 75444 131501 75445
rect 131435 75380 131436 75444
rect 131500 75380 131501 75444
rect 131435 75379 131501 75380
rect 131622 74085 131682 78371
rect 133091 78028 133157 78029
rect 131619 74084 131685 74085
rect 131619 74020 131620 74084
rect 131684 74020 131685 74084
rect 131619 74019 131685 74020
rect 132294 61954 132914 78000
rect 133091 77964 133092 78028
rect 133156 77964 133157 78028
rect 133091 77963 133157 77964
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 131251 10300 131317 10301
rect 131251 10236 131252 10300
rect 131316 10236 131317 10300
rect 131251 10235 131317 10236
rect 131067 6356 131133 6357
rect 131067 6292 131068 6356
rect 131132 6292 131133 6356
rect 131067 6291 131133 6292
rect 128675 6220 128741 6221
rect 128675 6156 128676 6220
rect 128740 6156 128741 6220
rect 128675 6155 128741 6156
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 -5146 132914 25398
rect 133094 10437 133154 77963
rect 133275 77892 133341 77893
rect 133275 77828 133276 77892
rect 133340 77828 133341 77892
rect 133275 77827 133341 77828
rect 133278 44845 133338 77827
rect 133462 75581 133522 79867
rect 135299 79796 135365 79797
rect 135299 79732 135300 79796
rect 135364 79732 135365 79796
rect 135299 79731 135365 79732
rect 135483 79796 135549 79797
rect 135483 79732 135484 79796
rect 135548 79732 135549 79796
rect 135483 79731 135549 79732
rect 134011 78028 134077 78029
rect 134011 77964 134012 78028
rect 134076 77964 134077 78028
rect 134011 77963 134077 77964
rect 133459 75580 133525 75581
rect 133459 75516 133460 75580
rect 133524 75516 133525 75580
rect 133459 75515 133525 75516
rect 133275 44844 133341 44845
rect 133275 44780 133276 44844
rect 133340 44780 133341 44844
rect 133275 44779 133341 44780
rect 133091 10436 133157 10437
rect 133091 10372 133092 10436
rect 133156 10372 133157 10436
rect 133091 10371 133157 10372
rect 134014 7717 134074 77963
rect 134195 77892 134261 77893
rect 134195 77828 134196 77892
rect 134260 77828 134261 77892
rect 134195 77827 134261 77828
rect 134198 10573 134258 77827
rect 134379 75308 134445 75309
rect 134379 75244 134380 75308
rect 134444 75244 134445 75308
rect 134379 75243 134445 75244
rect 134195 10572 134261 10573
rect 134195 10508 134196 10572
rect 134260 10508 134261 10572
rect 134195 10507 134261 10508
rect 134011 7716 134077 7717
rect 134011 7652 134012 7716
rect 134076 7652 134077 7716
rect 134011 7651 134077 7652
rect 134382 7581 134442 75243
rect 135302 75173 135362 79731
rect 135486 78437 135546 79731
rect 135483 78436 135549 78437
rect 135483 78372 135484 78436
rect 135548 78372 135549 78436
rect 135483 78371 135549 78372
rect 135670 78301 135730 79867
rect 136403 79796 136469 79797
rect 136403 79732 136404 79796
rect 136468 79732 136469 79796
rect 136403 79731 136469 79732
rect 135667 78300 135733 78301
rect 135667 78236 135668 78300
rect 135732 78236 135733 78300
rect 135667 78235 135733 78236
rect 135667 75308 135733 75309
rect 135667 75244 135668 75308
rect 135732 75244 135733 75308
rect 135667 75243 135733 75244
rect 135299 75172 135365 75173
rect 135299 75108 135300 75172
rect 135364 75108 135365 75172
rect 135299 75107 135365 75108
rect 135670 22677 135730 75243
rect 135667 22676 135733 22677
rect 135667 22612 135668 22676
rect 135732 22612 135733 22676
rect 135667 22611 135733 22612
rect 134379 7580 134445 7581
rect 134379 7516 134380 7580
rect 134444 7516 134445 7580
rect 134379 7515 134445 7516
rect 136406 3501 136466 79731
rect 136590 78437 136650 79867
rect 136587 78436 136653 78437
rect 136587 78372 136588 78436
rect 136652 78372 136653 78436
rect 136587 78371 136653 78372
rect 136958 78165 137018 79867
rect 136955 78164 137021 78165
rect 136955 78100 136956 78164
rect 137020 78100 137021 78164
rect 136955 78099 137021 78100
rect 136794 66454 137414 78000
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136403 3500 136469 3501
rect 136403 3436 136404 3500
rect 136468 3436 136469 3500
rect 136403 3435 136469 3436
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 -6106 137414 29898
rect 137694 19957 137754 79867
rect 137875 78436 137941 78437
rect 137875 78372 137876 78436
rect 137940 78372 137941 78436
rect 137875 78371 137941 78372
rect 137691 19956 137757 19957
rect 137691 19892 137692 19956
rect 137756 19892 137757 19956
rect 137691 19891 137757 19892
rect 137878 4861 137938 78371
rect 138611 78300 138677 78301
rect 138611 78236 138612 78300
rect 138676 78236 138677 78300
rect 138611 78235 138677 78236
rect 138614 75853 138674 78235
rect 138611 75852 138677 75853
rect 138611 75788 138612 75852
rect 138676 75788 138677 75852
rect 138611 75787 138677 75788
rect 138798 68509 138858 79867
rect 139899 79796 139965 79797
rect 139899 79732 139900 79796
rect 139964 79732 139965 79796
rect 139899 79731 139965 79732
rect 139163 79660 139229 79661
rect 139163 79596 139164 79660
rect 139228 79596 139229 79660
rect 139163 79595 139229 79596
rect 138979 78436 139045 78437
rect 138979 78372 138980 78436
rect 139044 78372 139045 78436
rect 138979 78371 139045 78372
rect 138795 68508 138861 68509
rect 138795 68444 138796 68508
rect 138860 68444 138861 68508
rect 138795 68443 138861 68444
rect 138982 32605 139042 78371
rect 138979 32604 139045 32605
rect 138979 32540 138980 32604
rect 139044 32540 139045 32604
rect 138979 32539 139045 32540
rect 139166 4997 139226 79595
rect 139902 77893 139962 79731
rect 140083 79660 140149 79661
rect 140083 79596 140084 79660
rect 140148 79596 140149 79660
rect 140083 79595 140149 79596
rect 139899 77892 139965 77893
rect 139899 77828 139900 77892
rect 139964 77828 139965 77892
rect 139899 77827 139965 77828
rect 140086 74493 140146 79595
rect 140454 78434 140514 80003
rect 141371 79932 141437 79933
rect 141371 79868 141372 79932
rect 141436 79868 141437 79932
rect 141371 79867 141437 79868
rect 141923 79932 141989 79933
rect 141923 79868 141924 79932
rect 141988 79930 141989 79932
rect 142291 79932 142357 79933
rect 141988 79870 142170 79930
rect 141988 79868 141989 79870
rect 141923 79867 141989 79868
rect 141003 79796 141069 79797
rect 141003 79732 141004 79796
rect 141068 79732 141069 79796
rect 141003 79731 141069 79732
rect 140270 78374 140514 78434
rect 140083 74492 140149 74493
rect 140083 74428 140084 74492
rect 140148 74428 140149 74492
rect 140083 74427 140149 74428
rect 140270 68373 140330 78374
rect 140451 78300 140517 78301
rect 140451 78236 140452 78300
rect 140516 78236 140517 78300
rect 140451 78235 140517 78236
rect 140267 68372 140333 68373
rect 140267 68308 140268 68372
rect 140332 68308 140333 68372
rect 140267 68307 140333 68308
rect 140454 34101 140514 78235
rect 140635 78028 140701 78029
rect 140635 77964 140636 78028
rect 140700 77964 140701 78028
rect 140635 77963 140701 77964
rect 140451 34100 140517 34101
rect 140451 34036 140452 34100
rect 140516 34036 140517 34100
rect 140451 34035 140517 34036
rect 140638 25533 140698 77963
rect 140635 25532 140701 25533
rect 140635 25468 140636 25532
rect 140700 25468 140701 25532
rect 140635 25467 140701 25468
rect 141006 17645 141066 79731
rect 141374 78165 141434 79867
rect 141371 78164 141437 78165
rect 141371 78100 141372 78164
rect 141436 78100 141437 78164
rect 141371 78099 141437 78100
rect 141294 70954 141914 78000
rect 142110 76941 142170 79870
rect 142291 79868 142292 79932
rect 142356 79868 142357 79932
rect 142291 79867 142357 79868
rect 143027 79932 143093 79933
rect 143027 79868 143028 79932
rect 143092 79868 143093 79932
rect 143027 79867 143093 79868
rect 144131 79932 144197 79933
rect 144131 79868 144132 79932
rect 144196 79868 144197 79932
rect 144131 79867 144197 79868
rect 142294 78029 142354 79867
rect 142843 79796 142909 79797
rect 142843 79732 142844 79796
rect 142908 79732 142909 79796
rect 142843 79731 142909 79732
rect 142291 78028 142357 78029
rect 142291 77964 142292 78028
rect 142356 77964 142357 78028
rect 142291 77963 142357 77964
rect 142107 76940 142173 76941
rect 142107 76876 142108 76940
rect 142172 76876 142173 76940
rect 142107 76875 142173 76876
rect 142846 74357 142906 79731
rect 142843 74356 142909 74357
rect 142843 74292 142844 74356
rect 142908 74292 142909 74356
rect 142843 74291 142909 74292
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141003 17644 141069 17645
rect 141003 17580 141004 17644
rect 141068 17580 141069 17644
rect 141003 17579 141069 17580
rect 139163 4996 139229 4997
rect 139163 4932 139164 4996
rect 139228 4932 139229 4996
rect 139163 4931 139229 4932
rect 137875 4860 137941 4861
rect 137875 4796 137876 4860
rect 137940 4796 137941 4860
rect 137875 4795 137941 4796
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 -7066 141914 34398
rect 143030 33965 143090 79867
rect 143211 79796 143277 79797
rect 143211 79732 143212 79796
rect 143276 79732 143277 79796
rect 143211 79731 143277 79732
rect 143027 33964 143093 33965
rect 143027 33900 143028 33964
rect 143092 33900 143093 33964
rect 143027 33899 143093 33900
rect 143214 13429 143274 79731
rect 143395 78436 143461 78437
rect 143395 78372 143396 78436
rect 143460 78372 143461 78436
rect 143395 78371 143461 78372
rect 143211 13428 143277 13429
rect 143211 13364 143212 13428
rect 143276 13364 143277 13428
rect 143211 13363 143277 13364
rect 143398 6085 143458 78371
rect 144134 20093 144194 79867
rect 144499 79660 144565 79661
rect 144499 79596 144500 79660
rect 144564 79596 144565 79660
rect 144499 79595 144565 79596
rect 144502 58581 144562 79595
rect 144683 78436 144749 78437
rect 144683 78372 144684 78436
rect 144748 78372 144749 78436
rect 144683 78371 144749 78372
rect 144686 74221 144746 78371
rect 145235 77620 145301 77621
rect 145235 77556 145236 77620
rect 145300 77556 145301 77620
rect 145235 77555 145301 77556
rect 144683 74220 144749 74221
rect 144683 74156 144684 74220
rect 144748 74156 144749 74220
rect 144683 74155 144749 74156
rect 145238 62797 145298 77555
rect 145235 62796 145301 62797
rect 145235 62732 145236 62796
rect 145300 62732 145301 62796
rect 145235 62731 145301 62732
rect 144499 58580 144565 58581
rect 144499 58516 144500 58580
rect 144564 58516 144565 58580
rect 144499 58515 144565 58516
rect 145422 33829 145482 80139
rect 147075 79932 147141 79933
rect 147075 79868 147076 79932
rect 147140 79868 147141 79932
rect 148547 79932 148613 79933
rect 148547 79930 148548 79932
rect 147075 79867 147141 79868
rect 148366 79870 148548 79930
rect 145787 79660 145853 79661
rect 145787 79658 145788 79660
rect 145606 79598 145788 79658
rect 145419 33828 145485 33829
rect 145419 33764 145420 33828
rect 145484 33764 145485 33828
rect 145419 33763 145485 33764
rect 144131 20092 144197 20093
rect 144131 20028 144132 20092
rect 144196 20028 144197 20092
rect 144131 20027 144197 20028
rect 145606 9621 145666 79598
rect 145787 79596 145788 79598
rect 145852 79596 145853 79660
rect 145787 79595 145853 79596
rect 146891 79660 146957 79661
rect 146891 79596 146892 79660
rect 146956 79596 146957 79660
rect 146891 79595 146957 79596
rect 145794 75454 146414 78000
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145603 9620 145669 9621
rect 145603 9556 145604 9620
rect 145668 9556 145669 9620
rect 145603 9555 145669 9556
rect 143395 6084 143461 6085
rect 143395 6020 143396 6084
rect 143460 6020 143461 6084
rect 143395 6019 143461 6020
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 3454 146414 38898
rect 146894 6765 146954 79595
rect 147078 9485 147138 79867
rect 148366 78437 148426 79870
rect 148547 79868 148548 79870
rect 148612 79868 148613 79932
rect 148547 79867 148613 79868
rect 149283 79932 149349 79933
rect 149283 79868 149284 79932
rect 149348 79868 149349 79932
rect 149283 79867 149349 79868
rect 150019 79932 150085 79933
rect 150019 79868 150020 79932
rect 150084 79930 150085 79932
rect 151491 79932 151557 79933
rect 150084 79870 150266 79930
rect 150084 79868 150085 79870
rect 150019 79867 150085 79868
rect 148731 79796 148797 79797
rect 148731 79732 148732 79796
rect 148796 79732 148797 79796
rect 148731 79731 148797 79732
rect 147259 78436 147325 78437
rect 147259 78372 147260 78436
rect 147324 78372 147325 78436
rect 147259 78371 147325 78372
rect 148363 78436 148429 78437
rect 148363 78372 148364 78436
rect 148428 78372 148429 78436
rect 148363 78371 148429 78372
rect 147075 9484 147141 9485
rect 147075 9420 147076 9484
rect 147140 9420 147141 9484
rect 147075 9419 147141 9420
rect 147262 6901 147322 78371
rect 148363 78300 148429 78301
rect 148363 78236 148364 78300
rect 148428 78236 148429 78300
rect 148363 78235 148429 78236
rect 147259 6900 147325 6901
rect 147259 6836 147260 6900
rect 147324 6836 147325 6900
rect 147259 6835 147325 6836
rect 146891 6764 146957 6765
rect 146891 6700 146892 6764
rect 146956 6700 146957 6764
rect 146891 6699 146957 6700
rect 148366 6629 148426 78235
rect 148547 78164 148613 78165
rect 148547 78100 148548 78164
rect 148612 78100 148613 78164
rect 148547 78099 148613 78100
rect 148550 17509 148610 78099
rect 148547 17508 148613 17509
rect 148547 17444 148548 17508
rect 148612 17444 148613 17508
rect 148547 17443 148613 17444
rect 148734 9349 148794 79731
rect 149286 78437 149346 79867
rect 150019 79796 150085 79797
rect 150019 79794 150020 79796
rect 149654 79734 150020 79794
rect 149283 78436 149349 78437
rect 149283 78372 149284 78436
rect 149348 78372 149349 78436
rect 149283 78371 149349 78372
rect 149467 78300 149533 78301
rect 149467 78236 149468 78300
rect 149532 78236 149533 78300
rect 149467 78235 149533 78236
rect 148915 78028 148981 78029
rect 148915 77964 148916 78028
rect 148980 77964 148981 78028
rect 148915 77963 148981 77964
rect 148918 72453 148978 77963
rect 148915 72452 148981 72453
rect 148915 72388 148916 72452
rect 148980 72388 148981 72452
rect 148915 72387 148981 72388
rect 149470 29885 149530 78235
rect 149467 29884 149533 29885
rect 149467 29820 149468 29884
rect 149532 29820 149533 29884
rect 149467 29819 149533 29820
rect 149654 10437 149714 79734
rect 150019 79732 150020 79734
rect 150084 79732 150085 79796
rect 150019 79731 150085 79732
rect 150206 78570 150266 79870
rect 151491 79868 151492 79932
rect 151556 79868 151557 79932
rect 151491 79867 151557 79868
rect 152043 79932 152109 79933
rect 152043 79868 152044 79932
rect 152108 79868 152109 79932
rect 152043 79867 152109 79868
rect 152779 79932 152845 79933
rect 152779 79868 152780 79932
rect 152844 79868 152845 79932
rect 152779 79867 152845 79868
rect 153331 79932 153397 79933
rect 153331 79868 153332 79932
rect 153396 79868 153397 79932
rect 153331 79867 153397 79868
rect 153883 79932 153949 79933
rect 153883 79868 153884 79932
rect 153948 79868 153949 79932
rect 153883 79867 153949 79868
rect 155723 79932 155789 79933
rect 155723 79868 155724 79932
rect 155788 79868 155789 79932
rect 155723 79867 155789 79868
rect 156091 79932 156157 79933
rect 156091 79868 156092 79932
rect 156156 79868 156157 79932
rect 156091 79867 156157 79868
rect 150022 78510 150266 78570
rect 149835 78436 149901 78437
rect 149835 78372 149836 78436
rect 149900 78372 149901 78436
rect 149835 78371 149901 78372
rect 149651 10436 149717 10437
rect 149651 10372 149652 10436
rect 149716 10372 149717 10436
rect 149651 10371 149717 10372
rect 148731 9348 148797 9349
rect 148731 9284 148732 9348
rect 148796 9284 148797 9348
rect 148731 9283 148797 9284
rect 149838 9213 149898 78371
rect 149835 9212 149901 9213
rect 149835 9148 149836 9212
rect 149900 9148 149901 9212
rect 149835 9147 149901 9148
rect 150022 7581 150082 78510
rect 151307 78164 151373 78165
rect 151307 78100 151308 78164
rect 151372 78100 151373 78164
rect 151307 78099 151373 78100
rect 150294 43954 150914 78000
rect 151310 75581 151370 78099
rect 151307 75580 151373 75581
rect 151307 75516 151308 75580
rect 151372 75516 151373 75580
rect 151307 75515 151373 75516
rect 151494 71093 151554 79867
rect 151675 79660 151741 79661
rect 151675 79596 151676 79660
rect 151740 79596 151741 79660
rect 151675 79595 151741 79596
rect 151678 75717 151738 79595
rect 152046 78165 152106 79867
rect 152411 78436 152477 78437
rect 152411 78372 152412 78436
rect 152476 78372 152477 78436
rect 152411 78371 152477 78372
rect 152043 78164 152109 78165
rect 152043 78100 152044 78164
rect 152108 78100 152109 78164
rect 152043 78099 152109 78100
rect 151675 75716 151741 75717
rect 151675 75652 151676 75716
rect 151740 75652 151741 75716
rect 151675 75651 151741 75652
rect 151491 71092 151557 71093
rect 151491 71028 151492 71092
rect 151556 71028 151557 71092
rect 151491 71027 151557 71028
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150019 7580 150085 7581
rect 150019 7516 150020 7580
rect 150084 7516 150085 7580
rect 150019 7515 150085 7516
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 148363 6628 148429 6629
rect 148363 6564 148364 6628
rect 148428 6564 148429 6628
rect 148363 6563 148429 6564
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 -1306 150914 7398
rect 152414 6493 152474 78371
rect 152595 78300 152661 78301
rect 152595 78236 152596 78300
rect 152660 78236 152661 78300
rect 152595 78235 152661 78236
rect 152598 51781 152658 78235
rect 152595 51780 152661 51781
rect 152595 51716 152596 51780
rect 152660 51716 152661 51780
rect 152595 51715 152661 51716
rect 152782 29749 152842 79867
rect 152963 79796 153029 79797
rect 152963 79732 152964 79796
rect 153028 79732 153029 79796
rect 152963 79731 153029 79732
rect 152966 68237 153026 79731
rect 153334 78029 153394 79867
rect 153886 79661 153946 79867
rect 154067 79796 154133 79797
rect 154067 79732 154068 79796
rect 154132 79732 154133 79796
rect 154067 79731 154133 79732
rect 154435 79796 154501 79797
rect 154435 79732 154436 79796
rect 154500 79732 154501 79796
rect 154435 79731 154501 79732
rect 153883 79660 153949 79661
rect 153883 79596 153884 79660
rect 153948 79596 153949 79660
rect 153883 79595 153949 79596
rect 154070 78301 154130 79731
rect 154251 79660 154317 79661
rect 154251 79596 154252 79660
rect 154316 79596 154317 79660
rect 154251 79595 154317 79596
rect 154067 78300 154133 78301
rect 154067 78236 154068 78300
rect 154132 78236 154133 78300
rect 154067 78235 154133 78236
rect 153883 78164 153949 78165
rect 153883 78100 153884 78164
rect 153948 78100 153949 78164
rect 153883 78099 153949 78100
rect 153331 78028 153397 78029
rect 153331 77964 153332 78028
rect 153396 77964 153397 78028
rect 153331 77963 153397 77964
rect 152963 68236 153029 68237
rect 152963 68172 152964 68236
rect 153028 68172 153029 68236
rect 152963 68171 153029 68172
rect 153886 35189 153946 78099
rect 154067 77892 154133 77893
rect 154067 77828 154068 77892
rect 154132 77828 154133 77892
rect 154067 77827 154133 77828
rect 153883 35188 153949 35189
rect 153883 35124 153884 35188
rect 153948 35124 153949 35188
rect 153883 35123 153949 35124
rect 152779 29748 152845 29749
rect 152779 29684 152780 29748
rect 152844 29684 152845 29748
rect 152779 29683 152845 29684
rect 154070 15877 154130 77827
rect 154067 15876 154133 15877
rect 154067 15812 154068 15876
rect 154132 15812 154133 15876
rect 154067 15811 154133 15812
rect 154254 13157 154314 79595
rect 154438 13293 154498 79731
rect 154794 48454 155414 78000
rect 155726 75445 155786 79867
rect 155907 79796 155973 79797
rect 155907 79732 155908 79796
rect 155972 79732 155973 79796
rect 155907 79731 155973 79732
rect 155723 75444 155789 75445
rect 155723 75380 155724 75444
rect 155788 75380 155789 75444
rect 155723 75379 155789 75380
rect 155910 74085 155970 79731
rect 156094 78029 156154 79867
rect 156278 78709 156338 80139
rect 157563 80068 157629 80069
rect 157563 80004 157564 80068
rect 157628 80004 157629 80068
rect 157563 80003 157629 80004
rect 158851 80068 158917 80069
rect 158851 80004 158852 80068
rect 158916 80004 158917 80068
rect 158851 80003 158917 80004
rect 156459 79932 156525 79933
rect 156459 79868 156460 79932
rect 156524 79868 156525 79932
rect 157195 79932 157261 79933
rect 157195 79930 157196 79932
rect 156459 79867 156525 79868
rect 156830 79870 157196 79930
rect 156275 78708 156341 78709
rect 156275 78644 156276 78708
rect 156340 78644 156341 78708
rect 156275 78643 156341 78644
rect 156091 78028 156157 78029
rect 156091 77964 156092 78028
rect 156156 77964 156157 78028
rect 156091 77963 156157 77964
rect 156462 77757 156522 79867
rect 156643 78708 156709 78709
rect 156643 78644 156644 78708
rect 156708 78644 156709 78708
rect 156643 78643 156709 78644
rect 156459 77756 156525 77757
rect 156459 77692 156460 77756
rect 156524 77692 156525 77756
rect 156459 77691 156525 77692
rect 155907 74084 155973 74085
rect 155907 74020 155908 74084
rect 155972 74020 155973 74084
rect 155907 74019 155973 74020
rect 156646 72589 156706 78643
rect 156830 73949 156890 79870
rect 157195 79868 157196 79870
rect 157260 79868 157261 79932
rect 157195 79867 157261 79868
rect 157011 79796 157077 79797
rect 157011 79732 157012 79796
rect 157076 79732 157077 79796
rect 157011 79731 157077 79732
rect 157014 74085 157074 79731
rect 157379 78708 157445 78709
rect 157379 78644 157380 78708
rect 157444 78644 157445 78708
rect 157379 78643 157445 78644
rect 157382 75930 157442 78643
rect 157566 78437 157626 80003
rect 157931 79796 157997 79797
rect 157931 79732 157932 79796
rect 157996 79732 157997 79796
rect 157931 79731 157997 79732
rect 158299 79796 158365 79797
rect 158299 79732 158300 79796
rect 158364 79732 158365 79796
rect 158299 79731 158365 79732
rect 157934 78437 157994 79731
rect 158115 79660 158181 79661
rect 158115 79596 158116 79660
rect 158180 79596 158181 79660
rect 158115 79595 158181 79596
rect 157563 78436 157629 78437
rect 157563 78372 157564 78436
rect 157628 78372 157629 78436
rect 157563 78371 157629 78372
rect 157931 78436 157997 78437
rect 157931 78372 157932 78436
rect 157996 78372 157997 78436
rect 157931 78371 157997 78372
rect 157747 78028 157813 78029
rect 157747 77964 157748 78028
rect 157812 77964 157813 78028
rect 157747 77963 157813 77964
rect 157198 75870 157442 75930
rect 157198 75581 157258 75870
rect 157195 75580 157261 75581
rect 157195 75516 157196 75580
rect 157260 75516 157261 75580
rect 157195 75515 157261 75516
rect 157011 74084 157077 74085
rect 157011 74020 157012 74084
rect 157076 74020 157077 74084
rect 157011 74019 157077 74020
rect 156827 73948 156893 73949
rect 156827 73884 156828 73948
rect 156892 73884 156893 73948
rect 156827 73883 156893 73884
rect 156643 72588 156709 72589
rect 156643 72524 156644 72588
rect 156708 72524 156709 72588
rect 156643 72523 156709 72524
rect 157750 70410 157810 77963
rect 157750 70350 157994 70410
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154435 13292 154501 13293
rect 154435 13228 154436 13292
rect 154500 13228 154501 13292
rect 154435 13227 154501 13228
rect 154251 13156 154317 13157
rect 154251 13092 154252 13156
rect 154316 13092 154317 13156
rect 154251 13091 154317 13092
rect 154794 12454 155414 47898
rect 157934 22677 157994 70350
rect 157931 22676 157997 22677
rect 157931 22612 157932 22676
rect 157996 22612 157997 22676
rect 157931 22611 157997 22612
rect 158118 17373 158178 79595
rect 158302 78301 158362 79731
rect 158299 78300 158365 78301
rect 158299 78236 158300 78300
rect 158364 78236 158365 78300
rect 158299 78235 158365 78236
rect 158483 77076 158549 77077
rect 158483 77012 158484 77076
rect 158548 77012 158549 77076
rect 158483 77011 158549 77012
rect 158299 75308 158365 75309
rect 158299 75244 158300 75308
rect 158364 75244 158365 75308
rect 158299 75243 158365 75244
rect 158115 17372 158181 17373
rect 158115 17308 158116 17372
rect 158180 17308 158181 17372
rect 158115 17307 158181 17308
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 158302 11933 158362 75243
rect 152411 6492 152477 6493
rect 152411 6428 152412 6492
rect 152476 6428 152477 6492
rect 152411 6427 152477 6428
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 -2266 155414 11898
rect 158299 11932 158365 11933
rect 158299 11868 158300 11932
rect 158364 11868 158365 11932
rect 158299 11867 158365 11868
rect 158486 10301 158546 77011
rect 158854 14789 158914 80003
rect 159771 79932 159837 79933
rect 159771 79868 159772 79932
rect 159836 79868 159837 79932
rect 159771 79867 159837 79868
rect 160875 79932 160941 79933
rect 160875 79868 160876 79932
rect 160940 79868 160941 79932
rect 160875 79867 160941 79868
rect 161427 79932 161493 79933
rect 161427 79868 161428 79932
rect 161492 79868 161493 79932
rect 161427 79867 161493 79868
rect 161795 79932 161861 79933
rect 161795 79868 161796 79932
rect 161860 79868 161861 79932
rect 162715 79932 162781 79933
rect 162715 79930 162716 79932
rect 161795 79867 161861 79868
rect 162350 79870 162716 79930
rect 159403 79796 159469 79797
rect 159403 79732 159404 79796
rect 159468 79732 159469 79796
rect 159403 79731 159469 79732
rect 159035 79660 159101 79661
rect 159035 79596 159036 79660
rect 159100 79596 159101 79660
rect 159035 79595 159101 79596
rect 158851 14788 158917 14789
rect 158851 14724 158852 14788
rect 158916 14724 158917 14788
rect 158851 14723 158917 14724
rect 159038 14653 159098 79595
rect 159406 78301 159466 79731
rect 159774 78301 159834 79867
rect 160139 79796 160205 79797
rect 160139 79732 160140 79796
rect 160204 79732 160205 79796
rect 160139 79731 160205 79732
rect 160691 79796 160757 79797
rect 160691 79732 160692 79796
rect 160756 79732 160757 79796
rect 160691 79731 160757 79732
rect 159403 78300 159469 78301
rect 159403 78236 159404 78300
rect 159468 78236 159469 78300
rect 159403 78235 159469 78236
rect 159771 78300 159837 78301
rect 159771 78236 159772 78300
rect 159836 78236 159837 78300
rect 159771 78235 159837 78236
rect 159294 52954 159914 78000
rect 160142 75173 160202 79731
rect 160694 78165 160754 79731
rect 160691 78164 160757 78165
rect 160691 78100 160692 78164
rect 160756 78100 160757 78164
rect 160691 78099 160757 78100
rect 160691 77484 160757 77485
rect 160691 77420 160692 77484
rect 160756 77420 160757 77484
rect 160691 77419 160757 77420
rect 160139 75172 160205 75173
rect 160139 75108 160140 75172
rect 160204 75108 160205 75172
rect 160139 75107 160205 75108
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159035 14652 159101 14653
rect 159035 14588 159036 14652
rect 159100 14588 159101 14652
rect 159035 14587 159101 14588
rect 158483 10300 158549 10301
rect 158483 10236 158484 10300
rect 158548 10236 158549 10300
rect 158483 10235 158549 10236
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 -3226 159914 16398
rect 160694 6357 160754 77419
rect 160878 9077 160938 79867
rect 161430 77077 161490 79867
rect 161798 78165 161858 79867
rect 161979 79796 162045 79797
rect 161979 79732 161980 79796
rect 162044 79732 162045 79796
rect 161979 79731 162045 79732
rect 161795 78164 161861 78165
rect 161795 78100 161796 78164
rect 161860 78100 161861 78164
rect 161795 78099 161861 78100
rect 161427 77076 161493 77077
rect 161427 77012 161428 77076
rect 161492 77012 161493 77076
rect 161427 77011 161493 77012
rect 161982 75309 162042 79731
rect 162163 79660 162229 79661
rect 162163 79596 162164 79660
rect 162228 79596 162229 79660
rect 162163 79595 162229 79596
rect 161059 75308 161125 75309
rect 161059 75244 161060 75308
rect 161124 75244 161125 75308
rect 161059 75243 161125 75244
rect 161979 75308 162045 75309
rect 161979 75244 161980 75308
rect 162044 75244 162045 75308
rect 161979 75243 162045 75244
rect 160875 9076 160941 9077
rect 160875 9012 160876 9076
rect 160940 9012 160941 9076
rect 160875 9011 160941 9012
rect 161062 8941 161122 75243
rect 162166 11797 162226 79595
rect 162350 77485 162410 79870
rect 162715 79868 162716 79870
rect 162780 79868 162781 79932
rect 162715 79867 162781 79868
rect 165475 79932 165541 79933
rect 165475 79868 165476 79932
rect 165540 79868 165541 79932
rect 165475 79867 165541 79868
rect 166211 79932 166277 79933
rect 166211 79868 166212 79932
rect 166276 79868 166277 79932
rect 166211 79867 166277 79868
rect 162715 79660 162781 79661
rect 162715 79596 162716 79660
rect 162780 79596 162781 79660
rect 162715 79595 162781 79596
rect 165291 79660 165357 79661
rect 165291 79596 165292 79660
rect 165356 79596 165357 79660
rect 165291 79595 165357 79596
rect 162531 77892 162597 77893
rect 162531 77828 162532 77892
rect 162596 77828 162597 77892
rect 162531 77827 162597 77828
rect 162347 77484 162413 77485
rect 162347 77420 162348 77484
rect 162412 77420 162413 77484
rect 162347 77419 162413 77420
rect 162347 75308 162413 75309
rect 162347 75244 162348 75308
rect 162412 75244 162413 75308
rect 162347 75243 162413 75244
rect 162163 11796 162229 11797
rect 162163 11732 162164 11796
rect 162228 11732 162229 11796
rect 162163 11731 162229 11732
rect 162350 11661 162410 75243
rect 162347 11660 162413 11661
rect 162347 11596 162348 11660
rect 162412 11596 162413 11660
rect 162347 11595 162413 11596
rect 161059 8940 161125 8941
rect 161059 8876 161060 8940
rect 161124 8876 161125 8940
rect 161059 8875 161125 8876
rect 160691 6356 160757 6357
rect 160691 6292 160692 6356
rect 160756 6292 160757 6356
rect 160691 6291 160757 6292
rect 162534 3773 162594 77827
rect 162531 3772 162597 3773
rect 162531 3708 162532 3772
rect 162596 3708 162597 3772
rect 162531 3707 162597 3708
rect 162718 3637 162778 79595
rect 165107 78436 165173 78437
rect 165107 78372 165108 78436
rect 165172 78372 165173 78436
rect 165107 78371 165173 78372
rect 163451 75988 163517 75989
rect 163451 75924 163452 75988
rect 163516 75924 163517 75988
rect 163451 75923 163517 75924
rect 163454 65517 163514 75923
rect 163635 75308 163701 75309
rect 163635 75244 163636 75308
rect 163700 75244 163701 75308
rect 163635 75243 163701 75244
rect 163451 65516 163517 65517
rect 163451 65452 163452 65516
rect 163516 65452 163517 65516
rect 163451 65451 163517 65452
rect 163638 17237 163698 75243
rect 163794 57454 164414 78000
rect 164923 77892 164989 77893
rect 164923 77828 164924 77892
rect 164988 77828 164989 77892
rect 164923 77827 164989 77828
rect 164926 64157 164986 77827
rect 164923 64156 164989 64157
rect 164923 64092 164924 64156
rect 164988 64092 164989 64156
rect 164923 64091 164989 64092
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 165110 32469 165170 78371
rect 165107 32468 165173 32469
rect 165107 32404 165108 32468
rect 165172 32404 165173 32468
rect 165107 32403 165173 32404
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163635 17236 163701 17237
rect 163635 17172 163636 17236
rect 163700 17172 163701 17236
rect 163635 17171 163701 17172
rect 162715 3636 162781 3637
rect 162715 3572 162716 3636
rect 162780 3572 162781 3636
rect 162715 3571 162781 3572
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 -4186 164414 20898
rect 165294 19957 165354 79595
rect 165478 77893 165538 79867
rect 166027 79660 166093 79661
rect 166027 79596 166028 79660
rect 166092 79596 166093 79660
rect 166027 79595 166093 79596
rect 165475 77892 165541 77893
rect 165475 77828 165476 77892
rect 165540 77828 165541 77892
rect 165475 77827 165541 77828
rect 165475 77484 165541 77485
rect 165475 77420 165476 77484
rect 165540 77420 165541 77484
rect 165475 77419 165541 77420
rect 165291 19956 165357 19957
rect 165291 19892 165292 19956
rect 165356 19892 165357 19956
rect 165291 19891 165357 19892
rect 165478 14517 165538 77419
rect 166030 76533 166090 79595
rect 166214 77485 166274 79867
rect 166395 78436 166461 78437
rect 166395 78372 166396 78436
rect 166460 78372 166461 78436
rect 166395 78371 166461 78372
rect 166211 77484 166277 77485
rect 166211 77420 166212 77484
rect 166276 77420 166277 77484
rect 166211 77419 166277 77420
rect 166211 77348 166277 77349
rect 166211 77284 166212 77348
rect 166276 77284 166277 77348
rect 166211 77283 166277 77284
rect 166027 76532 166093 76533
rect 166027 76468 166028 76532
rect 166092 76468 166093 76532
rect 166027 76467 166093 76468
rect 166214 67013 166274 77283
rect 166211 67012 166277 67013
rect 166211 66948 166212 67012
rect 166276 66948 166277 67012
rect 166211 66947 166277 66948
rect 166398 21317 166458 78371
rect 166395 21316 166461 21317
rect 166395 21252 166396 21316
rect 166460 21252 166461 21316
rect 166395 21251 166461 21252
rect 165475 14516 165541 14517
rect 165475 14452 165476 14516
rect 165540 14452 165541 14516
rect 165475 14451 165541 14452
rect 166582 13021 166642 80139
rect 173203 80068 173269 80069
rect 173203 80004 173204 80068
rect 173268 80066 173269 80068
rect 173571 80068 173637 80069
rect 173571 80066 173572 80068
rect 173268 80006 173572 80066
rect 173268 80004 173269 80006
rect 173203 80003 173269 80004
rect 173571 80004 173572 80006
rect 173636 80004 173637 80068
rect 173571 80003 173637 80004
rect 186294 79954 186914 115398
rect 166763 79932 166829 79933
rect 166763 79868 166764 79932
rect 166828 79868 166829 79932
rect 166763 79867 166829 79868
rect 168051 79932 168117 79933
rect 168051 79868 168052 79932
rect 168116 79868 168117 79932
rect 168051 79867 168117 79868
rect 169155 79932 169221 79933
rect 169155 79868 169156 79932
rect 169220 79930 169221 79932
rect 170075 79932 170141 79933
rect 169220 79870 169402 79930
rect 169220 79868 169221 79870
rect 169155 79867 169221 79868
rect 166579 13020 166645 13021
rect 166579 12956 166580 13020
rect 166644 12956 166645 13020
rect 166579 12955 166645 12956
rect 166766 5133 166826 79867
rect 167315 79796 167381 79797
rect 167315 79732 167316 79796
rect 167380 79732 167381 79796
rect 167315 79731 167381 79732
rect 167683 79796 167749 79797
rect 167683 79732 167684 79796
rect 167748 79732 167749 79796
rect 167683 79731 167749 79732
rect 167318 77349 167378 79731
rect 167315 77348 167381 77349
rect 167315 77284 167316 77348
rect 167380 77284 167381 77348
rect 167315 77283 167381 77284
rect 167686 66877 167746 79731
rect 168054 78029 168114 79867
rect 168971 79660 169037 79661
rect 168971 79596 168972 79660
rect 169036 79658 169037 79660
rect 169036 79598 169218 79658
rect 169036 79596 169037 79598
rect 168971 79595 169037 79596
rect 168051 78028 168117 78029
rect 168051 77964 168052 78028
rect 168116 77964 168117 78028
rect 168051 77963 168117 77964
rect 167867 77620 167933 77621
rect 167867 77556 167868 77620
rect 167932 77556 167933 77620
rect 167867 77555 167933 77556
rect 167683 66876 167749 66877
rect 167683 66812 167684 66876
rect 167748 66812 167749 66876
rect 167683 66811 167749 66812
rect 167870 18597 167930 77555
rect 168051 77348 168117 77349
rect 168051 77284 168052 77348
rect 168116 77284 168117 77348
rect 168051 77283 168117 77284
rect 167867 18596 167933 18597
rect 167867 18532 167868 18596
rect 167932 18532 167933 18596
rect 167867 18531 167933 18532
rect 168054 6221 168114 77283
rect 168294 61954 168914 78000
rect 169158 75037 169218 79598
rect 169342 78029 169402 79870
rect 170075 79868 170076 79932
rect 170140 79868 170141 79932
rect 170075 79867 170141 79868
rect 170627 79932 170693 79933
rect 170627 79868 170628 79932
rect 170692 79868 170693 79932
rect 170627 79867 170693 79868
rect 170995 79932 171061 79933
rect 170995 79868 170996 79932
rect 171060 79868 171061 79932
rect 170995 79867 171061 79868
rect 171547 79932 171613 79933
rect 171547 79868 171548 79932
rect 171612 79930 171613 79932
rect 172651 79932 172717 79933
rect 171612 79870 172162 79930
rect 171612 79868 171613 79870
rect 171547 79867 171613 79868
rect 169523 79796 169589 79797
rect 169523 79732 169524 79796
rect 169588 79732 169589 79796
rect 169523 79731 169589 79732
rect 169339 78028 169405 78029
rect 169339 77964 169340 78028
rect 169404 77964 169405 78028
rect 169339 77963 169405 77964
rect 169155 75036 169221 75037
rect 169155 74972 169156 75036
rect 169220 74972 169221 75036
rect 169155 74971 169221 74972
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 169526 29613 169586 79731
rect 169707 78844 169773 78845
rect 169707 78780 169708 78844
rect 169772 78780 169773 78844
rect 169707 78779 169773 78780
rect 169710 76533 169770 78779
rect 170078 77349 170138 79867
rect 170443 79796 170509 79797
rect 170443 79732 170444 79796
rect 170508 79732 170509 79796
rect 170443 79731 170509 79732
rect 170075 77348 170141 77349
rect 170075 77284 170076 77348
rect 170140 77284 170141 77348
rect 170075 77283 170141 77284
rect 169707 76532 169773 76533
rect 169707 76468 169708 76532
rect 169772 76468 169773 76532
rect 169707 76467 169773 76468
rect 170446 75173 170506 79731
rect 170630 76261 170690 79867
rect 170998 79117 171058 79867
rect 172102 79661 172162 79870
rect 172651 79868 172652 79932
rect 172716 79930 172717 79932
rect 172716 79870 172898 79930
rect 172716 79868 172717 79870
rect 172651 79867 172717 79868
rect 171915 79660 171981 79661
rect 171915 79596 171916 79660
rect 171980 79596 171981 79660
rect 171915 79595 171981 79596
rect 172099 79660 172165 79661
rect 172099 79596 172100 79660
rect 172164 79596 172165 79660
rect 172099 79595 172165 79596
rect 170995 79116 171061 79117
rect 170995 79052 170996 79116
rect 171060 79052 171061 79116
rect 170995 79051 171061 79052
rect 170998 78510 171242 78570
rect 170998 78437 171058 78510
rect 170995 78436 171061 78437
rect 170995 78372 170996 78436
rect 171060 78372 171061 78436
rect 170995 78371 171061 78372
rect 170811 78300 170877 78301
rect 170811 78236 170812 78300
rect 170876 78236 170877 78300
rect 170811 78235 170877 78236
rect 170627 76260 170693 76261
rect 170627 76196 170628 76260
rect 170692 76196 170693 76260
rect 170627 76195 170693 76196
rect 170443 75172 170509 75173
rect 170443 75108 170444 75172
rect 170508 75108 170509 75172
rect 170443 75107 170509 75108
rect 169523 29612 169589 29613
rect 169523 29548 169524 29612
rect 169588 29548 169589 29612
rect 169523 29547 169589 29548
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168051 6220 168117 6221
rect 168051 6156 168052 6220
rect 168116 6156 168117 6220
rect 168051 6155 168117 6156
rect 166763 5132 166829 5133
rect 166763 5068 166764 5132
rect 166828 5068 166829 5132
rect 166763 5067 166829 5068
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 -5146 168914 25398
rect 170814 4861 170874 78235
rect 171182 77349 171242 78510
rect 171918 78165 171978 79595
rect 172838 79250 172898 79870
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 173387 79252 173453 79253
rect 173387 79250 173388 79252
rect 172838 79190 173388 79250
rect 173387 79188 173388 79190
rect 173452 79188 173453 79252
rect 173387 79187 173453 79188
rect 171731 78164 171797 78165
rect 171731 78100 171732 78164
rect 171796 78100 171797 78164
rect 171731 78099 171797 78100
rect 171915 78164 171981 78165
rect 171915 78100 171916 78164
rect 171980 78100 171981 78164
rect 171915 78099 171981 78100
rect 171179 77348 171245 77349
rect 171179 77284 171180 77348
rect 171244 77284 171245 77348
rect 171179 77283 171245 77284
rect 170995 76396 171061 76397
rect 170995 76332 170996 76396
rect 171060 76332 171061 76396
rect 170995 76331 171061 76332
rect 170998 4997 171058 76331
rect 171734 42125 171794 78099
rect 172099 77756 172165 77757
rect 172099 77692 172100 77756
rect 172164 77692 172165 77756
rect 172099 77691 172165 77692
rect 171915 77484 171981 77485
rect 171915 77420 171916 77484
rect 171980 77420 171981 77484
rect 171915 77419 171981 77420
rect 171918 47565 171978 77419
rect 172102 48925 172162 77691
rect 172283 77348 172349 77349
rect 172283 77284 172284 77348
rect 172348 77284 172349 77348
rect 172283 77283 172349 77284
rect 172286 61437 172346 77283
rect 172794 66454 173414 78000
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172283 61436 172349 61437
rect 172283 61372 172284 61436
rect 172348 61372 172349 61436
rect 172283 61371 172349 61372
rect 172099 48924 172165 48925
rect 172099 48860 172100 48924
rect 172164 48860 172165 48924
rect 172099 48859 172165 48860
rect 171915 47564 171981 47565
rect 171915 47500 171916 47564
rect 171980 47500 171981 47564
rect 171915 47499 171981 47500
rect 171731 42124 171797 42125
rect 171731 42060 171732 42124
rect 171796 42060 171797 42124
rect 171731 42059 171797 42060
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 170995 4996 171061 4997
rect 170995 4932 170996 4996
rect 171060 4932 171061 4996
rect 170995 4931 171061 4932
rect 170811 4860 170877 4861
rect 170811 4796 170812 4860
rect 170876 4796 170877 4860
rect 170811 4795 170877 4796
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 70954 177914 78000
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 75454 182414 78000
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 228454 191414 263898
rect 190794 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 191414 228454
rect 190794 228134 191414 228218
rect 190794 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 191414 228134
rect 190794 192454 191414 227898
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 232954 195914 268398
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 241954 204914 277398
rect 204294 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 204914 241954
rect 204294 241634 204914 241718
rect 204294 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 204914 241634
rect 204294 205954 204914 241398
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 210454 209414 245898
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 214954 213914 250398
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 223954 222914 259398
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 151954 222914 187398
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 228454 227414 263898
rect 226794 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 227414 228454
rect 226794 228134 227414 228218
rect 226794 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 227414 228134
rect 226794 192454 227414 227898
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 376954 231914 412398
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 232954 231914 268398
rect 231294 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 231914 232954
rect 231294 232634 231914 232718
rect 231294 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 231914 232634
rect 231294 196954 231914 232398
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 124954 231914 160398
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 457954 240914 493398
rect 240294 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 240914 457954
rect 240294 457634 240914 457718
rect 240294 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 240914 457634
rect 240294 421954 240914 457398
rect 240294 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 240914 421954
rect 240294 421634 240914 421718
rect 240294 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 240914 421634
rect 240294 385954 240914 421398
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 349954 240914 385398
rect 240294 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 240914 349954
rect 240294 349634 240914 349718
rect 240294 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 240914 349634
rect 240294 313954 240914 349398
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 241954 240914 277398
rect 240294 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 240914 241954
rect 240294 241634 240914 241718
rect 240294 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 240914 241634
rect 240294 205954 240914 241398
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 426454 245414 461898
rect 244794 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 245414 426454
rect 244794 426134 245414 426218
rect 244794 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 245414 426134
rect 244794 390454 245414 425898
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 354454 245414 389898
rect 244794 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 245414 354454
rect 244794 354134 245414 354218
rect 244794 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 245414 354134
rect 244794 318454 245414 353898
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 246454 245414 281898
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 210454 245414 245898
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 322954 249914 358398
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 214954 249914 250398
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 223954 258914 259398
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 228454 263414 263898
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 262794 192454 263414 227898
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 232954 267914 268398
rect 267294 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 267914 232954
rect 267294 232634 267914 232718
rect 267294 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 267914 232634
rect 267294 196954 267914 232398
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 241954 276914 277398
rect 276294 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 276914 241954
rect 276294 241634 276914 241718
rect 276294 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 276914 241634
rect 276294 205954 276914 241398
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 210454 281414 245898
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 214954 285914 250398
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 223954 294914 259398
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 298794 372454 299414 407898
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 298794 336454 299414 371898
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 228454 299414 263898
rect 298794 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 299414 228454
rect 298794 228134 299414 228218
rect 298794 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 299414 228134
rect 298794 192454 299414 227898
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 232954 303914 268398
rect 303294 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 303914 232954
rect 303294 232634 303914 232718
rect 303294 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 303914 232634
rect 303294 196954 303914 232398
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 124954 303914 160398
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 241954 312914 277398
rect 312294 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 312914 241954
rect 312294 241634 312914 241718
rect 312294 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 312914 241634
rect 312294 205954 312914 241398
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 169954 312914 205398
rect 312294 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 312914 169954
rect 312294 169634 312914 169718
rect 312294 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 312914 169634
rect 312294 133954 312914 169398
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 210454 317414 245898
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 174454 317414 209898
rect 316794 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 317414 174454
rect 316794 174134 317414 174218
rect 316794 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 317414 174134
rect 316794 138454 317414 173898
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 214954 321914 250398
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 321294 178954 321914 214398
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 142954 321914 178398
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 223954 330914 259398
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 330294 187954 330914 223398
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 330294 151954 330914 187398
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 228454 335414 263898
rect 334794 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 335414 228454
rect 334794 228134 335414 228218
rect 334794 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 335414 228134
rect 334794 192454 335414 227898
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 334794 156454 335414 191898
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 376954 339914 412398
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 232954 339914 268398
rect 339294 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 339914 232954
rect 339294 232634 339914 232718
rect 339294 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 339914 232634
rect 339294 196954 339914 232398
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 124954 339914 160398
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 385954 348914 421398
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 241954 348914 277398
rect 348294 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 348914 241954
rect 348294 241634 348914 241718
rect 348294 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 348914 241634
rect 348294 205954 348914 241398
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 210454 353414 245898
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 214954 357914 250398
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 100826 246218 101062 246454
rect 101146 246218 101382 246454
rect 100826 245898 101062 246134
rect 101146 245898 101382 246134
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 118826 228218 119062 228454
rect 119146 228218 119382 228454
rect 118826 227898 119062 228134
rect 119146 227898 119382 228134
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 123326 232718 123562 232954
rect 123646 232718 123882 232954
rect 123326 232398 123562 232634
rect 123646 232398 123882 232634
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 132326 241718 132562 241954
rect 132646 241718 132882 241954
rect 132326 241398 132562 241634
rect 132646 241398 132882 241634
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 132326 169718 132562 169954
rect 132646 169718 132882 169954
rect 132326 169398 132562 169634
rect 132646 169398 132882 169634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 136826 246218 137062 246454
rect 137146 246218 137382 246454
rect 136826 245898 137062 246134
rect 137146 245898 137382 246134
rect 136826 210218 137062 210454
rect 137146 210218 137382 210454
rect 136826 209898 137062 210134
rect 137146 209898 137382 210134
rect 136826 174218 137062 174454
rect 137146 174218 137382 174454
rect 136826 173898 137062 174134
rect 137146 173898 137382 174134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 141326 214718 141562 214954
rect 141646 214718 141882 214954
rect 141326 214398 141562 214634
rect 141646 214398 141882 214634
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 141326 142718 141562 142954
rect 141646 142718 141882 142954
rect 141326 142398 141562 142634
rect 141646 142398 141882 142634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 150326 223718 150562 223954
rect 150646 223718 150882 223954
rect 150326 223398 150562 223634
rect 150646 223398 150882 223634
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 150326 151718 150562 151954
rect 150646 151718 150882 151954
rect 150326 151398 150562 151634
rect 150646 151398 150882 151634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 154826 228218 155062 228454
rect 155146 228218 155382 228454
rect 154826 227898 155062 228134
rect 155146 227898 155382 228134
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 159326 232718 159562 232954
rect 159646 232718 159882 232954
rect 159326 232398 159562 232634
rect 159646 232398 159882 232634
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 159326 160718 159562 160954
rect 159646 160718 159882 160954
rect 159326 160398 159562 160634
rect 159646 160398 159882 160634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 168326 241718 168562 241954
rect 168646 241718 168882 241954
rect 168326 241398 168562 241634
rect 168646 241398 168882 241634
rect 168326 205718 168562 205954
rect 168646 205718 168882 205954
rect 168326 205398 168562 205634
rect 168646 205398 168882 205634
rect 168326 169718 168562 169954
rect 168646 169718 168882 169954
rect 168326 169398 168562 169634
rect 168646 169398 168882 169634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 172826 246218 173062 246454
rect 173146 246218 173382 246454
rect 172826 245898 173062 246134
rect 173146 245898 173382 246134
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 139610 115718 139846 115954
rect 139610 115398 139846 115634
rect 170330 115718 170566 115954
rect 170330 115398 170566 115634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 124250 111218 124486 111454
rect 124250 110898 124486 111134
rect 154970 111218 155206 111454
rect 154970 110898 155206 111134
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 190826 228218 191062 228454
rect 191146 228218 191382 228454
rect 190826 227898 191062 228134
rect 191146 227898 191382 228134
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 204326 241718 204562 241954
rect 204646 241718 204882 241954
rect 204326 241398 204562 241634
rect 204646 241398 204882 241634
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 226826 228218 227062 228454
rect 227146 228218 227382 228454
rect 226826 227898 227062 228134
rect 227146 227898 227382 228134
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 231326 232718 231562 232954
rect 231646 232718 231882 232954
rect 231326 232398 231562 232634
rect 231646 232398 231882 232634
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 240326 457718 240562 457954
rect 240646 457718 240882 457954
rect 240326 457398 240562 457634
rect 240646 457398 240882 457634
rect 240326 421718 240562 421954
rect 240646 421718 240882 421954
rect 240326 421398 240562 421634
rect 240646 421398 240882 421634
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 240326 349718 240562 349954
rect 240646 349718 240882 349954
rect 240326 349398 240562 349634
rect 240646 349398 240882 349634
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 240326 241718 240562 241954
rect 240646 241718 240882 241954
rect 240326 241398 240562 241634
rect 240646 241398 240882 241634
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 244826 426218 245062 426454
rect 245146 426218 245382 426454
rect 244826 425898 245062 426134
rect 245146 425898 245382 426134
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 244826 354218 245062 354454
rect 245146 354218 245382 354454
rect 244826 353898 245062 354134
rect 245146 353898 245382 354134
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 267326 232718 267562 232954
rect 267646 232718 267882 232954
rect 267326 232398 267562 232634
rect 267646 232398 267882 232634
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 276326 241718 276562 241954
rect 276646 241718 276882 241954
rect 276326 241398 276562 241634
rect 276646 241398 276882 241634
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 298826 228218 299062 228454
rect 299146 228218 299382 228454
rect 298826 227898 299062 228134
rect 299146 227898 299382 228134
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 303326 232718 303562 232954
rect 303646 232718 303882 232954
rect 303326 232398 303562 232634
rect 303646 232398 303882 232634
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 312326 241718 312562 241954
rect 312646 241718 312882 241954
rect 312326 241398 312562 241634
rect 312646 241398 312882 241634
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 312326 169718 312562 169954
rect 312646 169718 312882 169954
rect 312326 169398 312562 169634
rect 312646 169398 312882 169634
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 316826 174218 317062 174454
rect 317146 174218 317382 174454
rect 316826 173898 317062 174134
rect 317146 173898 317382 174134
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 334826 228218 335062 228454
rect 335146 228218 335382 228454
rect 334826 227898 335062 228134
rect 335146 227898 335382 228134
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 339326 232718 339562 232954
rect 339646 232718 339882 232954
rect 339326 232398 339562 232634
rect 339646 232398 339882 232634
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 348326 241718 348562 241954
rect 348646 241718 348882 241954
rect 348326 241398 348562 241634
rect 348646 241398 348882 241634
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 139610 115954
rect 139846 115718 170330 115954
rect 170566 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 139610 115634
rect 139846 115398 170330 115634
rect 170566 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 124250 111454
rect 124486 111218 154970 111454
rect 155206 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 124250 111134
rect 124486 110898 154970 111134
rect 155206 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use rlbp_macro  rlbp_macro0
timestamp 0
transform 1 0 120000 0 1 80000
box 0 0 60000 60000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 78000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 142000 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 78000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 142000 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 142000 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 142000 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 78000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 142000 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 78000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 142000 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 78000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 142000 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 78000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 142000 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 78000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 142000 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 78000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 142000 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 78000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 142000 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 78000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 142000 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 78000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 142000 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 78000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 142000 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 78000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 142000 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
